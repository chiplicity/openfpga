magic
tech sky130A
magscale 1 2
timestamp 1605123412
<< locali >>
rect 3341 9911 3375 10149
rect 13737 9435 13771 9605
rect 8677 8347 8711 8585
rect 17693 4063 17727 4233
<< viali >>
rect 1593 24361 1627 24395
rect 1409 24225 1443 24259
rect 2329 23817 2363 23851
rect 2697 23817 2731 23851
rect 3801 23817 3835 23851
rect 19993 23817 20027 23851
rect 1409 23613 1443 23647
rect 2513 23613 2547 23647
rect 3065 23613 3099 23647
rect 3617 23613 3651 23647
rect 1593 23477 1627 23511
rect 2053 23477 2087 23511
rect 4261 23477 4295 23511
rect 8309 23273 8343 23307
rect 1961 23205 1995 23239
rect 1685 23137 1719 23171
rect 8125 23137 8159 23171
rect 4261 22729 4295 22763
rect 7481 22729 7515 22763
rect 8217 22729 8251 22763
rect 1869 22593 1903 22627
rect 8953 22593 8987 22627
rect 1685 22525 1719 22559
rect 2973 22525 3007 22559
rect 3525 22525 3559 22559
rect 4077 22525 4111 22559
rect 7297 22525 7331 22559
rect 8769 22525 8803 22559
rect 2513 22389 2547 22423
rect 2881 22389 2915 22423
rect 3157 22389 3191 22423
rect 4721 22389 4755 22423
rect 7941 22389 7975 22423
rect 9597 22389 9631 22423
rect 1409 22049 1443 22083
rect 2513 22049 2547 22083
rect 4077 22049 4111 22083
rect 5457 22049 5491 22083
rect 8125 22049 8159 22083
rect 1961 21981 1995 22015
rect 8309 21981 8343 22015
rect 1593 21913 1627 21947
rect 4261 21913 4295 21947
rect 5641 21913 5675 21947
rect 2329 21845 2363 21879
rect 2697 21845 2731 21879
rect 4905 21641 4939 21675
rect 5273 21641 5307 21675
rect 6009 21641 6043 21675
rect 1869 21505 1903 21539
rect 8125 21505 8159 21539
rect 1593 21437 1627 21471
rect 2881 21437 2915 21471
rect 3433 21437 3467 21471
rect 3985 21437 4019 21471
rect 4537 21437 4571 21471
rect 5089 21437 5123 21471
rect 5641 21437 5675 21471
rect 7941 21437 7975 21471
rect 8677 21437 8711 21471
rect 2513 21301 2547 21335
rect 3065 21301 3099 21335
rect 4169 21301 4203 21335
rect 7849 21301 7883 21335
rect 9229 21301 9263 21335
rect 9689 21097 9723 21131
rect 10057 21097 10091 21131
rect 1961 21029 1995 21063
rect 4445 21029 4479 21063
rect 6377 21029 6411 21063
rect 1685 20961 1719 20995
rect 4169 20961 4203 20995
rect 6101 20961 6135 20995
rect 7389 20893 7423 20927
rect 10149 20893 10183 20927
rect 10333 20893 10367 20927
rect 6929 20757 6963 20791
rect 10057 20553 10091 20587
rect 10425 20553 10459 20587
rect 9781 20485 9815 20519
rect 1961 20417 1995 20451
rect 3157 20417 3191 20451
rect 4537 20417 4571 20451
rect 1685 20349 1719 20383
rect 2421 20349 2455 20383
rect 2973 20349 3007 20383
rect 4261 20349 4295 20383
rect 5549 20349 5583 20383
rect 6101 20349 6135 20383
rect 6837 20349 6871 20383
rect 2789 20281 2823 20315
rect 6561 20281 6595 20315
rect 7082 20281 7116 20315
rect 3709 20213 3743 20247
rect 4169 20213 4203 20247
rect 5089 20213 5123 20247
rect 5365 20213 5399 20247
rect 5733 20213 5767 20247
rect 8217 20213 8251 20247
rect 8585 20213 8619 20247
rect 4905 20009 4939 20043
rect 6285 20009 6319 20043
rect 11069 20009 11103 20043
rect 1685 19941 1719 19975
rect 2973 19941 3007 19975
rect 4629 19941 4663 19975
rect 9934 19941 9968 19975
rect 1409 19873 1443 19907
rect 2697 19873 2731 19907
rect 3893 19873 3927 19907
rect 5273 19873 5307 19907
rect 7656 19873 7690 19907
rect 5365 19805 5399 19839
rect 5457 19805 5491 19839
rect 7389 19805 7423 19839
rect 9689 19805 9723 19839
rect 2145 19669 2179 19703
rect 2513 19669 2547 19703
rect 3525 19669 3559 19703
rect 4261 19669 4295 19703
rect 6009 19669 6043 19703
rect 6929 19669 6963 19703
rect 7297 19669 7331 19703
rect 8769 19669 8803 19703
rect 9045 19669 9079 19703
rect 9413 19669 9447 19703
rect 2329 19465 2363 19499
rect 4721 19465 4755 19499
rect 5181 19465 5215 19499
rect 6837 19465 6871 19499
rect 10609 19465 10643 19499
rect 8217 19397 8251 19431
rect 2697 19329 2731 19363
rect 4169 19329 4203 19363
rect 5641 19329 5675 19363
rect 5825 19329 5859 19363
rect 6193 19329 6227 19363
rect 7297 19329 7331 19363
rect 7389 19329 7423 19363
rect 11161 19329 11195 19363
rect 1593 19261 1627 19295
rect 1869 19261 1903 19295
rect 2881 19261 2915 19295
rect 3617 19261 3651 19295
rect 6653 19261 6687 19295
rect 7205 19261 7239 19295
rect 8401 19261 8435 19295
rect 8657 19261 8691 19295
rect 10517 19261 10551 19295
rect 11069 19261 11103 19295
rect 3157 19193 3191 19227
rect 4077 19193 4111 19227
rect 5089 19125 5123 19159
rect 5549 19125 5583 19159
rect 7941 19125 7975 19159
rect 9781 19125 9815 19159
rect 10149 19125 10183 19159
rect 10977 19125 11011 19159
rect 4997 18921 5031 18955
rect 6653 18921 6687 18955
rect 7481 18921 7515 18955
rect 9505 18921 9539 18955
rect 9689 18921 9723 18955
rect 10701 18853 10735 18887
rect 2329 18785 2363 18819
rect 4077 18785 4111 18819
rect 5540 18785 5574 18819
rect 7849 18785 7883 18819
rect 7941 18785 7975 18819
rect 10057 18785 10091 18819
rect 2421 18717 2455 18751
rect 2513 18717 2547 18751
rect 5273 18717 5307 18751
rect 8125 18717 8159 18751
rect 10149 18717 10183 18751
rect 10333 18717 10367 18751
rect 1869 18649 1903 18683
rect 1961 18581 1995 18615
rect 2973 18581 3007 18615
rect 3709 18581 3743 18615
rect 4261 18581 4295 18615
rect 7297 18581 7331 18615
rect 8493 18581 8527 18615
rect 8861 18581 8895 18615
rect 3617 18377 3651 18411
rect 5181 18377 5215 18411
rect 7205 18377 7239 18411
rect 9229 18377 9263 18411
rect 10977 18377 11011 18411
rect 10701 18309 10735 18343
rect 2605 18241 2639 18275
rect 4169 18241 4203 18275
rect 5825 18241 5859 18275
rect 6285 18241 6319 18275
rect 7757 18241 7791 18275
rect 8309 18173 8343 18207
rect 9321 18173 9355 18207
rect 9588 18173 9622 18207
rect 1869 18105 1903 18139
rect 3433 18105 3467 18139
rect 3985 18105 4019 18139
rect 5089 18105 5123 18139
rect 6653 18105 6687 18139
rect 7573 18105 7607 18139
rect 8861 18105 8895 18139
rect 1961 18037 1995 18071
rect 2329 18037 2363 18071
rect 2421 18037 2455 18071
rect 2973 18037 3007 18071
rect 4077 18037 4111 18071
rect 4629 18037 4663 18071
rect 5549 18037 5583 18071
rect 5641 18037 5675 18071
rect 7113 18037 7147 18071
rect 7665 18037 7699 18071
rect 11437 18037 11471 18071
rect 1409 17833 1443 17867
rect 5825 17833 5859 17867
rect 7665 17833 7699 17867
rect 8309 17833 8343 17867
rect 8585 17833 8619 17867
rect 9413 17833 9447 17867
rect 11161 17833 11195 17867
rect 3525 17765 3559 17799
rect 2789 17697 2823 17731
rect 4333 17697 4367 17731
rect 6541 17697 6575 17731
rect 10037 17697 10071 17731
rect 2881 17629 2915 17663
rect 2973 17629 3007 17663
rect 3801 17629 3835 17663
rect 4077 17629 4111 17663
rect 6285 17629 6319 17663
rect 9781 17629 9815 17663
rect 2421 17561 2455 17595
rect 7941 17561 7975 17595
rect 1961 17493 1995 17527
rect 5457 17493 5491 17527
rect 6193 17493 6227 17527
rect 4997 17289 5031 17323
rect 9689 17289 9723 17323
rect 4169 17221 4203 17255
rect 9321 17221 9355 17255
rect 5549 17153 5583 17187
rect 6009 17153 6043 17187
rect 6377 17153 6411 17187
rect 10333 17153 10367 17187
rect 11253 17153 11287 17187
rect 1409 17085 1443 17119
rect 1685 17085 1719 17119
rect 2789 17085 2823 17119
rect 6837 17085 6871 17119
rect 9505 17085 9539 17119
rect 11069 17085 11103 17119
rect 3056 17017 3090 17051
rect 5365 17017 5399 17051
rect 7104 17017 7138 17051
rect 8493 17017 8527 17051
rect 9229 17017 9263 17051
rect 10057 17017 10091 17051
rect 2513 16949 2547 16983
rect 4537 16949 4571 16983
rect 4905 16949 4939 16983
rect 5457 16949 5491 16983
rect 8217 16949 8251 16983
rect 10149 16949 10183 16983
rect 10701 16949 10735 16983
rect 11805 16949 11839 16983
rect 2145 16745 2179 16779
rect 3433 16745 3467 16779
rect 4077 16745 4111 16779
rect 7205 16745 7239 16779
rect 8033 16745 8067 16779
rect 9505 16745 9539 16779
rect 11345 16745 11379 16779
rect 2789 16677 2823 16711
rect 3065 16677 3099 16711
rect 6092 16677 6126 16711
rect 7481 16677 7515 16711
rect 7941 16677 7975 16711
rect 2053 16609 2087 16643
rect 3893 16609 3927 16643
rect 4445 16609 4479 16643
rect 5825 16609 5859 16643
rect 8401 16609 8435 16643
rect 10221 16609 10255 16643
rect 2237 16541 2271 16575
rect 4537 16541 4571 16575
rect 4629 16541 4663 16575
rect 8493 16541 8527 16575
rect 8677 16541 8711 16575
rect 9965 16541 9999 16575
rect 3709 16473 3743 16507
rect 5181 16473 5215 16507
rect 1685 16405 1719 16439
rect 5457 16405 5491 16439
rect 9137 16405 9171 16439
rect 2237 16201 2271 16235
rect 4169 16201 4203 16235
rect 5089 16201 5123 16235
rect 6101 16201 6135 16235
rect 10241 16201 10275 16235
rect 1685 16065 1719 16099
rect 5733 16065 5767 16099
rect 9413 16065 9447 16099
rect 10793 16065 10827 16099
rect 12449 16065 12483 16099
rect 1409 15997 1443 16031
rect 2789 15997 2823 16031
rect 4905 15997 4939 16031
rect 7389 15997 7423 16031
rect 7645 15997 7679 16031
rect 2697 15929 2731 15963
rect 3034 15929 3068 15963
rect 5549 15929 5583 15963
rect 10149 15929 10183 15963
rect 10701 15929 10735 15963
rect 4537 15861 4571 15895
rect 5457 15861 5491 15895
rect 6561 15861 6595 15895
rect 7297 15861 7331 15895
rect 8769 15861 8803 15895
rect 9781 15861 9815 15895
rect 10609 15861 10643 15895
rect 11253 15861 11287 15895
rect 11713 15861 11747 15895
rect 12081 15861 12115 15895
rect 2421 15657 2455 15691
rect 3801 15657 3835 15691
rect 4077 15657 4111 15691
rect 4537 15657 4571 15691
rect 6745 15657 6779 15691
rect 7297 15657 7331 15691
rect 8677 15657 8711 15691
rect 10057 15657 10091 15691
rect 11713 15657 11747 15691
rect 2329 15589 2363 15623
rect 4997 15589 5031 15623
rect 5334 15589 5368 15623
rect 10600 15589 10634 15623
rect 1409 15521 1443 15555
rect 2789 15521 2823 15555
rect 5089 15521 5123 15555
rect 7665 15521 7699 15555
rect 9321 15521 9355 15555
rect 10333 15521 10367 15555
rect 2881 15453 2915 15487
rect 2973 15453 3007 15487
rect 7757 15453 7791 15487
rect 7849 15453 7883 15487
rect 3525 15385 3559 15419
rect 1961 15317 1995 15351
rect 6469 15317 6503 15351
rect 7113 15317 7147 15351
rect 8401 15317 8435 15351
rect 9137 15317 9171 15351
rect 12081 15317 12115 15351
rect 12541 15317 12575 15351
rect 2053 15113 2087 15147
rect 3065 15113 3099 15147
rect 3617 15113 3651 15147
rect 5181 15113 5215 15147
rect 9965 15113 9999 15147
rect 11069 15113 11103 15147
rect 2605 14977 2639 15011
rect 4169 14977 4203 15011
rect 5733 14977 5767 15011
rect 6193 14977 6227 15011
rect 7757 14977 7791 15011
rect 10609 14977 10643 15011
rect 11897 14977 11931 15011
rect 13001 14977 13035 15011
rect 2421 14909 2455 14943
rect 12817 14909 12851 14943
rect 1961 14841 1995 14875
rect 2513 14841 2547 14875
rect 4077 14841 4111 14875
rect 5089 14841 5123 14875
rect 6653 14841 6687 14875
rect 8024 14841 8058 14875
rect 9505 14841 9539 14875
rect 10425 14841 10459 14875
rect 12173 14841 12207 14875
rect 12909 14841 12943 14875
rect 3525 14773 3559 14807
rect 3985 14773 4019 14807
rect 4629 14773 4663 14807
rect 5549 14773 5583 14807
rect 5641 14773 5675 14807
rect 7297 14773 7331 14807
rect 9137 14773 9171 14807
rect 9873 14773 9907 14807
rect 10333 14773 10367 14807
rect 11437 14773 11471 14807
rect 12449 14773 12483 14807
rect 1409 14569 1443 14603
rect 2421 14569 2455 14603
rect 3801 14569 3835 14603
rect 4261 14569 4295 14603
rect 6377 14569 6411 14603
rect 7205 14569 7239 14603
rect 8677 14569 8711 14603
rect 8769 14569 8803 14603
rect 9321 14569 9355 14603
rect 11621 14569 11655 14603
rect 11897 14569 11931 14603
rect 12265 14569 12299 14603
rect 12449 14569 12483 14603
rect 2145 14501 2179 14535
rect 2881 14501 2915 14535
rect 7573 14501 7607 14535
rect 8309 14501 8343 14535
rect 10057 14501 10091 14535
rect 10508 14501 10542 14535
rect 12817 14501 12851 14535
rect 2789 14433 2823 14467
rect 3433 14433 3467 14467
rect 4997 14433 5031 14467
rect 5264 14433 5298 14467
rect 8953 14433 8987 14467
rect 10241 14433 10275 14467
rect 23489 14433 23523 14467
rect 3065 14365 3099 14399
rect 4721 14365 4755 14399
rect 7665 14365 7699 14399
rect 7849 14365 7883 14399
rect 12909 14365 12943 14399
rect 13001 14365 13035 14399
rect 6653 14229 6687 14263
rect 7021 14229 7055 14263
rect 23673 14229 23707 14263
rect 3341 14025 3375 14059
rect 4077 14025 4111 14059
rect 6653 14025 6687 14059
rect 10057 14025 10091 14059
rect 11805 14025 11839 14059
rect 12265 14025 12299 14059
rect 13277 14025 13311 14059
rect 23489 14025 23523 14059
rect 5181 13957 5215 13991
rect 23857 13957 23891 13991
rect 1869 13889 1903 13923
rect 3709 13889 3743 13923
rect 5089 13889 5123 13923
rect 5825 13889 5859 13923
rect 9597 13889 9631 13923
rect 10609 13889 10643 13923
rect 1961 13821 1995 13855
rect 4721 13821 4755 13855
rect 7297 13821 7331 13855
rect 7757 13821 7791 13855
rect 7849 13821 7883 13855
rect 8116 13821 8150 13855
rect 12909 13821 12943 13855
rect 23673 13821 23707 13855
rect 24225 13821 24259 13855
rect 2228 13753 2262 13787
rect 4169 13753 4203 13787
rect 5641 13753 5675 13787
rect 9873 13753 9907 13787
rect 10517 13753 10551 13787
rect 5549 13685 5583 13719
rect 6285 13685 6319 13719
rect 6837 13685 6871 13719
rect 9229 13685 9263 13719
rect 10425 13685 10459 13719
rect 11161 13685 11195 13719
rect 11529 13685 11563 13719
rect 12449 13685 12483 13719
rect 3157 13481 3191 13515
rect 4261 13481 4295 13515
rect 5273 13481 5307 13515
rect 7573 13481 7607 13515
rect 8861 13481 8895 13515
rect 9137 13481 9171 13515
rect 10057 13481 10091 13515
rect 11621 13481 11655 13515
rect 11897 13481 11931 13515
rect 2022 13413 2056 13447
rect 3433 13413 3467 13447
rect 10508 13413 10542 13447
rect 1777 13345 1811 13379
rect 4077 13345 4111 13379
rect 5632 13345 5666 13379
rect 7941 13345 7975 13379
rect 9321 13345 9355 13379
rect 10241 13345 10275 13379
rect 22293 13345 22327 13379
rect 3893 13277 3927 13311
rect 5365 13277 5399 13311
rect 8033 13277 8067 13311
rect 8217 13277 8251 13311
rect 6745 13209 6779 13243
rect 1685 13141 1719 13175
rect 4721 13141 4755 13175
rect 7205 13141 7239 13175
rect 12357 13141 12391 13175
rect 12633 13141 12667 13175
rect 22477 13141 22511 13175
rect 2513 12937 2547 12971
rect 4721 12937 4755 12971
rect 11161 12937 11195 12971
rect 11437 12937 11471 12971
rect 11989 12937 12023 12971
rect 5457 12869 5491 12903
rect 8585 12869 8619 12903
rect 11897 12869 11931 12903
rect 2145 12801 2179 12835
rect 2881 12801 2915 12835
rect 7665 12801 7699 12835
rect 9781 12801 9815 12835
rect 1961 12733 1995 12767
rect 3065 12733 3099 12767
rect 3332 12733 3366 12767
rect 5273 12733 5307 12767
rect 12173 12733 12207 12767
rect 12633 12733 12667 12767
rect 13001 12733 13035 12767
rect 22293 12733 22327 12767
rect 6193 12665 6227 12699
rect 6653 12665 6687 12699
rect 7481 12665 7515 12699
rect 9229 12665 9263 12699
rect 9689 12665 9723 12699
rect 10048 12665 10082 12699
rect 1501 12597 1535 12631
rect 1869 12597 1903 12631
rect 4445 12597 4479 12631
rect 5089 12597 5123 12631
rect 5917 12597 5951 12631
rect 7113 12597 7147 12631
rect 7573 12597 7607 12631
rect 8217 12597 8251 12631
rect 8769 12597 8803 12631
rect 3433 12393 3467 12427
rect 4261 12393 4295 12427
rect 5181 12393 5215 12427
rect 6929 12393 6963 12427
rect 7297 12393 7331 12427
rect 8033 12393 8067 12427
rect 8401 12393 8435 12427
rect 11069 12393 11103 12427
rect 9505 12325 9539 12359
rect 9956 12325 9990 12359
rect 1869 12257 1903 12291
rect 4077 12257 4111 12291
rect 5365 12257 5399 12291
rect 5816 12257 5850 12291
rect 9689 12257 9723 12291
rect 11713 12257 11747 12291
rect 12256 12257 12290 12291
rect 21741 12257 21775 12291
rect 1961 12189 1995 12223
rect 2145 12189 2179 12223
rect 3065 12189 3099 12223
rect 5549 12189 5583 12223
rect 8493 12189 8527 12223
rect 8677 12189 8711 12223
rect 9137 12189 9171 12223
rect 11989 12189 12023 12223
rect 1501 12053 1535 12087
rect 2789 12053 2823 12087
rect 3893 12053 3927 12087
rect 4629 12053 4663 12087
rect 5089 12053 5123 12087
rect 7665 12053 7699 12087
rect 11345 12053 11379 12087
rect 13369 12053 13403 12087
rect 21925 12053 21959 12087
rect 2697 11849 2731 11883
rect 4353 11849 4387 11883
rect 5917 11849 5951 11883
rect 7757 11849 7791 11883
rect 8125 11849 8159 11883
rect 13369 11849 13403 11883
rect 13737 11849 13771 11883
rect 14105 11849 14139 11883
rect 21741 11781 21775 11815
rect 1685 11713 1719 11747
rect 3249 11713 3283 11747
rect 3709 11713 3743 11747
rect 10701 11713 10735 11747
rect 1409 11645 1443 11679
rect 4537 11645 4571 11679
rect 4793 11645 4827 11679
rect 12725 11645 12759 11679
rect 2605 11577 2639 11611
rect 3157 11577 3191 11611
rect 6561 11577 6595 11611
rect 7389 11577 7423 11611
rect 8769 11577 8803 11611
rect 8861 11577 8895 11611
rect 10946 11577 10980 11611
rect 2237 11509 2271 11543
rect 3065 11509 3099 11543
rect 6285 11509 6319 11543
rect 6837 11509 6871 11543
rect 10149 11509 10183 11543
rect 12081 11509 12115 11543
rect 13093 11509 13127 11543
rect 3065 11305 3099 11339
rect 3341 11305 3375 11339
rect 4077 11305 4111 11339
rect 5273 11305 5307 11339
rect 7021 11305 7055 11339
rect 9689 11305 9723 11339
rect 11253 11305 11287 11339
rect 11713 11305 11747 11339
rect 12817 11305 12851 11339
rect 5908 11237 5942 11271
rect 7757 11237 7791 11271
rect 8116 11237 8150 11271
rect 1685 11169 1719 11203
rect 1941 11169 1975 11203
rect 4445 11169 4479 11203
rect 5641 11169 5675 11203
rect 7849 11169 7883 11203
rect 10057 11169 10091 11203
rect 11069 11169 11103 11203
rect 11621 11169 11655 11203
rect 13185 11169 13219 11203
rect 13277 11169 13311 11203
rect 3893 11101 3927 11135
rect 4537 11101 4571 11135
rect 4629 11101 4663 11135
rect 10149 11101 10183 11135
rect 10333 11101 10367 11135
rect 11805 11101 11839 11135
rect 13369 11101 13403 11135
rect 9229 11033 9263 11067
rect 10793 11033 10827 11067
rect 7389 10965 7423 10999
rect 12541 10965 12575 10999
rect 3065 10761 3099 10795
rect 4169 10761 4203 10795
rect 5641 10761 5675 10795
rect 6009 10761 6043 10795
rect 7297 10761 7331 10795
rect 7849 10761 7883 10795
rect 10701 10761 10735 10795
rect 12449 10761 12483 10795
rect 14197 10761 14231 10795
rect 7757 10693 7791 10727
rect 8401 10625 8435 10659
rect 9689 10625 9723 10659
rect 11253 10625 11287 10659
rect 12909 10625 12943 10659
rect 13093 10625 13127 10659
rect 13829 10625 13863 10659
rect 1409 10557 1443 10591
rect 1676 10557 1710 10591
rect 4261 10557 4295 10591
rect 8217 10557 8251 10591
rect 12173 10557 12207 10591
rect 12817 10557 12851 10591
rect 3801 10489 3835 10523
rect 4528 10489 4562 10523
rect 8309 10489 8343 10523
rect 9045 10489 9079 10523
rect 10609 10489 10643 10523
rect 2789 10421 2823 10455
rect 6561 10421 6595 10455
rect 9137 10421 9171 10455
rect 9505 10421 9539 10455
rect 9597 10421 9631 10455
rect 10149 10421 10183 10455
rect 11069 10421 11103 10455
rect 11161 10421 11195 10455
rect 11713 10421 11747 10455
rect 13461 10421 13495 10455
rect 1777 10217 1811 10251
rect 4077 10217 4111 10251
rect 5641 10217 5675 10251
rect 7573 10217 7607 10251
rect 7941 10217 7975 10251
rect 8677 10217 8711 10251
rect 9965 10217 9999 10251
rect 10333 10217 10367 10251
rect 12357 10217 12391 10251
rect 12909 10217 12943 10251
rect 2513 10149 2547 10183
rect 3065 10149 3099 10183
rect 3341 10149 3375 10183
rect 3525 10149 3559 10183
rect 6009 10149 6043 10183
rect 10793 10149 10827 10183
rect 2421 10081 2455 10115
rect 2605 10013 2639 10047
rect 4445 10081 4479 10115
rect 7113 10081 7147 10115
rect 8033 10081 8067 10115
rect 11244 10081 11278 10115
rect 4537 10013 4571 10047
rect 4721 10013 4755 10047
rect 6101 10013 6135 10047
rect 6193 10013 6227 10047
rect 7205 10013 7239 10047
rect 7297 10013 7331 10047
rect 8125 10013 8159 10047
rect 10977 10013 11011 10047
rect 13185 10013 13219 10047
rect 3801 9945 3835 9979
rect 6745 9945 6779 9979
rect 2053 9877 2087 9911
rect 3341 9877 3375 9911
rect 5181 9877 5215 9911
rect 5457 9877 5491 9911
rect 9137 9877 9171 9911
rect 13645 9877 13679 9911
rect 1685 9673 1719 9707
rect 3249 9673 3283 9707
rect 9597 9673 9631 9707
rect 11529 9673 11563 9707
rect 11805 9673 11839 9707
rect 4077 9605 4111 9639
rect 5457 9605 5491 9639
rect 12449 9605 12483 9639
rect 13737 9605 13771 9639
rect 1869 9537 1903 9571
rect 4721 9537 4755 9571
rect 5089 9537 5123 9571
rect 5641 9537 5675 9571
rect 13001 9537 13035 9571
rect 2136 9469 2170 9503
rect 4445 9469 4479 9503
rect 7573 9469 7607 9503
rect 10149 9469 10183 9503
rect 12173 9469 12207 9503
rect 12909 9469 12943 9503
rect 4537 9401 4571 9435
rect 7818 9401 7852 9435
rect 9229 9401 9263 9435
rect 10394 9401 10428 9435
rect 13737 9401 13771 9435
rect 13829 9401 13863 9435
rect 3525 9333 3559 9367
rect 3893 9333 3927 9367
rect 6101 9333 6135 9367
rect 6469 9333 6503 9367
rect 7113 9333 7147 9367
rect 7389 9333 7423 9367
rect 8953 9333 8987 9367
rect 10057 9333 10091 9367
rect 12817 9333 12851 9367
rect 13461 9333 13495 9367
rect 1501 9129 1535 9163
rect 1961 9129 1995 9163
rect 2605 9129 2639 9163
rect 2973 9129 3007 9163
rect 3617 9129 3651 9163
rect 6745 9129 6779 9163
rect 7297 9129 7331 9163
rect 9413 9129 9447 9163
rect 10425 9129 10459 9163
rect 12817 9129 12851 9163
rect 14013 9129 14047 9163
rect 4353 9061 4387 9095
rect 8401 9061 8435 9095
rect 12449 9061 12483 9095
rect 13369 9061 13403 9095
rect 1869 8993 1903 9027
rect 3893 8993 3927 9027
rect 4077 8993 4111 9027
rect 5621 8993 5655 9027
rect 7941 8993 7975 9027
rect 10793 8993 10827 9027
rect 11060 8993 11094 9027
rect 2053 8925 2087 8959
rect 5365 8925 5399 8959
rect 7665 8925 7699 8959
rect 8493 8925 8527 8959
rect 8585 8925 8619 8959
rect 9781 8925 9815 8959
rect 13461 8925 13495 8959
rect 13645 8925 13679 8959
rect 3709 8789 3743 8823
rect 4813 8789 4847 8823
rect 5273 8789 5307 8823
rect 7757 8789 7791 8823
rect 8033 8789 8067 8823
rect 9137 8789 9171 8823
rect 12173 8789 12207 8823
rect 13001 8789 13035 8823
rect 3341 8585 3375 8619
rect 3709 8585 3743 8619
rect 3985 8585 4019 8619
rect 4721 8585 4755 8619
rect 8309 8585 8343 8619
rect 8677 8585 8711 8619
rect 8861 8585 8895 8619
rect 11897 8585 11931 8619
rect 13829 8585 13863 8619
rect 5181 8517 5215 8551
rect 6837 8517 6871 8551
rect 8401 8517 8435 8551
rect 1961 8449 1995 8483
rect 4169 8449 4203 8483
rect 5089 8449 5123 8483
rect 5733 8449 5767 8483
rect 6285 8449 6319 8483
rect 7389 8449 7423 8483
rect 5549 8381 5583 8415
rect 8585 8381 8619 8415
rect 10425 8517 10459 8551
rect 12449 8517 12483 8551
rect 17141 8517 17175 8551
rect 9505 8449 9539 8483
rect 9965 8449 9999 8483
rect 10977 8449 11011 8483
rect 13001 8449 13035 8483
rect 14473 8449 14507 8483
rect 10793 8381 10827 8415
rect 11529 8381 11563 8415
rect 12265 8381 12299 8415
rect 12817 8381 12851 8415
rect 12909 8381 12943 8415
rect 14013 8381 14047 8415
rect 15761 8381 15795 8415
rect 2228 8313 2262 8347
rect 5641 8313 5675 8347
rect 7297 8313 7331 8347
rect 7941 8313 7975 8347
rect 8677 8313 8711 8347
rect 9229 8313 9263 8347
rect 10241 8313 10275 8347
rect 10885 8313 10919 8347
rect 16006 8313 16040 8347
rect 1869 8245 1903 8279
rect 6561 8245 6595 8279
rect 7205 8245 7239 8279
rect 9321 8245 9355 8279
rect 12081 8245 12115 8279
rect 13461 8245 13495 8279
rect 15669 8245 15703 8279
rect 3433 8041 3467 8075
rect 4353 8041 4387 8075
rect 4721 8041 4755 8075
rect 6193 8041 6227 8075
rect 6561 8041 6595 8075
rect 9873 8041 9907 8075
rect 12909 8041 12943 8075
rect 3801 7973 3835 8007
rect 5080 7973 5114 8007
rect 11428 7973 11462 8007
rect 14749 7973 14783 8007
rect 15761 7973 15795 8007
rect 1409 7905 1443 7939
rect 1676 7905 1710 7939
rect 3157 7905 3191 7939
rect 7472 7905 7506 7939
rect 11161 7905 11195 7939
rect 13737 7905 13771 7939
rect 4813 7837 4847 7871
rect 7205 7837 7239 7871
rect 10149 7837 10183 7871
rect 10793 7837 10827 7871
rect 13829 7837 13863 7871
rect 13921 7837 13955 7871
rect 16037 7837 16071 7871
rect 2789 7769 2823 7803
rect 12541 7769 12575 7803
rect 6929 7701 6963 7735
rect 8585 7701 8619 7735
rect 8953 7701 8987 7735
rect 9321 7701 9355 7735
rect 13185 7701 13219 7735
rect 13369 7701 13403 7735
rect 14381 7701 14415 7735
rect 1409 7497 1443 7531
rect 4629 7497 4663 7531
rect 6285 7497 6319 7531
rect 7389 7497 7423 7531
rect 9689 7497 9723 7531
rect 11897 7497 11931 7531
rect 13001 7497 13035 7531
rect 15117 7497 15151 7531
rect 15853 7497 15887 7531
rect 2053 7361 2087 7395
rect 5825 7361 5859 7395
rect 6837 7361 6871 7395
rect 8033 7361 8067 7395
rect 10149 7361 10183 7395
rect 11437 7361 11471 7395
rect 12541 7361 12575 7395
rect 13737 7361 13771 7395
rect 16497 7361 16531 7395
rect 1777 7293 1811 7327
rect 2789 7293 2823 7327
rect 2973 7293 3007 7327
rect 3229 7293 3263 7327
rect 5549 7293 5583 7327
rect 8300 7293 8334 7327
rect 10425 7293 10459 7327
rect 11161 7293 11195 7327
rect 11253 7293 11287 7327
rect 12173 7293 12207 7327
rect 16313 7293 16347 7327
rect 5089 7225 5123 7259
rect 5641 7225 5675 7259
rect 7941 7225 7975 7259
rect 14004 7225 14038 7259
rect 15485 7225 15519 7259
rect 1869 7157 1903 7191
rect 2513 7157 2547 7191
rect 4353 7157 4387 7191
rect 5181 7157 5215 7191
rect 6653 7157 6687 7191
rect 9413 7157 9447 7191
rect 10241 7157 10275 7191
rect 10793 7157 10827 7191
rect 13369 7157 13403 7191
rect 15945 7157 15979 7191
rect 16405 7157 16439 7191
rect 16957 7157 16991 7191
rect 2881 6953 2915 6987
rect 4077 6953 4111 6987
rect 4905 6953 4939 6987
rect 12909 6953 12943 6987
rect 14657 6953 14691 6987
rect 3893 6885 3927 6919
rect 1777 6817 1811 6851
rect 5365 6817 5399 6851
rect 5457 6817 5491 6851
rect 5724 6817 5758 6851
rect 7113 6817 7147 6851
rect 8125 6817 8159 6851
rect 8217 6817 8251 6851
rect 10324 6817 10358 6851
rect 12173 6817 12207 6851
rect 13257 6817 13291 6851
rect 15925 6817 15959 6851
rect 17877 6817 17911 6851
rect 1869 6749 1903 6783
rect 2053 6749 2087 6783
rect 2973 6749 3007 6783
rect 8401 6749 8435 6783
rect 10057 6749 10091 6783
rect 13001 6749 13035 6783
rect 15117 6749 15151 6783
rect 15676 6749 15710 6783
rect 18153 6749 18187 6783
rect 7757 6681 7791 6715
rect 1409 6613 1443 6647
rect 2421 6613 2455 6647
rect 3525 6613 3559 6647
rect 5181 6613 5215 6647
rect 6837 6613 6871 6647
rect 7481 6613 7515 6647
rect 8769 6613 8803 6647
rect 9137 6613 9171 6647
rect 9873 6613 9907 6647
rect 11437 6613 11471 6647
rect 11713 6613 11747 6647
rect 12449 6613 12483 6647
rect 14381 6613 14415 6647
rect 17049 6613 17083 6647
rect 1961 6409 1995 6443
rect 4997 6409 5031 6443
rect 6837 6409 6871 6443
rect 7941 6409 7975 6443
rect 8309 6409 8343 6443
rect 10149 6409 10183 6443
rect 10425 6409 10459 6443
rect 11713 6409 11747 6443
rect 15025 6409 15059 6443
rect 16405 6409 16439 6443
rect 18521 6409 18555 6443
rect 4077 6341 4111 6375
rect 5181 6341 5215 6375
rect 6285 6341 6319 6375
rect 2789 6273 2823 6307
rect 5641 6273 5675 6307
rect 5825 6273 5859 6307
rect 6653 6273 6687 6307
rect 7389 6273 7423 6307
rect 8677 6273 8711 6307
rect 12817 6273 12851 6307
rect 15669 6273 15703 6307
rect 7205 6205 7239 6239
rect 8769 6205 8803 6239
rect 9036 6205 9070 6239
rect 13084 6205 13118 6239
rect 15393 6205 15427 6239
rect 16589 6205 16623 6239
rect 17325 6205 17359 6239
rect 19533 6205 19567 6239
rect 20269 6205 20303 6239
rect 2605 6137 2639 6171
rect 3617 6137 3651 6171
rect 4169 6137 4203 6171
rect 4721 6137 4755 6171
rect 5549 6137 5583 6171
rect 7297 6137 7331 6171
rect 12725 6137 12759 6171
rect 15485 6137 15519 6171
rect 16865 6137 16899 6171
rect 19809 6137 19843 6171
rect 1593 6069 1627 6103
rect 2237 6069 2271 6103
rect 2697 6069 2731 6103
rect 3249 6069 3283 6103
rect 10793 6069 10827 6103
rect 11161 6069 11195 6103
rect 12265 6069 12299 6103
rect 14197 6069 14231 6103
rect 14841 6069 14875 6103
rect 16129 6069 16163 6103
rect 18061 6069 18095 6103
rect 1409 5865 1443 5899
rect 2421 5865 2455 5899
rect 2789 5865 2823 5899
rect 4629 5865 4663 5899
rect 5365 5865 5399 5899
rect 5733 5865 5767 5899
rect 7389 5865 7423 5899
rect 8217 5865 8251 5899
rect 8769 5865 8803 5899
rect 9137 5865 9171 5899
rect 13093 5865 13127 5899
rect 13737 5865 13771 5899
rect 17693 5865 17727 5899
rect 6254 5797 6288 5831
rect 11958 5797 11992 5831
rect 15025 5797 15059 5831
rect 3525 5729 3559 5763
rect 3893 5729 3927 5763
rect 6009 5729 6043 5763
rect 7849 5729 7883 5763
rect 10057 5729 10091 5763
rect 11161 5729 11195 5763
rect 11437 5729 11471 5763
rect 13921 5729 13955 5763
rect 16580 5729 16614 5763
rect 18521 5729 18555 5763
rect 19625 5729 19659 5763
rect 2881 5661 2915 5695
rect 2973 5661 3007 5695
rect 4721 5661 4755 5695
rect 4813 5661 4847 5695
rect 10149 5661 10183 5695
rect 10241 5661 10275 5695
rect 11713 5661 11747 5695
rect 14105 5661 14139 5695
rect 15301 5661 15335 5695
rect 16313 5661 16347 5695
rect 2329 5593 2363 5627
rect 9413 5593 9447 5627
rect 1961 5525 1995 5559
rect 4261 5525 4295 5559
rect 9689 5525 9723 5559
rect 10793 5525 10827 5559
rect 11253 5525 11287 5559
rect 13369 5525 13403 5559
rect 15761 5525 15795 5559
rect 16221 5525 16255 5559
rect 18705 5525 18739 5559
rect 19809 5525 19843 5559
rect 4629 5321 4663 5355
rect 5181 5321 5215 5355
rect 7941 5321 7975 5355
rect 8309 5321 8343 5355
rect 12449 5321 12483 5355
rect 13921 5321 13955 5355
rect 15025 5321 15059 5355
rect 18797 5321 18831 5355
rect 11805 5253 11839 5287
rect 5733 5185 5767 5219
rect 7389 5185 7423 5219
rect 8585 5185 8619 5219
rect 13001 5185 13035 5219
rect 13461 5185 13495 5219
rect 14565 5185 14599 5219
rect 16037 5185 16071 5219
rect 16773 5185 16807 5219
rect 1961 5117 1995 5151
rect 3709 5117 3743 5151
rect 5089 5117 5123 5151
rect 5641 5117 5675 5151
rect 7205 5117 7239 5151
rect 9597 5117 9631 5151
rect 12817 5117 12851 5151
rect 14381 5117 14415 5151
rect 17877 5117 17911 5151
rect 18061 5117 18095 5151
rect 19349 5117 19383 5151
rect 19901 5117 19935 5151
rect 20545 5117 20579 5151
rect 21097 5117 21131 5151
rect 2228 5049 2262 5083
rect 6653 5049 6687 5083
rect 7297 5049 7331 5083
rect 9137 5049 9171 5083
rect 9842 5049 9876 5083
rect 11253 5049 11287 5083
rect 14473 5049 14507 5083
rect 15669 5049 15703 5083
rect 16497 5049 16531 5083
rect 18337 5049 18371 5083
rect 1869 4981 1903 5015
rect 3341 4981 3375 5015
rect 4353 4981 4387 5015
rect 5549 4981 5583 5015
rect 6193 4981 6227 5015
rect 6837 4981 6871 5015
rect 9413 4981 9447 5015
rect 10977 4981 11011 5015
rect 12265 4981 12299 5015
rect 12909 4981 12943 5015
rect 14013 4981 14047 5015
rect 16129 4981 16163 5015
rect 16589 4981 16623 5015
rect 17233 4981 17267 5015
rect 19533 4981 19567 5015
rect 20361 4981 20395 5015
rect 20729 4981 20763 5015
rect 3157 4777 3191 4811
rect 3433 4777 3467 4811
rect 3893 4777 3927 4811
rect 6929 4777 6963 4811
rect 8033 4777 8067 4811
rect 9045 4777 9079 4811
rect 11621 4777 11655 4811
rect 12817 4777 12851 4811
rect 14105 4777 14139 4811
rect 14473 4777 14507 4811
rect 17417 4777 17451 4811
rect 2044 4709 2078 4743
rect 5794 4709 5828 4743
rect 13185 4709 13219 4743
rect 18061 4709 18095 4743
rect 8401 4641 8435 4675
rect 10057 4641 10091 4675
rect 11713 4641 11747 4675
rect 13277 4641 13311 4675
rect 16304 4641 16338 4675
rect 18245 4641 18279 4675
rect 19533 4641 19567 4675
rect 20913 4641 20947 4675
rect 22017 4641 22051 4675
rect 1777 4573 1811 4607
rect 4353 4573 4387 4607
rect 5549 4573 5583 4607
rect 8493 4573 8527 4607
rect 8677 4573 8711 4607
rect 10149 4573 10183 4607
rect 10241 4573 10275 4607
rect 11897 4573 11931 4607
rect 13369 4573 13403 4607
rect 16037 4573 16071 4607
rect 18521 4573 18555 4607
rect 19809 4573 19843 4607
rect 4721 4505 4755 4539
rect 9689 4505 9723 4539
rect 11069 4505 11103 4539
rect 1685 4437 1719 4471
rect 5181 4437 5215 4471
rect 7205 4437 7239 4471
rect 7573 4437 7607 4471
rect 9413 4437 9447 4471
rect 10793 4437 10827 4471
rect 11253 4437 11287 4471
rect 12449 4437 12483 4471
rect 14841 4437 14875 4471
rect 15485 4437 15519 4471
rect 15853 4437 15887 4471
rect 21097 4437 21131 4471
rect 22201 4437 22235 4471
rect 1593 4233 1627 4267
rect 2605 4233 2639 4267
rect 3065 4233 3099 4267
rect 4905 4233 4939 4267
rect 7941 4233 7975 4267
rect 8493 4233 8527 4267
rect 17693 4233 17727 4267
rect 17785 4233 17819 4267
rect 19073 4233 19107 4267
rect 19533 4233 19567 4267
rect 20821 4233 20855 4267
rect 2053 4097 2087 4131
rect 2237 4097 2271 4131
rect 6653 4097 6687 4131
rect 7297 4097 7331 4131
rect 7389 4097 7423 4131
rect 9137 4097 9171 4131
rect 10149 4097 10183 4131
rect 13093 4097 13127 4131
rect 13829 4097 13863 4131
rect 17417 4097 17451 4131
rect 18613 4097 18647 4131
rect 19901 4097 19935 4131
rect 22569 4097 22603 4131
rect 3157 4029 3191 4063
rect 6009 4029 6043 4063
rect 7205 4029 7239 4063
rect 8861 4029 8895 4063
rect 10416 4029 10450 4063
rect 12173 4029 12207 4063
rect 12817 4029 12851 4063
rect 14105 4029 14139 4063
rect 14841 4029 14875 4063
rect 15393 4029 15427 4063
rect 17693 4029 17727 4063
rect 18521 4029 18555 4063
rect 19625 4029 19659 4063
rect 20361 4029 20395 4063
rect 20913 4029 20947 4063
rect 21465 4029 21499 4063
rect 22017 4029 22051 4063
rect 1961 3961 1995 3995
rect 3402 3961 3436 3995
rect 5181 3961 5215 3995
rect 8401 3961 8435 3995
rect 9965 3961 9999 3995
rect 11805 3961 11839 3995
rect 12909 3961 12943 3995
rect 14381 3961 14415 3995
rect 15638 3961 15672 3995
rect 17141 3961 17175 3995
rect 18429 3961 18463 3995
rect 4537 3893 4571 3927
rect 5549 3893 5583 3927
rect 6837 3893 6871 3927
rect 8953 3893 8987 3927
rect 9505 3893 9539 3927
rect 11529 3893 11563 3927
rect 12449 3893 12483 3927
rect 13461 3893 13495 3927
rect 15301 3893 15335 3927
rect 16773 3893 16807 3927
rect 18061 3893 18095 3927
rect 21097 3893 21131 3927
rect 21833 3893 21867 3927
rect 22201 3893 22235 3927
rect 1685 3689 1719 3723
rect 3157 3689 3191 3723
rect 3433 3689 3467 3723
rect 4721 3689 4755 3723
rect 5549 3689 5583 3723
rect 6745 3689 6779 3723
rect 8125 3689 8159 3723
rect 8493 3689 8527 3723
rect 9505 3689 9539 3723
rect 10701 3689 10735 3723
rect 11069 3689 11103 3723
rect 12541 3689 12575 3723
rect 12817 3689 12851 3723
rect 13185 3689 13219 3723
rect 13829 3689 13863 3723
rect 15945 3689 15979 3723
rect 16313 3689 16347 3723
rect 17509 3689 17543 3723
rect 17877 3689 17911 3723
rect 18889 3689 18923 3723
rect 5089 3621 5123 3655
rect 6653 3621 6687 3655
rect 7113 3621 7147 3655
rect 11428 3621 11462 3655
rect 16405 3621 16439 3655
rect 19349 3621 19383 3655
rect 1777 3553 1811 3587
rect 2044 3553 2078 3587
rect 5641 3553 5675 3587
rect 7205 3553 7239 3587
rect 9873 3553 9907 3587
rect 11161 3553 11195 3587
rect 13737 3553 13771 3587
rect 19073 3553 19107 3587
rect 20913 3553 20947 3587
rect 22017 3553 22051 3587
rect 23949 3553 23983 3587
rect 4169 3485 4203 3519
rect 5733 3485 5767 3519
rect 7297 3485 7331 3519
rect 8585 3485 8619 3519
rect 10149 3485 10183 3519
rect 14013 3485 14047 3519
rect 16589 3485 16623 3519
rect 17969 3485 18003 3519
rect 18153 3485 18187 3519
rect 16957 3417 16991 3451
rect 3801 3349 3835 3383
rect 5181 3349 5215 3383
rect 6285 3349 6319 3383
rect 9045 3349 9079 3383
rect 13369 3349 13403 3383
rect 14381 3349 14415 3383
rect 14749 3349 14783 3383
rect 15485 3349 15519 3383
rect 17325 3349 17359 3383
rect 18613 3349 18647 3383
rect 21097 3349 21131 3383
rect 22201 3349 22235 3383
rect 24133 3349 24167 3383
rect 1409 3145 1443 3179
rect 2421 3145 2455 3179
rect 2973 3145 3007 3179
rect 4445 3145 4479 3179
rect 5917 3145 5951 3179
rect 6653 3145 6687 3179
rect 10425 3145 10459 3179
rect 14105 3145 14139 3179
rect 14473 3145 14507 3179
rect 16681 3145 16715 3179
rect 17601 3145 17635 3179
rect 18061 3145 18095 3179
rect 19073 3145 19107 3179
rect 21373 3145 21407 3179
rect 22109 3145 22143 3179
rect 24777 3145 24811 3179
rect 9597 3077 9631 3111
rect 9965 3077 9999 3111
rect 11529 3077 11563 3111
rect 17049 3077 17083 3111
rect 1869 3009 1903 3043
rect 2053 3009 2087 3043
rect 3617 3009 3651 3043
rect 4537 3009 4571 3043
rect 7205 3009 7239 3043
rect 8125 3009 8159 3043
rect 10885 3009 10919 3043
rect 10977 3009 11011 3043
rect 12265 3009 12299 3043
rect 16405 3009 16439 3043
rect 18521 3009 18555 3043
rect 18613 3009 18647 3043
rect 19441 3009 19475 3043
rect 20545 3009 20579 3043
rect 1777 2941 1811 2975
rect 2881 2941 2915 2975
rect 3341 2941 3375 2975
rect 3433 2941 3467 2975
rect 6193 2941 6227 2975
rect 7757 2941 7791 2975
rect 8217 2941 8251 2975
rect 8484 2941 8518 2975
rect 11805 2941 11839 2975
rect 12449 2941 12483 2975
rect 12705 2941 12739 2975
rect 14657 2941 14691 2975
rect 16865 2941 16899 2975
rect 20269 2941 20303 2975
rect 21005 2941 21039 2975
rect 21557 2941 21591 2975
rect 24593 2941 24627 2975
rect 3985 2873 4019 2907
rect 4782 2873 4816 2907
rect 14902 2873 14936 2907
rect 25237 2873 25271 2907
rect 7021 2805 7055 2839
rect 10241 2805 10275 2839
rect 10793 2805 10827 2839
rect 13829 2805 13863 2839
rect 16037 2805 16071 2839
rect 18429 2805 18463 2839
rect 21741 2805 21775 2839
rect 23949 2805 23983 2839
rect 1685 2601 1719 2635
rect 2605 2601 2639 2635
rect 3249 2601 3283 2635
rect 5733 2601 5767 2635
rect 6009 2601 6043 2635
rect 8861 2601 8895 2635
rect 10517 2601 10551 2635
rect 11437 2601 11471 2635
rect 12449 2601 12483 2635
rect 14197 2601 14231 2635
rect 15301 2601 15335 2635
rect 15853 2601 15887 2635
rect 16589 2601 16623 2635
rect 17693 2601 17727 2635
rect 18153 2601 18187 2635
rect 20913 2601 20947 2635
rect 24777 2601 24811 2635
rect 3893 2533 3927 2567
rect 4598 2533 4632 2567
rect 7389 2533 7423 2567
rect 7726 2533 7760 2567
rect 10793 2533 10827 2567
rect 11345 2533 11379 2567
rect 12081 2533 12115 2567
rect 13084 2533 13118 2567
rect 15945 2533 15979 2567
rect 19901 2533 19935 2567
rect 21465 2533 21499 2567
rect 2513 2465 2547 2499
rect 4353 2465 4387 2499
rect 7481 2465 7515 2499
rect 9229 2465 9263 2499
rect 9873 2465 9907 2499
rect 12817 2465 12851 2499
rect 14473 2465 14507 2499
rect 16957 2465 16991 2499
rect 17049 2465 17083 2499
rect 18337 2465 18371 2499
rect 19073 2465 19107 2499
rect 19625 2465 19659 2499
rect 20361 2465 20395 2499
rect 21189 2465 21223 2499
rect 21925 2465 21959 2499
rect 22477 2465 22511 2499
rect 23029 2465 23063 2499
rect 2789 2397 2823 2431
rect 6377 2397 6411 2431
rect 9597 2397 9631 2431
rect 11621 2397 11655 2431
rect 14933 2397 14967 2431
rect 16037 2397 16071 2431
rect 18521 2397 18555 2431
rect 2145 2329 2179 2363
rect 10057 2329 10091 2363
rect 15485 2329 15519 2363
rect 17233 2329 17267 2363
rect 2053 2261 2087 2295
rect 10977 2261 11011 2295
rect 22661 2261 22695 2295
<< metal1 >>
rect 4062 26528 4068 26580
rect 4120 26568 4126 26580
rect 5534 26568 5540 26580
rect 4120 26540 5540 26568
rect 4120 26528 4126 26540
rect 5534 26528 5540 26540
rect 5592 26528 5598 26580
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1578 24392 1584 24404
rect 1539 24364 1584 24392
rect 1578 24352 1584 24364
rect 1636 24352 1642 24404
rect 1394 24256 1400 24268
rect 1355 24228 1400 24256
rect 1394 24216 1400 24228
rect 1452 24216 1458 24268
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1394 23808 1400 23860
rect 1452 23848 1458 23860
rect 1854 23848 1860 23860
rect 1452 23820 1860 23848
rect 1452 23808 1458 23820
rect 1854 23808 1860 23820
rect 1912 23848 1918 23860
rect 2317 23851 2375 23857
rect 2317 23848 2329 23851
rect 1912 23820 2329 23848
rect 1912 23808 1918 23820
rect 2317 23817 2329 23820
rect 2363 23817 2375 23851
rect 2682 23848 2688 23860
rect 2643 23820 2688 23848
rect 2317 23811 2375 23817
rect 2682 23808 2688 23820
rect 2740 23808 2746 23860
rect 3786 23848 3792 23860
rect 3747 23820 3792 23848
rect 3786 23808 3792 23820
rect 3844 23808 3850 23860
rect 19981 23851 20039 23857
rect 19981 23817 19993 23851
rect 20027 23848 20039 23851
rect 20990 23848 20996 23860
rect 20027 23820 20996 23848
rect 20027 23817 20039 23820
rect 19981 23811 20039 23817
rect 20990 23808 20996 23820
rect 21048 23808 21054 23860
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23613 1455 23647
rect 1397 23607 1455 23613
rect 1412 23576 1440 23607
rect 1946 23604 1952 23656
rect 2004 23644 2010 23656
rect 2501 23647 2559 23653
rect 2501 23644 2513 23647
rect 2004 23616 2513 23644
rect 2004 23604 2010 23616
rect 2501 23613 2513 23616
rect 2547 23644 2559 23647
rect 3053 23647 3111 23653
rect 3053 23644 3065 23647
rect 2547 23616 3065 23644
rect 2547 23613 2559 23616
rect 2501 23607 2559 23613
rect 3053 23613 3065 23616
rect 3099 23613 3111 23647
rect 3053 23607 3111 23613
rect 3605 23647 3663 23653
rect 3605 23613 3617 23647
rect 3651 23644 3663 23647
rect 3651 23616 4292 23644
rect 3651 23613 3663 23616
rect 3605 23607 3663 23613
rect 1412 23548 2084 23576
rect 1578 23508 1584 23520
rect 1539 23480 1584 23508
rect 1578 23468 1584 23480
rect 1636 23468 1642 23520
rect 2056 23517 2084 23548
rect 2041 23511 2099 23517
rect 2041 23477 2053 23511
rect 2087 23508 2099 23511
rect 2590 23508 2596 23520
rect 2087 23480 2596 23508
rect 2087 23477 2099 23480
rect 2041 23471 2099 23477
rect 2590 23468 2596 23480
rect 2648 23468 2654 23520
rect 4264 23517 4292 23616
rect 4249 23511 4307 23517
rect 4249 23477 4261 23511
rect 4295 23508 4307 23511
rect 4430 23508 4436 23520
rect 4295 23480 4436 23508
rect 4295 23477 4307 23480
rect 4249 23471 4307 23477
rect 4430 23468 4436 23480
rect 4488 23468 4494 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 8294 23304 8300 23316
rect 8255 23276 8300 23304
rect 8294 23264 8300 23276
rect 8352 23264 8358 23316
rect 1946 23236 1952 23248
rect 1907 23208 1952 23236
rect 1946 23196 1952 23208
rect 2004 23196 2010 23248
rect 1673 23171 1731 23177
rect 1673 23137 1685 23171
rect 1719 23168 1731 23171
rect 2866 23168 2872 23180
rect 1719 23140 2872 23168
rect 1719 23137 1731 23140
rect 1673 23131 1731 23137
rect 2866 23128 2872 23140
rect 2924 23128 2930 23180
rect 8110 23168 8116 23180
rect 8071 23140 8116 23168
rect 8110 23128 8116 23140
rect 8168 23128 8174 23180
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 4154 22720 4160 22772
rect 4212 22760 4218 22772
rect 4249 22763 4307 22769
rect 4249 22760 4261 22763
rect 4212 22732 4261 22760
rect 4212 22720 4218 22732
rect 4249 22729 4261 22732
rect 4295 22729 4307 22763
rect 7466 22760 7472 22772
rect 7427 22732 7472 22760
rect 4249 22723 4307 22729
rect 7466 22720 7472 22732
rect 7524 22720 7530 22772
rect 8110 22720 8116 22772
rect 8168 22760 8174 22772
rect 8205 22763 8263 22769
rect 8205 22760 8217 22763
rect 8168 22732 8217 22760
rect 8168 22720 8174 22732
rect 8205 22729 8217 22732
rect 8251 22760 8263 22763
rect 8251 22732 8984 22760
rect 8251 22729 8263 22732
rect 8205 22723 8263 22729
rect 1854 22624 1860 22636
rect 1815 22596 1860 22624
rect 1854 22584 1860 22596
rect 1912 22584 1918 22636
rect 8956 22633 8984 22732
rect 8941 22627 8999 22633
rect 8941 22593 8953 22627
rect 8987 22593 8999 22627
rect 8941 22587 8999 22593
rect 1673 22559 1731 22565
rect 1673 22525 1685 22559
rect 1719 22556 1731 22559
rect 1719 22528 2544 22556
rect 1719 22525 1731 22528
rect 1673 22519 1731 22525
rect 2516 22432 2544 22528
rect 2774 22516 2780 22568
rect 2832 22556 2838 22568
rect 2961 22559 3019 22565
rect 2961 22556 2973 22559
rect 2832 22528 2973 22556
rect 2832 22516 2838 22528
rect 2961 22525 2973 22528
rect 3007 22556 3019 22559
rect 3513 22559 3571 22565
rect 3513 22556 3525 22559
rect 3007 22528 3525 22556
rect 3007 22525 3019 22528
rect 2961 22519 3019 22525
rect 3513 22525 3525 22528
rect 3559 22525 3571 22559
rect 3513 22519 3571 22525
rect 4065 22559 4123 22565
rect 4065 22525 4077 22559
rect 4111 22556 4123 22559
rect 7285 22559 7343 22565
rect 4111 22528 4752 22556
rect 4111 22525 4123 22528
rect 4065 22519 4123 22525
rect 4724 22432 4752 22528
rect 7285 22525 7297 22559
rect 7331 22556 7343 22559
rect 8757 22559 8815 22565
rect 7331 22528 7972 22556
rect 7331 22525 7343 22528
rect 7285 22519 7343 22525
rect 2498 22420 2504 22432
rect 2459 22392 2504 22420
rect 2498 22380 2504 22392
rect 2556 22380 2562 22432
rect 2866 22420 2872 22432
rect 2827 22392 2872 22420
rect 2866 22380 2872 22392
rect 2924 22380 2930 22432
rect 3142 22420 3148 22432
rect 3103 22392 3148 22420
rect 3142 22380 3148 22392
rect 3200 22380 3206 22432
rect 4706 22420 4712 22432
rect 4667 22392 4712 22420
rect 4706 22380 4712 22392
rect 4764 22380 4770 22432
rect 7944 22429 7972 22528
rect 8757 22525 8769 22559
rect 8803 22525 8815 22559
rect 8757 22519 8815 22525
rect 7929 22423 7987 22429
rect 7929 22389 7941 22423
rect 7975 22420 7987 22423
rect 8110 22420 8116 22432
rect 7975 22392 8116 22420
rect 7975 22389 7987 22392
rect 7929 22383 7987 22389
rect 8110 22380 8116 22392
rect 8168 22380 8174 22432
rect 8772 22420 8800 22519
rect 9582 22420 9588 22432
rect 8772 22392 9588 22420
rect 9582 22380 9588 22392
rect 9640 22380 9646 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1397 22083 1455 22089
rect 1397 22049 1409 22083
rect 1443 22080 1455 22083
rect 2038 22080 2044 22092
rect 1443 22052 2044 22080
rect 1443 22049 1455 22052
rect 1397 22043 1455 22049
rect 2038 22040 2044 22052
rect 2096 22040 2102 22092
rect 2498 22080 2504 22092
rect 2459 22052 2504 22080
rect 2498 22040 2504 22052
rect 2556 22040 2562 22092
rect 4062 22080 4068 22092
rect 4023 22052 4068 22080
rect 4062 22040 4068 22052
rect 4120 22040 4126 22092
rect 5445 22083 5503 22089
rect 5445 22049 5457 22083
rect 5491 22080 5503 22083
rect 5994 22080 6000 22092
rect 5491 22052 6000 22080
rect 5491 22049 5503 22052
rect 5445 22043 5503 22049
rect 5994 22040 6000 22052
rect 6052 22040 6058 22092
rect 7834 22040 7840 22092
rect 7892 22080 7898 22092
rect 8113 22083 8171 22089
rect 8113 22080 8125 22083
rect 7892 22052 8125 22080
rect 7892 22040 7898 22052
rect 8113 22049 8125 22052
rect 8159 22049 8171 22083
rect 8113 22043 8171 22049
rect 1949 22015 2007 22021
rect 1949 21981 1961 22015
rect 1995 22012 2007 22015
rect 2130 22012 2136 22024
rect 1995 21984 2136 22012
rect 1995 21981 2007 21984
rect 1949 21975 2007 21981
rect 2130 21972 2136 21984
rect 2188 21972 2194 22024
rect 8294 22012 8300 22024
rect 8255 21984 8300 22012
rect 8294 21972 8300 21984
rect 8352 21972 8358 22024
rect 1581 21947 1639 21953
rect 1581 21913 1593 21947
rect 1627 21944 1639 21947
rect 2222 21944 2228 21956
rect 1627 21916 2228 21944
rect 1627 21913 1639 21916
rect 1581 21907 1639 21913
rect 2222 21904 2228 21916
rect 2280 21904 2286 21956
rect 4246 21944 4252 21956
rect 4207 21916 4252 21944
rect 4246 21904 4252 21916
rect 4304 21904 4310 21956
rect 5534 21904 5540 21956
rect 5592 21944 5598 21956
rect 5629 21947 5687 21953
rect 5629 21944 5641 21947
rect 5592 21916 5641 21944
rect 5592 21904 5598 21916
rect 5629 21913 5641 21916
rect 5675 21913 5687 21947
rect 5629 21907 5687 21913
rect 2038 21836 2044 21888
rect 2096 21876 2102 21888
rect 2317 21879 2375 21885
rect 2317 21876 2329 21879
rect 2096 21848 2329 21876
rect 2096 21836 2102 21848
rect 2317 21845 2329 21848
rect 2363 21845 2375 21879
rect 2317 21839 2375 21845
rect 2685 21879 2743 21885
rect 2685 21845 2697 21879
rect 2731 21876 2743 21879
rect 2866 21876 2872 21888
rect 2731 21848 2872 21876
rect 2731 21845 2743 21848
rect 2685 21839 2743 21845
rect 2866 21836 2872 21848
rect 2924 21836 2930 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 4062 21632 4068 21684
rect 4120 21672 4126 21684
rect 4522 21672 4528 21684
rect 4120 21644 4528 21672
rect 4120 21632 4126 21644
rect 4522 21632 4528 21644
rect 4580 21672 4586 21684
rect 4893 21675 4951 21681
rect 4893 21672 4905 21675
rect 4580 21644 4905 21672
rect 4580 21632 4586 21644
rect 4893 21641 4905 21644
rect 4939 21641 4951 21675
rect 5258 21672 5264 21684
rect 5219 21644 5264 21672
rect 4893 21635 4951 21641
rect 5258 21632 5264 21644
rect 5316 21632 5322 21684
rect 5994 21672 6000 21684
rect 5955 21644 6000 21672
rect 5994 21632 6000 21644
rect 6052 21632 6058 21684
rect 1857 21539 1915 21545
rect 1857 21505 1869 21539
rect 1903 21536 1915 21539
rect 2682 21536 2688 21548
rect 1903 21508 2688 21536
rect 1903 21505 1915 21508
rect 1857 21499 1915 21505
rect 2682 21496 2688 21508
rect 2740 21496 2746 21548
rect 8110 21536 8116 21548
rect 8071 21508 8116 21536
rect 8110 21496 8116 21508
rect 8168 21496 8174 21548
rect 1581 21471 1639 21477
rect 1581 21437 1593 21471
rect 1627 21468 1639 21471
rect 2130 21468 2136 21480
rect 1627 21440 2136 21468
rect 1627 21437 1639 21440
rect 1581 21431 1639 21437
rect 2130 21428 2136 21440
rect 2188 21428 2194 21480
rect 2774 21428 2780 21480
rect 2832 21468 2838 21480
rect 2869 21471 2927 21477
rect 2869 21468 2881 21471
rect 2832 21440 2881 21468
rect 2832 21428 2838 21440
rect 2869 21437 2881 21440
rect 2915 21468 2927 21471
rect 3421 21471 3479 21477
rect 3421 21468 3433 21471
rect 2915 21440 3433 21468
rect 2915 21437 2927 21440
rect 2869 21431 2927 21437
rect 3421 21437 3433 21440
rect 3467 21437 3479 21471
rect 3970 21468 3976 21480
rect 3931 21440 3976 21468
rect 3421 21431 3479 21437
rect 3970 21428 3976 21440
rect 4028 21468 4034 21480
rect 4525 21471 4583 21477
rect 4525 21468 4537 21471
rect 4028 21440 4537 21468
rect 4028 21428 4034 21440
rect 4525 21437 4537 21440
rect 4571 21437 4583 21471
rect 5074 21468 5080 21480
rect 5035 21440 5080 21468
rect 4525 21431 4583 21437
rect 5074 21428 5080 21440
rect 5132 21468 5138 21480
rect 5629 21471 5687 21477
rect 5629 21468 5641 21471
rect 5132 21440 5641 21468
rect 5132 21428 5138 21440
rect 5629 21437 5641 21440
rect 5675 21437 5687 21471
rect 7926 21468 7932 21480
rect 7887 21440 7932 21468
rect 5629 21431 5687 21437
rect 7926 21428 7932 21440
rect 7984 21468 7990 21480
rect 8665 21471 8723 21477
rect 8665 21468 8677 21471
rect 7984 21440 8677 21468
rect 7984 21428 7990 21440
rect 8665 21437 8677 21440
rect 8711 21437 8723 21471
rect 8665 21431 8723 21437
rect 2498 21332 2504 21344
rect 2459 21304 2504 21332
rect 2498 21292 2504 21304
rect 2556 21292 2562 21344
rect 3050 21332 3056 21344
rect 3011 21304 3056 21332
rect 3050 21292 3056 21304
rect 3108 21292 3114 21344
rect 4154 21332 4160 21344
rect 4115 21304 4160 21332
rect 4154 21292 4160 21304
rect 4212 21292 4218 21344
rect 7834 21332 7840 21344
rect 7795 21304 7840 21332
rect 7834 21292 7840 21304
rect 7892 21292 7898 21344
rect 9217 21335 9275 21341
rect 9217 21301 9229 21335
rect 9263 21332 9275 21335
rect 10042 21332 10048 21344
rect 9263 21304 10048 21332
rect 9263 21301 9275 21304
rect 9217 21295 9275 21301
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 9674 21128 9680 21140
rect 9635 21100 9680 21128
rect 9674 21088 9680 21100
rect 9732 21088 9738 21140
rect 10042 21128 10048 21140
rect 10003 21100 10048 21128
rect 10042 21088 10048 21100
rect 10100 21088 10106 21140
rect 1946 21060 1952 21072
rect 1907 21032 1952 21060
rect 1946 21020 1952 21032
rect 2004 21020 2010 21072
rect 4430 21060 4436 21072
rect 4391 21032 4436 21060
rect 4430 21020 4436 21032
rect 4488 21020 4494 21072
rect 5994 21020 6000 21072
rect 6052 21060 6058 21072
rect 6365 21063 6423 21069
rect 6365 21060 6377 21063
rect 6052 21032 6377 21060
rect 6052 21020 6058 21032
rect 6365 21029 6377 21032
rect 6411 21029 6423 21063
rect 6365 21023 6423 21029
rect 1670 20992 1676 21004
rect 1631 20964 1676 20992
rect 1670 20952 1676 20964
rect 1728 20952 1734 21004
rect 4157 20995 4215 21001
rect 4157 20961 4169 20995
rect 4203 20992 4215 20995
rect 4246 20992 4252 21004
rect 4203 20964 4252 20992
rect 4203 20961 4215 20964
rect 4157 20955 4215 20961
rect 4246 20952 4252 20964
rect 4304 20952 4310 21004
rect 6086 20992 6092 21004
rect 6047 20964 6092 20992
rect 6086 20952 6092 20964
rect 6144 20952 6150 21004
rect 7190 20884 7196 20936
rect 7248 20924 7254 20936
rect 7377 20927 7435 20933
rect 7377 20924 7389 20927
rect 7248 20896 7389 20924
rect 7248 20884 7254 20896
rect 7377 20893 7389 20896
rect 7423 20893 7435 20927
rect 10134 20924 10140 20936
rect 10095 20896 10140 20924
rect 7377 20887 7435 20893
rect 10134 20884 10140 20896
rect 10192 20884 10198 20936
rect 10321 20927 10379 20933
rect 10321 20893 10333 20927
rect 10367 20924 10379 20927
rect 10686 20924 10692 20936
rect 10367 20896 10692 20924
rect 10367 20893 10379 20896
rect 10321 20887 10379 20893
rect 10686 20884 10692 20896
rect 10744 20884 10750 20936
rect 6914 20788 6920 20800
rect 6875 20760 6920 20788
rect 6914 20748 6920 20760
rect 6972 20748 6978 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 10042 20584 10048 20596
rect 10003 20556 10048 20584
rect 10042 20544 10048 20556
rect 10100 20544 10106 20596
rect 10134 20544 10140 20596
rect 10192 20584 10198 20596
rect 10413 20587 10471 20593
rect 10413 20584 10425 20587
rect 10192 20556 10425 20584
rect 10192 20544 10198 20556
rect 10413 20553 10425 20556
rect 10459 20553 10471 20587
rect 10413 20547 10471 20553
rect 9769 20519 9827 20525
rect 9769 20485 9781 20519
rect 9815 20516 9827 20519
rect 10686 20516 10692 20528
rect 9815 20488 10692 20516
rect 9815 20485 9827 20488
rect 9769 20479 9827 20485
rect 10686 20476 10692 20488
rect 10744 20476 10750 20528
rect 1946 20448 1952 20460
rect 1907 20420 1952 20448
rect 1946 20408 1952 20420
rect 2004 20408 2010 20460
rect 2590 20408 2596 20460
rect 2648 20448 2654 20460
rect 3145 20451 3203 20457
rect 3145 20448 3157 20451
rect 2648 20420 3157 20448
rect 2648 20408 2654 20420
rect 3145 20417 3157 20420
rect 3191 20417 3203 20451
rect 4522 20448 4528 20460
rect 4483 20420 4528 20448
rect 3145 20411 3203 20417
rect 4522 20408 4528 20420
rect 4580 20408 4586 20460
rect 1673 20383 1731 20389
rect 1673 20349 1685 20383
rect 1719 20380 1731 20383
rect 1762 20380 1768 20392
rect 1719 20352 1768 20380
rect 1719 20349 1731 20352
rect 1673 20343 1731 20349
rect 1762 20340 1768 20352
rect 1820 20380 1826 20392
rect 2409 20383 2467 20389
rect 2409 20380 2421 20383
rect 1820 20352 2421 20380
rect 1820 20340 1826 20352
rect 2409 20349 2421 20352
rect 2455 20349 2467 20383
rect 2409 20343 2467 20349
rect 2961 20383 3019 20389
rect 2961 20349 2973 20383
rect 3007 20380 3019 20383
rect 4249 20383 4307 20389
rect 3007 20352 3648 20380
rect 3007 20349 3019 20352
rect 2961 20343 3019 20349
rect 2314 20272 2320 20324
rect 2372 20312 2378 20324
rect 2777 20315 2835 20321
rect 2777 20312 2789 20315
rect 2372 20284 2789 20312
rect 2372 20272 2378 20284
rect 2777 20281 2789 20284
rect 2823 20281 2835 20315
rect 2777 20275 2835 20281
rect 3620 20256 3648 20352
rect 4249 20349 4261 20383
rect 4295 20380 4307 20383
rect 5534 20380 5540 20392
rect 4295 20352 5120 20380
rect 5495 20352 5540 20380
rect 4295 20349 4307 20352
rect 4249 20343 4307 20349
rect 5092 20256 5120 20352
rect 5534 20340 5540 20352
rect 5592 20380 5598 20392
rect 6089 20383 6147 20389
rect 6089 20380 6101 20383
rect 5592 20352 6101 20380
rect 5592 20340 5598 20352
rect 6089 20349 6101 20352
rect 6135 20349 6147 20383
rect 6089 20343 6147 20349
rect 6825 20383 6883 20389
rect 6825 20349 6837 20383
rect 6871 20380 6883 20383
rect 6914 20380 6920 20392
rect 6871 20352 6920 20380
rect 6871 20349 6883 20352
rect 6825 20343 6883 20349
rect 6914 20340 6920 20352
rect 6972 20380 6978 20392
rect 7374 20380 7380 20392
rect 6972 20352 7380 20380
rect 6972 20340 6978 20352
rect 7374 20340 7380 20352
rect 7432 20340 7438 20392
rect 5442 20272 5448 20324
rect 5500 20312 5506 20324
rect 6549 20315 6607 20321
rect 6549 20312 6561 20315
rect 5500 20284 6561 20312
rect 5500 20272 5506 20284
rect 6549 20281 6561 20284
rect 6595 20312 6607 20315
rect 7070 20315 7128 20321
rect 7070 20312 7082 20315
rect 6595 20284 7082 20312
rect 6595 20281 6607 20284
rect 6549 20275 6607 20281
rect 7070 20281 7082 20284
rect 7116 20281 7128 20315
rect 7070 20275 7128 20281
rect 2406 20204 2412 20256
rect 2464 20244 2470 20256
rect 2590 20244 2596 20256
rect 2464 20216 2596 20244
rect 2464 20204 2470 20216
rect 2590 20204 2596 20216
rect 2648 20204 2654 20256
rect 3602 20204 3608 20256
rect 3660 20244 3666 20256
rect 3697 20247 3755 20253
rect 3697 20244 3709 20247
rect 3660 20216 3709 20244
rect 3660 20204 3666 20216
rect 3697 20213 3709 20216
rect 3743 20213 3755 20247
rect 4154 20244 4160 20256
rect 4115 20216 4160 20244
rect 3697 20207 3755 20213
rect 4154 20204 4160 20216
rect 4212 20204 4218 20256
rect 5074 20244 5080 20256
rect 5035 20216 5080 20244
rect 5074 20204 5080 20216
rect 5132 20204 5138 20256
rect 5350 20244 5356 20256
rect 5311 20216 5356 20244
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 5718 20244 5724 20256
rect 5679 20216 5724 20244
rect 5718 20204 5724 20216
rect 5776 20204 5782 20256
rect 8202 20244 8208 20256
rect 8163 20216 8208 20244
rect 8202 20204 8208 20216
rect 8260 20204 8266 20256
rect 8573 20247 8631 20253
rect 8573 20213 8585 20247
rect 8619 20244 8631 20247
rect 9306 20244 9312 20256
rect 8619 20216 9312 20244
rect 8619 20213 8631 20216
rect 8573 20207 8631 20213
rect 9306 20204 9312 20216
rect 9364 20204 9370 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 2682 20040 2688 20052
rect 1688 20012 2688 20040
rect 1688 19981 1716 20012
rect 2682 20000 2688 20012
rect 2740 20000 2746 20052
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 4893 20043 4951 20049
rect 4893 20040 4905 20043
rect 4212 20012 4905 20040
rect 4212 20000 4218 20012
rect 4893 20009 4905 20012
rect 4939 20009 4951 20043
rect 4893 20003 4951 20009
rect 6086 20000 6092 20052
rect 6144 20040 6150 20052
rect 6273 20043 6331 20049
rect 6273 20040 6285 20043
rect 6144 20012 6285 20040
rect 6144 20000 6150 20012
rect 6273 20009 6285 20012
rect 6319 20009 6331 20043
rect 6273 20003 6331 20009
rect 10686 20000 10692 20052
rect 10744 20040 10750 20052
rect 11057 20043 11115 20049
rect 11057 20040 11069 20043
rect 10744 20012 11069 20040
rect 10744 20000 10750 20012
rect 11057 20009 11069 20012
rect 11103 20009 11115 20043
rect 11057 20003 11115 20009
rect 1673 19975 1731 19981
rect 1673 19941 1685 19975
rect 1719 19941 1731 19975
rect 1673 19935 1731 19941
rect 2961 19975 3019 19981
rect 2961 19941 2973 19975
rect 3007 19972 3019 19975
rect 3970 19972 3976 19984
rect 3007 19944 3976 19972
rect 3007 19941 3019 19944
rect 2961 19935 3019 19941
rect 3970 19932 3976 19944
rect 4028 19932 4034 19984
rect 4617 19975 4675 19981
rect 4617 19941 4629 19975
rect 4663 19972 4675 19975
rect 5074 19972 5080 19984
rect 4663 19944 5080 19972
rect 4663 19941 4675 19944
rect 4617 19935 4675 19941
rect 1394 19904 1400 19916
rect 1355 19876 1400 19904
rect 1394 19864 1400 19876
rect 1452 19864 1458 19916
rect 2682 19904 2688 19916
rect 2643 19876 2688 19904
rect 2682 19864 2688 19876
rect 2740 19864 2746 19916
rect 3881 19907 3939 19913
rect 3881 19873 3893 19907
rect 3927 19904 3939 19907
rect 4632 19904 4660 19935
rect 5074 19932 5080 19944
rect 5132 19972 5138 19984
rect 5350 19972 5356 19984
rect 5132 19944 5356 19972
rect 5132 19932 5138 19944
rect 5350 19932 5356 19944
rect 5408 19932 5414 19984
rect 9858 19932 9864 19984
rect 9916 19981 9922 19984
rect 9916 19975 9980 19981
rect 9916 19941 9934 19975
rect 9968 19941 9980 19975
rect 9916 19935 9980 19941
rect 9916 19932 9922 19935
rect 3927 19876 4660 19904
rect 3927 19873 3939 19876
rect 3881 19867 3939 19873
rect 4706 19864 4712 19916
rect 4764 19904 4770 19916
rect 5261 19907 5319 19913
rect 5261 19904 5273 19907
rect 4764 19876 5273 19904
rect 4764 19864 4770 19876
rect 5261 19873 5273 19876
rect 5307 19873 5319 19907
rect 5261 19867 5319 19873
rect 7644 19907 7702 19913
rect 7644 19873 7656 19907
rect 7690 19904 7702 19907
rect 8202 19904 8208 19916
rect 7690 19876 8208 19904
rect 7690 19873 7702 19876
rect 7644 19867 7702 19873
rect 8202 19864 8208 19876
rect 8260 19864 8266 19916
rect 5350 19836 5356 19848
rect 5311 19808 5356 19836
rect 5350 19796 5356 19808
rect 5408 19796 5414 19848
rect 5442 19796 5448 19848
rect 5500 19836 5506 19848
rect 7374 19836 7380 19848
rect 5500 19808 5545 19836
rect 7287 19808 7380 19836
rect 5500 19796 5506 19808
rect 7374 19796 7380 19808
rect 7432 19796 7438 19848
rect 9677 19839 9735 19845
rect 9677 19836 9689 19839
rect 9416 19808 9689 19836
rect 1670 19660 1676 19712
rect 1728 19700 1734 19712
rect 2130 19700 2136 19712
rect 1728 19672 2136 19700
rect 1728 19660 1734 19672
rect 2130 19660 2136 19672
rect 2188 19660 2194 19712
rect 2406 19660 2412 19712
rect 2464 19700 2470 19712
rect 2501 19703 2559 19709
rect 2501 19700 2513 19703
rect 2464 19672 2513 19700
rect 2464 19660 2470 19672
rect 2501 19669 2513 19672
rect 2547 19669 2559 19703
rect 3510 19700 3516 19712
rect 3471 19672 3516 19700
rect 2501 19663 2559 19669
rect 3510 19660 3516 19672
rect 3568 19660 3574 19712
rect 4154 19660 4160 19712
rect 4212 19700 4218 19712
rect 4249 19703 4307 19709
rect 4249 19700 4261 19703
rect 4212 19672 4261 19700
rect 4212 19660 4218 19672
rect 4249 19669 4261 19672
rect 4295 19669 4307 19703
rect 5994 19700 6000 19712
rect 5955 19672 6000 19700
rect 4249 19663 4307 19669
rect 5994 19660 6000 19672
rect 6052 19660 6058 19712
rect 6914 19700 6920 19712
rect 6875 19672 6920 19700
rect 6914 19660 6920 19672
rect 6972 19660 6978 19712
rect 7282 19700 7288 19712
rect 7243 19672 7288 19700
rect 7282 19660 7288 19672
rect 7340 19660 7346 19712
rect 7392 19700 7420 19796
rect 8312 19740 9076 19768
rect 8312 19700 8340 19740
rect 9048 19712 9076 19740
rect 7392 19672 8340 19700
rect 8662 19660 8668 19712
rect 8720 19700 8726 19712
rect 8757 19703 8815 19709
rect 8757 19700 8769 19703
rect 8720 19672 8769 19700
rect 8720 19660 8726 19672
rect 8757 19669 8769 19672
rect 8803 19669 8815 19703
rect 9030 19700 9036 19712
rect 8991 19672 9036 19700
rect 8757 19663 8815 19669
rect 9030 19660 9036 19672
rect 9088 19660 9094 19712
rect 9306 19660 9312 19712
rect 9364 19700 9370 19712
rect 9416 19709 9444 19808
rect 9677 19805 9689 19808
rect 9723 19805 9735 19839
rect 9677 19799 9735 19805
rect 9401 19703 9459 19709
rect 9401 19700 9413 19703
rect 9364 19672 9413 19700
rect 9364 19660 9370 19672
rect 9401 19669 9413 19672
rect 9447 19669 9459 19703
rect 9401 19663 9459 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1394 19456 1400 19508
rect 1452 19496 1458 19508
rect 2317 19499 2375 19505
rect 2317 19496 2329 19499
rect 1452 19468 2329 19496
rect 1452 19456 1458 19468
rect 2317 19465 2329 19468
rect 2363 19465 2375 19499
rect 4706 19496 4712 19508
rect 4667 19468 4712 19496
rect 2317 19459 2375 19465
rect 4706 19456 4712 19468
rect 4764 19456 4770 19508
rect 5166 19496 5172 19508
rect 5127 19468 5172 19496
rect 5166 19456 5172 19468
rect 5224 19456 5230 19508
rect 6086 19456 6092 19508
rect 6144 19496 6150 19508
rect 6825 19499 6883 19505
rect 6825 19496 6837 19499
rect 6144 19468 6837 19496
rect 6144 19456 6150 19468
rect 6825 19465 6837 19468
rect 6871 19465 6883 19499
rect 6825 19459 6883 19465
rect 10134 19456 10140 19508
rect 10192 19496 10198 19508
rect 10597 19499 10655 19505
rect 10597 19496 10609 19499
rect 10192 19468 10609 19496
rect 10192 19456 10198 19468
rect 10597 19465 10609 19468
rect 10643 19465 10655 19499
rect 10597 19459 10655 19465
rect 1486 19320 1492 19372
rect 1544 19360 1550 19372
rect 2682 19360 2688 19372
rect 1544 19332 2688 19360
rect 1544 19320 1550 19332
rect 2682 19320 2688 19332
rect 2740 19320 2746 19372
rect 4157 19363 4215 19369
rect 4157 19329 4169 19363
rect 4203 19360 4215 19363
rect 4724 19360 4752 19456
rect 5994 19428 6000 19440
rect 5644 19400 6000 19428
rect 5644 19369 5672 19400
rect 5994 19388 6000 19400
rect 6052 19428 6058 19440
rect 6730 19428 6736 19440
rect 6052 19400 6736 19428
rect 6052 19388 6058 19400
rect 6730 19388 6736 19400
rect 6788 19388 6794 19440
rect 6914 19388 6920 19440
rect 6972 19428 6978 19440
rect 8205 19431 8263 19437
rect 8205 19428 8217 19431
rect 6972 19400 8217 19428
rect 6972 19388 6978 19400
rect 4203 19332 4752 19360
rect 5629 19363 5687 19369
rect 4203 19329 4215 19332
rect 4157 19323 4215 19329
rect 5629 19329 5641 19363
rect 5675 19329 5687 19363
rect 5629 19323 5687 19329
rect 5813 19363 5871 19369
rect 5813 19329 5825 19363
rect 5859 19360 5871 19363
rect 6181 19363 6239 19369
rect 6181 19360 6193 19363
rect 5859 19332 6193 19360
rect 5859 19329 5871 19332
rect 5813 19323 5871 19329
rect 6181 19329 6193 19332
rect 6227 19360 6239 19363
rect 6822 19360 6828 19372
rect 6227 19332 6828 19360
rect 6227 19329 6239 19332
rect 6181 19323 6239 19329
rect 6822 19320 6828 19332
rect 6880 19320 6886 19372
rect 7282 19360 7288 19372
rect 7243 19332 7288 19360
rect 7282 19320 7288 19332
rect 7340 19320 7346 19372
rect 7392 19369 7420 19400
rect 8205 19397 8217 19400
rect 8251 19397 8263 19431
rect 8205 19391 8263 19397
rect 7377 19363 7435 19369
rect 7377 19329 7389 19363
rect 7423 19329 7435 19363
rect 8220 19360 8248 19391
rect 8220 19332 8524 19360
rect 7377 19323 7435 19329
rect 1578 19292 1584 19304
rect 1539 19264 1584 19292
rect 1578 19252 1584 19264
rect 1636 19252 1642 19304
rect 1857 19295 1915 19301
rect 1857 19261 1869 19295
rect 1903 19292 1915 19295
rect 2038 19292 2044 19304
rect 1903 19264 2044 19292
rect 1903 19261 1915 19264
rect 1857 19255 1915 19261
rect 2038 19252 2044 19264
rect 2096 19252 2102 19304
rect 2866 19292 2872 19304
rect 2779 19264 2872 19292
rect 2866 19252 2872 19264
rect 2924 19292 2930 19304
rect 3605 19295 3663 19301
rect 3605 19292 3617 19295
rect 2924 19264 3617 19292
rect 2924 19252 2930 19264
rect 3605 19261 3617 19264
rect 3651 19261 3663 19295
rect 3605 19255 3663 19261
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19292 6699 19295
rect 7190 19292 7196 19304
rect 6687 19264 7196 19292
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 7190 19252 7196 19264
rect 7248 19252 7254 19304
rect 8389 19295 8447 19301
rect 8389 19261 8401 19295
rect 8435 19261 8447 19295
rect 8496 19292 8524 19332
rect 9858 19320 9864 19372
rect 9916 19360 9922 19372
rect 11149 19363 11207 19369
rect 11149 19360 11161 19363
rect 9916 19332 11161 19360
rect 9916 19320 9922 19332
rect 11149 19329 11161 19332
rect 11195 19329 11207 19363
rect 11149 19323 11207 19329
rect 8662 19301 8668 19304
rect 8645 19295 8668 19301
rect 8645 19292 8657 19295
rect 8496 19264 8657 19292
rect 8389 19255 8447 19261
rect 8645 19261 8657 19264
rect 8720 19292 8726 19304
rect 10505 19295 10563 19301
rect 8720 19264 8793 19292
rect 8645 19255 8668 19261
rect 2498 19184 2504 19236
rect 2556 19224 2562 19236
rect 3145 19227 3203 19233
rect 3145 19224 3157 19227
rect 2556 19196 3157 19224
rect 2556 19184 2562 19196
rect 3145 19193 3157 19196
rect 3191 19193 3203 19227
rect 3145 19187 3203 19193
rect 4065 19227 4123 19233
rect 4065 19193 4077 19227
rect 4111 19224 4123 19227
rect 5350 19224 5356 19236
rect 4111 19196 5356 19224
rect 4111 19193 4123 19196
rect 4065 19187 4123 19193
rect 5350 19184 5356 19196
rect 5408 19184 5414 19236
rect 8404 19224 8432 19255
rect 8662 19252 8668 19255
rect 8720 19252 8726 19264
rect 10505 19261 10517 19295
rect 10551 19292 10563 19295
rect 10962 19292 10968 19304
rect 10551 19264 10968 19292
rect 10551 19261 10563 19264
rect 10505 19255 10563 19261
rect 10962 19252 10968 19264
rect 11020 19292 11026 19304
rect 11057 19295 11115 19301
rect 11057 19292 11069 19295
rect 11020 19264 11069 19292
rect 11020 19252 11026 19264
rect 11057 19261 11069 19264
rect 11103 19261 11115 19295
rect 11057 19255 11115 19261
rect 9306 19224 9312 19236
rect 8404 19196 9312 19224
rect 9306 19184 9312 19196
rect 9364 19184 9370 19236
rect 2130 19116 2136 19168
rect 2188 19156 2194 19168
rect 2590 19156 2596 19168
rect 2188 19128 2596 19156
rect 2188 19116 2194 19128
rect 2590 19116 2596 19128
rect 2648 19116 2654 19168
rect 5077 19159 5135 19165
rect 5077 19125 5089 19159
rect 5123 19156 5135 19159
rect 5537 19159 5595 19165
rect 5537 19156 5549 19159
rect 5123 19128 5549 19156
rect 5123 19125 5135 19128
rect 5077 19119 5135 19125
rect 5537 19125 5549 19128
rect 5583 19156 5595 19159
rect 5626 19156 5632 19168
rect 5583 19128 5632 19156
rect 5583 19125 5595 19128
rect 5537 19119 5595 19125
rect 5626 19116 5632 19128
rect 5684 19116 5690 19168
rect 7929 19159 7987 19165
rect 7929 19125 7941 19159
rect 7975 19156 7987 19159
rect 8202 19156 8208 19168
rect 7975 19128 8208 19156
rect 7975 19125 7987 19128
rect 7929 19119 7987 19125
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 9490 19116 9496 19168
rect 9548 19156 9554 19168
rect 9769 19159 9827 19165
rect 9769 19156 9781 19159
rect 9548 19128 9781 19156
rect 9548 19116 9554 19128
rect 9769 19125 9781 19128
rect 9815 19156 9827 19159
rect 9858 19156 9864 19168
rect 9815 19128 9864 19156
rect 9815 19125 9827 19128
rect 9769 19119 9827 19125
rect 9858 19116 9864 19128
rect 9916 19116 9922 19168
rect 10042 19116 10048 19168
rect 10100 19156 10106 19168
rect 10137 19159 10195 19165
rect 10137 19156 10149 19159
rect 10100 19128 10149 19156
rect 10100 19116 10106 19128
rect 10137 19125 10149 19128
rect 10183 19156 10195 19159
rect 10965 19159 11023 19165
rect 10965 19156 10977 19159
rect 10183 19128 10977 19156
rect 10183 19125 10195 19128
rect 10137 19119 10195 19125
rect 10965 19125 10977 19128
rect 11011 19156 11023 19159
rect 12802 19156 12808 19168
rect 11011 19128 12808 19156
rect 11011 19125 11023 19128
rect 10965 19119 11023 19125
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 4985 18955 5043 18961
rect 4985 18921 4997 18955
rect 5031 18952 5043 18955
rect 5442 18952 5448 18964
rect 5031 18924 5448 18952
rect 5031 18921 5043 18924
rect 4985 18915 5043 18921
rect 5442 18912 5448 18924
rect 5500 18952 5506 18964
rect 6641 18955 6699 18961
rect 6641 18952 6653 18955
rect 5500 18924 6653 18952
rect 5500 18912 5506 18924
rect 6641 18921 6653 18924
rect 6687 18921 6699 18955
rect 6641 18915 6699 18921
rect 7282 18912 7288 18964
rect 7340 18952 7346 18964
rect 7469 18955 7527 18961
rect 7469 18952 7481 18955
rect 7340 18924 7481 18952
rect 7340 18912 7346 18924
rect 7469 18921 7481 18924
rect 7515 18921 7527 18955
rect 9490 18952 9496 18964
rect 9451 18924 9496 18952
rect 7469 18915 7527 18921
rect 9490 18912 9496 18924
rect 9548 18912 9554 18964
rect 9677 18955 9735 18961
rect 9677 18921 9689 18955
rect 9723 18952 9735 18955
rect 9766 18952 9772 18964
rect 9723 18924 9772 18952
rect 9723 18921 9735 18924
rect 9677 18915 9735 18921
rect 9766 18912 9772 18924
rect 9824 18912 9830 18964
rect 9508 18884 9536 18912
rect 10689 18887 10747 18893
rect 10689 18884 10701 18887
rect 9508 18856 10701 18884
rect 10689 18853 10701 18856
rect 10735 18853 10747 18887
rect 10689 18847 10747 18853
rect 2038 18776 2044 18828
rect 2096 18816 2102 18828
rect 2314 18816 2320 18828
rect 2096 18788 2320 18816
rect 2096 18776 2102 18788
rect 2314 18776 2320 18788
rect 2372 18776 2378 18828
rect 4062 18816 4068 18828
rect 4023 18788 4068 18816
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 5534 18825 5540 18828
rect 5528 18816 5540 18825
rect 5495 18788 5540 18816
rect 5528 18779 5540 18788
rect 5534 18776 5540 18779
rect 5592 18776 5598 18828
rect 7374 18776 7380 18828
rect 7432 18816 7438 18828
rect 7837 18819 7895 18825
rect 7837 18816 7849 18819
rect 7432 18788 7849 18816
rect 7432 18776 7438 18788
rect 7837 18785 7849 18788
rect 7883 18785 7895 18819
rect 7837 18779 7895 18785
rect 7929 18819 7987 18825
rect 7929 18785 7941 18819
rect 7975 18816 7987 18819
rect 8386 18816 8392 18828
rect 7975 18788 8392 18816
rect 7975 18785 7987 18788
rect 7929 18779 7987 18785
rect 8386 18776 8392 18788
rect 8444 18776 8450 18828
rect 9214 18776 9220 18828
rect 9272 18816 9278 18828
rect 10045 18819 10103 18825
rect 10045 18816 10057 18819
rect 9272 18788 10057 18816
rect 9272 18776 9278 18788
rect 10045 18785 10057 18788
rect 10091 18785 10103 18819
rect 10045 18779 10103 18785
rect 2406 18748 2412 18760
rect 2367 18720 2412 18748
rect 2406 18708 2412 18720
rect 2464 18708 2470 18760
rect 2498 18708 2504 18760
rect 2556 18748 2562 18760
rect 2556 18720 2601 18748
rect 2556 18708 2562 18720
rect 5166 18708 5172 18760
rect 5224 18748 5230 18760
rect 5261 18751 5319 18757
rect 5261 18748 5273 18751
rect 5224 18720 5273 18748
rect 5224 18708 5230 18720
rect 5261 18717 5273 18720
rect 5307 18717 5319 18751
rect 5261 18711 5319 18717
rect 8113 18751 8171 18757
rect 8113 18717 8125 18751
rect 8159 18748 8171 18751
rect 8202 18748 8208 18760
rect 8159 18720 8208 18748
rect 8159 18717 8171 18720
rect 8113 18711 8171 18717
rect 8202 18708 8208 18720
rect 8260 18708 8266 18760
rect 10134 18748 10140 18760
rect 10095 18720 10140 18748
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 10318 18748 10324 18760
rect 10231 18720 10324 18748
rect 10318 18708 10324 18720
rect 10376 18748 10382 18760
rect 10962 18748 10968 18760
rect 10376 18720 10968 18748
rect 10376 18708 10382 18720
rect 10962 18708 10968 18720
rect 11020 18708 11026 18760
rect 1857 18683 1915 18689
rect 1857 18649 1869 18683
rect 1903 18680 1915 18683
rect 2516 18680 2544 18708
rect 1903 18652 2544 18680
rect 1903 18649 1915 18652
rect 1857 18643 1915 18649
rect 1946 18612 1952 18624
rect 1907 18584 1952 18612
rect 1946 18572 1952 18584
rect 2004 18572 2010 18624
rect 2958 18612 2964 18624
rect 2919 18584 2964 18612
rect 2958 18572 2964 18584
rect 3016 18572 3022 18624
rect 3694 18612 3700 18624
rect 3655 18584 3700 18612
rect 3694 18572 3700 18584
rect 3752 18572 3758 18624
rect 4246 18612 4252 18624
rect 4207 18584 4252 18612
rect 4246 18572 4252 18584
rect 4304 18572 4310 18624
rect 7285 18615 7343 18621
rect 7285 18581 7297 18615
rect 7331 18612 7343 18615
rect 7374 18612 7380 18624
rect 7331 18584 7380 18612
rect 7331 18581 7343 18584
rect 7285 18575 7343 18581
rect 7374 18572 7380 18584
rect 7432 18572 7438 18624
rect 8478 18612 8484 18624
rect 8439 18584 8484 18612
rect 8478 18572 8484 18584
rect 8536 18612 8542 18624
rect 8849 18615 8907 18621
rect 8849 18612 8861 18615
rect 8536 18584 8861 18612
rect 8536 18572 8542 18584
rect 8849 18581 8861 18584
rect 8895 18612 8907 18615
rect 9030 18612 9036 18624
rect 8895 18584 9036 18612
rect 8895 18581 8907 18584
rect 8849 18575 8907 18581
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 3602 18408 3608 18420
rect 3563 18380 3608 18408
rect 3602 18368 3608 18380
rect 3660 18368 3666 18420
rect 5169 18411 5227 18417
rect 5169 18377 5181 18411
rect 5215 18408 5227 18411
rect 5350 18408 5356 18420
rect 5215 18380 5356 18408
rect 5215 18377 5227 18380
rect 5169 18371 5227 18377
rect 5350 18368 5356 18380
rect 5408 18368 5414 18420
rect 6730 18368 6736 18420
rect 6788 18408 6794 18420
rect 7193 18411 7251 18417
rect 7193 18408 7205 18411
rect 6788 18380 7205 18408
rect 6788 18368 6794 18380
rect 7193 18377 7205 18380
rect 7239 18377 7251 18411
rect 9214 18408 9220 18420
rect 9175 18380 9220 18408
rect 7193 18371 7251 18377
rect 9214 18368 9220 18380
rect 9272 18368 9278 18420
rect 10226 18368 10232 18420
rect 10284 18408 10290 18420
rect 10965 18411 11023 18417
rect 10965 18408 10977 18411
rect 10284 18380 10977 18408
rect 10284 18368 10290 18380
rect 10965 18377 10977 18380
rect 11011 18377 11023 18411
rect 10965 18371 11023 18377
rect 10686 18340 10692 18352
rect 10647 18312 10692 18340
rect 10686 18300 10692 18312
rect 10744 18300 10750 18352
rect 2498 18232 2504 18284
rect 2556 18272 2562 18284
rect 2593 18275 2651 18281
rect 2593 18272 2605 18275
rect 2556 18244 2605 18272
rect 2556 18232 2562 18244
rect 2593 18241 2605 18244
rect 2639 18272 2651 18275
rect 2639 18244 2728 18272
rect 2639 18241 2651 18244
rect 2593 18235 2651 18241
rect 1857 18139 1915 18145
rect 1857 18105 1869 18139
rect 1903 18136 1915 18139
rect 1903 18108 2452 18136
rect 1903 18105 1915 18108
rect 1857 18099 1915 18105
rect 1949 18071 2007 18077
rect 1949 18037 1961 18071
rect 1995 18068 2007 18071
rect 2130 18068 2136 18080
rect 1995 18040 2136 18068
rect 1995 18037 2007 18040
rect 1949 18031 2007 18037
rect 2130 18028 2136 18040
rect 2188 18028 2194 18080
rect 2314 18068 2320 18080
rect 2275 18040 2320 18068
rect 2314 18028 2320 18040
rect 2372 18028 2378 18080
rect 2424 18077 2452 18108
rect 2409 18071 2467 18077
rect 2409 18037 2421 18071
rect 2455 18068 2467 18071
rect 2498 18068 2504 18080
rect 2455 18040 2504 18068
rect 2455 18037 2467 18040
rect 2409 18031 2467 18037
rect 2498 18028 2504 18040
rect 2556 18028 2562 18080
rect 2700 18068 2728 18244
rect 3694 18232 3700 18284
rect 3752 18272 3758 18284
rect 4157 18275 4215 18281
rect 4157 18272 4169 18275
rect 3752 18244 4169 18272
rect 3752 18232 3758 18244
rect 4157 18241 4169 18244
rect 4203 18241 4215 18275
rect 4157 18235 4215 18241
rect 5534 18232 5540 18284
rect 5592 18272 5598 18284
rect 5810 18272 5816 18284
rect 5592 18244 5816 18272
rect 5592 18232 5598 18244
rect 5810 18232 5816 18244
rect 5868 18272 5874 18284
rect 6270 18272 6276 18284
rect 5868 18244 6276 18272
rect 5868 18232 5874 18244
rect 6270 18232 6276 18244
rect 6328 18232 6334 18284
rect 7742 18272 7748 18284
rect 7703 18244 7748 18272
rect 7742 18232 7748 18244
rect 7800 18232 7806 18284
rect 8297 18207 8355 18213
rect 8297 18173 8309 18207
rect 8343 18204 8355 18207
rect 8386 18204 8392 18216
rect 8343 18176 8392 18204
rect 8343 18173 8355 18176
rect 8297 18167 8355 18173
rect 8386 18164 8392 18176
rect 8444 18164 8450 18216
rect 9306 18204 9312 18216
rect 9267 18176 9312 18204
rect 9306 18164 9312 18176
rect 9364 18164 9370 18216
rect 9398 18164 9404 18216
rect 9456 18204 9462 18216
rect 9576 18207 9634 18213
rect 9576 18204 9588 18207
rect 9456 18176 9588 18204
rect 9456 18164 9462 18176
rect 9576 18173 9588 18176
rect 9622 18204 9634 18207
rect 10318 18204 10324 18216
rect 9622 18176 10324 18204
rect 9622 18173 9634 18176
rect 9576 18167 9634 18173
rect 10318 18164 10324 18176
rect 10376 18164 10382 18216
rect 2774 18096 2780 18148
rect 2832 18136 2838 18148
rect 3421 18139 3479 18145
rect 3421 18136 3433 18139
rect 2832 18108 3433 18136
rect 2832 18096 2838 18108
rect 3421 18105 3433 18108
rect 3467 18136 3479 18139
rect 3973 18139 4031 18145
rect 3973 18136 3985 18139
rect 3467 18108 3985 18136
rect 3467 18105 3479 18108
rect 3421 18099 3479 18105
rect 3973 18105 3985 18108
rect 4019 18105 4031 18139
rect 3973 18099 4031 18105
rect 5077 18139 5135 18145
rect 5077 18105 5089 18139
rect 5123 18136 5135 18139
rect 6641 18139 6699 18145
rect 5123 18108 5672 18136
rect 5123 18105 5135 18108
rect 5077 18099 5135 18105
rect 2961 18071 3019 18077
rect 2961 18068 2973 18071
rect 2700 18040 2973 18068
rect 2961 18037 2973 18040
rect 3007 18068 3019 18071
rect 3326 18068 3332 18080
rect 3007 18040 3332 18068
rect 3007 18037 3019 18040
rect 2961 18031 3019 18037
rect 3326 18028 3332 18040
rect 3384 18028 3390 18080
rect 4062 18068 4068 18080
rect 4023 18040 4068 18068
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 4614 18068 4620 18080
rect 4575 18040 4620 18068
rect 4614 18028 4620 18040
rect 4672 18068 4678 18080
rect 5644 18077 5672 18108
rect 6641 18105 6653 18139
rect 6687 18136 6699 18139
rect 7374 18136 7380 18148
rect 6687 18108 7380 18136
rect 6687 18105 6699 18108
rect 6641 18099 6699 18105
rect 7374 18096 7380 18108
rect 7432 18136 7438 18148
rect 7561 18139 7619 18145
rect 7561 18136 7573 18139
rect 7432 18108 7573 18136
rect 7432 18096 7438 18108
rect 7561 18105 7573 18108
rect 7607 18105 7619 18139
rect 7561 18099 7619 18105
rect 8849 18139 8907 18145
rect 8849 18105 8861 18139
rect 8895 18136 8907 18139
rect 9416 18136 9444 18164
rect 8895 18108 9444 18136
rect 8895 18105 8907 18108
rect 8849 18099 8907 18105
rect 5537 18071 5595 18077
rect 5537 18068 5549 18071
rect 4672 18040 5549 18068
rect 4672 18028 4678 18040
rect 5537 18037 5549 18040
rect 5583 18037 5595 18071
rect 5537 18031 5595 18037
rect 5629 18071 5687 18077
rect 5629 18037 5641 18071
rect 5675 18068 5687 18071
rect 5994 18068 6000 18080
rect 5675 18040 6000 18068
rect 5675 18037 5687 18040
rect 5629 18031 5687 18037
rect 5994 18028 6000 18040
rect 6052 18028 6058 18080
rect 7101 18071 7159 18077
rect 7101 18037 7113 18071
rect 7147 18068 7159 18071
rect 7650 18068 7656 18080
rect 7147 18040 7656 18068
rect 7147 18037 7159 18040
rect 7101 18031 7159 18037
rect 7650 18028 7656 18040
rect 7708 18028 7714 18080
rect 11425 18071 11483 18077
rect 11425 18037 11437 18071
rect 11471 18068 11483 18071
rect 12066 18068 12072 18080
rect 11471 18040 12072 18068
rect 11471 18037 11483 18040
rect 11425 18031 11483 18037
rect 12066 18028 12072 18040
rect 12124 18028 12130 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1397 17867 1455 17873
rect 1397 17833 1409 17867
rect 1443 17864 1455 17867
rect 2682 17864 2688 17876
rect 1443 17836 2688 17864
rect 1443 17833 1455 17836
rect 1397 17827 1455 17833
rect 2682 17824 2688 17836
rect 2740 17824 2746 17876
rect 5810 17864 5816 17876
rect 5771 17836 5816 17864
rect 5810 17824 5816 17836
rect 5868 17824 5874 17876
rect 6086 17824 6092 17876
rect 6144 17864 6150 17876
rect 7653 17867 7711 17873
rect 7653 17864 7665 17867
rect 6144 17836 7665 17864
rect 6144 17824 6150 17836
rect 7653 17833 7665 17836
rect 7699 17833 7711 17867
rect 8294 17864 8300 17876
rect 8255 17836 8300 17864
rect 7653 17827 7711 17833
rect 8294 17824 8300 17836
rect 8352 17824 8358 17876
rect 8573 17867 8631 17873
rect 8573 17833 8585 17867
rect 8619 17864 8631 17867
rect 9214 17864 9220 17876
rect 8619 17836 9220 17864
rect 8619 17833 8631 17836
rect 8573 17827 8631 17833
rect 9214 17824 9220 17836
rect 9272 17824 9278 17876
rect 9398 17864 9404 17876
rect 9359 17836 9404 17864
rect 9398 17824 9404 17836
rect 9456 17824 9462 17876
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 11149 17867 11207 17873
rect 11149 17864 11161 17867
rect 11112 17836 11161 17864
rect 11112 17824 11118 17836
rect 11149 17833 11161 17836
rect 11195 17833 11207 17867
rect 11149 17827 11207 17833
rect 3513 17799 3571 17805
rect 3513 17765 3525 17799
rect 3559 17796 3571 17799
rect 4062 17796 4068 17808
rect 3559 17768 4068 17796
rect 3559 17765 3571 17768
rect 3513 17759 3571 17765
rect 4062 17756 4068 17768
rect 4120 17756 4126 17808
rect 2774 17688 2780 17740
rect 2832 17728 2838 17740
rect 4321 17731 4379 17737
rect 4321 17728 4333 17731
rect 2832 17700 2877 17728
rect 3804 17700 4333 17728
rect 2832 17688 2838 17700
rect 3804 17672 3832 17700
rect 4321 17697 4333 17700
rect 4367 17697 4379 17731
rect 4321 17691 4379 17697
rect 6362 17688 6368 17740
rect 6420 17728 6426 17740
rect 6529 17731 6587 17737
rect 6529 17728 6541 17731
rect 6420 17700 6541 17728
rect 6420 17688 6426 17700
rect 6529 17697 6541 17700
rect 6575 17697 6587 17731
rect 6529 17691 6587 17697
rect 9858 17688 9864 17740
rect 9916 17728 9922 17740
rect 10025 17731 10083 17737
rect 10025 17728 10037 17731
rect 9916 17700 10037 17728
rect 9916 17688 9922 17700
rect 10025 17697 10037 17700
rect 10071 17697 10083 17731
rect 10025 17691 10083 17697
rect 2866 17660 2872 17672
rect 2827 17632 2872 17660
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 2958 17620 2964 17672
rect 3016 17660 3022 17672
rect 3786 17660 3792 17672
rect 3016 17632 3792 17660
rect 3016 17620 3022 17632
rect 3786 17620 3792 17632
rect 3844 17620 3850 17672
rect 3970 17620 3976 17672
rect 4028 17660 4034 17672
rect 4065 17663 4123 17669
rect 4065 17660 4077 17663
rect 4028 17632 4077 17660
rect 4028 17620 4034 17632
rect 4065 17629 4077 17632
rect 4111 17629 4123 17663
rect 6273 17663 6331 17669
rect 6273 17660 6285 17663
rect 4065 17623 4123 17629
rect 6196 17632 6285 17660
rect 1486 17552 1492 17604
rect 1544 17592 1550 17604
rect 2409 17595 2467 17601
rect 2409 17592 2421 17595
rect 1544 17564 2421 17592
rect 1544 17552 1550 17564
rect 2409 17561 2421 17564
rect 2455 17561 2467 17595
rect 2409 17555 2467 17561
rect 6196 17536 6224 17632
rect 6273 17629 6285 17632
rect 6319 17629 6331 17663
rect 9766 17660 9772 17672
rect 9727 17632 9772 17660
rect 6273 17623 6331 17629
rect 9766 17620 9772 17632
rect 9824 17620 9830 17672
rect 7742 17592 7748 17604
rect 7208 17564 7748 17592
rect 7208 17536 7236 17564
rect 7742 17552 7748 17564
rect 7800 17592 7806 17604
rect 7929 17595 7987 17601
rect 7929 17592 7941 17595
rect 7800 17564 7941 17592
rect 7800 17552 7806 17564
rect 7929 17561 7941 17564
rect 7975 17561 7987 17595
rect 7929 17555 7987 17561
rect 1394 17484 1400 17536
rect 1452 17524 1458 17536
rect 1949 17527 2007 17533
rect 1949 17524 1961 17527
rect 1452 17496 1961 17524
rect 1452 17484 1458 17496
rect 1949 17493 1961 17496
rect 1995 17524 2007 17527
rect 2314 17524 2320 17536
rect 1995 17496 2320 17524
rect 1995 17493 2007 17496
rect 1949 17487 2007 17493
rect 2314 17484 2320 17496
rect 2372 17484 2378 17536
rect 5442 17524 5448 17536
rect 5403 17496 5448 17524
rect 5442 17484 5448 17496
rect 5500 17484 5506 17536
rect 6178 17524 6184 17536
rect 6139 17496 6184 17524
rect 6178 17484 6184 17496
rect 6236 17484 6242 17536
rect 7190 17484 7196 17536
rect 7248 17484 7254 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 4062 17280 4068 17332
rect 4120 17320 4126 17332
rect 4985 17323 5043 17329
rect 4985 17320 4997 17323
rect 4120 17292 4997 17320
rect 4120 17280 4126 17292
rect 4985 17289 4997 17292
rect 5031 17289 5043 17323
rect 4985 17283 5043 17289
rect 9677 17323 9735 17329
rect 9677 17289 9689 17323
rect 9723 17320 9735 17323
rect 9950 17320 9956 17332
rect 9723 17292 9956 17320
rect 9723 17289 9735 17292
rect 9677 17283 9735 17289
rect 9950 17280 9956 17292
rect 10008 17280 10014 17332
rect 3786 17212 3792 17264
rect 3844 17252 3850 17264
rect 4157 17255 4215 17261
rect 4157 17252 4169 17255
rect 3844 17224 4169 17252
rect 3844 17212 3850 17224
rect 4157 17221 4169 17224
rect 4203 17221 4215 17255
rect 4157 17215 4215 17221
rect 8110 17212 8116 17264
rect 8168 17252 8174 17264
rect 9306 17252 9312 17264
rect 8168 17224 9312 17252
rect 8168 17212 8174 17224
rect 9306 17212 9312 17224
rect 9364 17252 9370 17264
rect 9766 17252 9772 17264
rect 9364 17224 9772 17252
rect 9364 17212 9370 17224
rect 9766 17212 9772 17224
rect 9824 17212 9830 17264
rect 5442 17144 5448 17196
rect 5500 17184 5506 17196
rect 5537 17187 5595 17193
rect 5537 17184 5549 17187
rect 5500 17156 5549 17184
rect 5500 17144 5506 17156
rect 5537 17153 5549 17156
rect 5583 17184 5595 17187
rect 5997 17187 6055 17193
rect 5997 17184 6009 17187
rect 5583 17156 6009 17184
rect 5583 17153 5595 17156
rect 5537 17147 5595 17153
rect 5997 17153 6009 17156
rect 6043 17184 6055 17187
rect 6362 17184 6368 17196
rect 6043 17156 6368 17184
rect 6043 17153 6055 17156
rect 5997 17147 6055 17153
rect 6362 17144 6368 17156
rect 6420 17144 6426 17196
rect 10321 17187 10379 17193
rect 10321 17153 10333 17187
rect 10367 17184 10379 17187
rect 10686 17184 10692 17196
rect 10367 17156 10692 17184
rect 10367 17153 10379 17156
rect 10321 17147 10379 17153
rect 10686 17144 10692 17156
rect 10744 17144 10750 17196
rect 11238 17184 11244 17196
rect 11199 17156 11244 17184
rect 11238 17144 11244 17156
rect 11296 17144 11302 17196
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 1578 17116 1584 17128
rect 1443 17088 1584 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 1578 17076 1584 17088
rect 1636 17076 1642 17128
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17116 1731 17119
rect 2498 17116 2504 17128
rect 1719 17088 2504 17116
rect 1719 17085 1731 17088
rect 1673 17079 1731 17085
rect 2498 17076 2504 17088
rect 2556 17076 2562 17128
rect 2777 17119 2835 17125
rect 2777 17085 2789 17119
rect 2823 17116 2835 17119
rect 3970 17116 3976 17128
rect 2823 17088 3976 17116
rect 2823 17085 2835 17088
rect 2777 17079 2835 17085
rect 3970 17076 3976 17088
rect 4028 17076 4034 17128
rect 5810 17076 5816 17128
rect 5868 17116 5874 17128
rect 6178 17116 6184 17128
rect 5868 17088 6184 17116
rect 5868 17076 5874 17088
rect 6178 17076 6184 17088
rect 6236 17116 6242 17128
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6236 17088 6837 17116
rect 6236 17076 6242 17088
rect 6825 17085 6837 17088
rect 6871 17116 6883 17119
rect 8202 17116 8208 17128
rect 6871 17088 8208 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 9306 17076 9312 17128
rect 9364 17116 9370 17128
rect 9493 17119 9551 17125
rect 9493 17116 9505 17119
rect 9364 17088 9505 17116
rect 9364 17076 9370 17088
rect 9493 17085 9505 17088
rect 9539 17085 9551 17119
rect 9493 17079 9551 17085
rect 9858 17076 9864 17128
rect 9916 17116 9922 17128
rect 11057 17119 11115 17125
rect 11057 17116 11069 17119
rect 9916 17088 11069 17116
rect 9916 17076 9922 17088
rect 11057 17085 11069 17088
rect 11103 17116 11115 17119
rect 11330 17116 11336 17128
rect 11103 17088 11336 17116
rect 11103 17085 11115 17088
rect 11057 17079 11115 17085
rect 11330 17076 11336 17088
rect 11388 17076 11394 17128
rect 3050 17057 3056 17060
rect 3044 17011 3056 17057
rect 3108 17048 3114 17060
rect 5353 17051 5411 17057
rect 5353 17048 5365 17051
rect 3108 17020 3144 17048
rect 4632 17020 5365 17048
rect 3050 17008 3056 17011
rect 3108 17008 3114 17020
rect 4632 16992 4660 17020
rect 5353 17017 5365 17020
rect 5399 17017 5411 17051
rect 5353 17011 5411 17017
rect 7092 17051 7150 17057
rect 7092 17017 7104 17051
rect 7138 17048 7150 17051
rect 7190 17048 7196 17060
rect 7138 17020 7196 17048
rect 7138 17017 7150 17020
rect 7092 17011 7150 17017
rect 7190 17008 7196 17020
rect 7248 17048 7254 17060
rect 8481 17051 8539 17057
rect 8481 17048 8493 17051
rect 7248 17020 8493 17048
rect 7248 17008 7254 17020
rect 8481 17017 8493 17020
rect 8527 17017 8539 17051
rect 8481 17011 8539 17017
rect 9217 17051 9275 17057
rect 9217 17017 9229 17051
rect 9263 17048 9275 17051
rect 10045 17051 10103 17057
rect 10045 17048 10057 17051
rect 9263 17020 10057 17048
rect 9263 17017 9275 17020
rect 9217 17011 9275 17017
rect 10045 17017 10057 17020
rect 10091 17048 10103 17051
rect 10778 17048 10784 17060
rect 10091 17020 10784 17048
rect 10091 17017 10103 17020
rect 10045 17011 10103 17017
rect 10778 17008 10784 17020
rect 10836 17008 10842 17060
rect 2501 16983 2559 16989
rect 2501 16949 2513 16983
rect 2547 16980 2559 16983
rect 2774 16980 2780 16992
rect 2547 16952 2780 16980
rect 2547 16949 2559 16952
rect 2501 16943 2559 16949
rect 2774 16940 2780 16952
rect 2832 16980 2838 16992
rect 4062 16980 4068 16992
rect 2832 16952 4068 16980
rect 2832 16940 2838 16952
rect 4062 16940 4068 16952
rect 4120 16940 4126 16992
rect 4525 16983 4583 16989
rect 4525 16949 4537 16983
rect 4571 16980 4583 16983
rect 4614 16980 4620 16992
rect 4571 16952 4620 16980
rect 4571 16949 4583 16952
rect 4525 16943 4583 16949
rect 4614 16940 4620 16952
rect 4672 16940 4678 16992
rect 4893 16983 4951 16989
rect 4893 16949 4905 16983
rect 4939 16980 4951 16983
rect 5445 16983 5503 16989
rect 5445 16980 5457 16983
rect 4939 16952 5457 16980
rect 4939 16949 4951 16952
rect 4893 16943 4951 16949
rect 5445 16949 5457 16952
rect 5491 16980 5503 16983
rect 5994 16980 6000 16992
rect 5491 16952 6000 16980
rect 5491 16949 5503 16952
rect 5445 16943 5503 16949
rect 5994 16940 6000 16952
rect 6052 16940 6058 16992
rect 6914 16940 6920 16992
rect 6972 16980 6978 16992
rect 8205 16983 8263 16989
rect 8205 16980 8217 16983
rect 6972 16952 8217 16980
rect 6972 16940 6978 16952
rect 8205 16949 8217 16952
rect 8251 16949 8263 16983
rect 10134 16980 10140 16992
rect 10095 16952 10140 16980
rect 8205 16943 8263 16949
rect 10134 16940 10140 16952
rect 10192 16940 10198 16992
rect 10686 16980 10692 16992
rect 10647 16952 10692 16980
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 11793 16983 11851 16989
rect 11793 16949 11805 16983
rect 11839 16980 11851 16983
rect 12066 16980 12072 16992
rect 11839 16952 12072 16980
rect 11839 16949 11851 16952
rect 11793 16943 11851 16949
rect 12066 16940 12072 16952
rect 12124 16940 12130 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1946 16736 1952 16788
rect 2004 16776 2010 16788
rect 2133 16779 2191 16785
rect 2133 16776 2145 16779
rect 2004 16748 2145 16776
rect 2004 16736 2010 16748
rect 2133 16745 2145 16748
rect 2179 16776 2191 16779
rect 2682 16776 2688 16788
rect 2179 16748 2688 16776
rect 2179 16745 2191 16748
rect 2133 16739 2191 16745
rect 2682 16736 2688 16748
rect 2740 16736 2746 16788
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 3421 16779 3479 16785
rect 3421 16776 3433 16779
rect 2924 16748 3433 16776
rect 2924 16736 2930 16748
rect 3421 16745 3433 16748
rect 3467 16776 3479 16779
rect 4065 16779 4123 16785
rect 4065 16776 4077 16779
rect 3467 16748 4077 16776
rect 3467 16745 3479 16748
rect 3421 16739 3479 16745
rect 4065 16745 4077 16748
rect 4111 16745 4123 16779
rect 7190 16776 7196 16788
rect 7151 16748 7196 16776
rect 4065 16739 4123 16745
rect 7190 16736 7196 16748
rect 7248 16736 7254 16788
rect 8018 16776 8024 16788
rect 7979 16748 8024 16776
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 9493 16779 9551 16785
rect 9493 16745 9505 16779
rect 9539 16776 9551 16779
rect 10134 16776 10140 16788
rect 9539 16748 10140 16776
rect 9539 16745 9551 16748
rect 9493 16739 9551 16745
rect 10134 16736 10140 16748
rect 10192 16736 10198 16788
rect 11330 16776 11336 16788
rect 11291 16748 11336 16776
rect 11330 16736 11336 16748
rect 11388 16736 11394 16788
rect 2777 16711 2835 16717
rect 2777 16677 2789 16711
rect 2823 16708 2835 16711
rect 2958 16708 2964 16720
rect 2823 16680 2964 16708
rect 2823 16677 2835 16680
rect 2777 16671 2835 16677
rect 2958 16668 2964 16680
rect 3016 16668 3022 16720
rect 3050 16668 3056 16720
rect 3108 16708 3114 16720
rect 4154 16708 4160 16720
rect 3108 16680 4160 16708
rect 3108 16668 3114 16680
rect 4154 16668 4160 16680
rect 4212 16668 4218 16720
rect 6086 16717 6092 16720
rect 6080 16708 6092 16717
rect 4264 16680 5580 16708
rect 6047 16680 6092 16708
rect 2041 16643 2099 16649
rect 2041 16609 2053 16643
rect 2087 16640 2099 16643
rect 2130 16640 2136 16652
rect 2087 16612 2136 16640
rect 2087 16609 2099 16612
rect 2041 16603 2099 16609
rect 2130 16600 2136 16612
rect 2188 16640 2194 16652
rect 3142 16640 3148 16652
rect 2188 16612 3148 16640
rect 2188 16600 2194 16612
rect 3142 16600 3148 16612
rect 3200 16600 3206 16652
rect 3881 16643 3939 16649
rect 3881 16609 3893 16643
rect 3927 16640 3939 16643
rect 4264 16640 4292 16680
rect 4430 16640 4436 16652
rect 3927 16612 4292 16640
rect 4391 16612 4436 16640
rect 3927 16609 3939 16612
rect 3881 16603 3939 16609
rect 4430 16600 4436 16612
rect 4488 16600 4494 16652
rect 5552 16584 5580 16680
rect 6080 16671 6092 16680
rect 6086 16668 6092 16671
rect 6144 16668 6150 16720
rect 6914 16668 6920 16720
rect 6972 16708 6978 16720
rect 7466 16708 7472 16720
rect 6972 16680 7472 16708
rect 6972 16668 6978 16680
rect 7466 16668 7472 16680
rect 7524 16668 7530 16720
rect 7929 16711 7987 16717
rect 7929 16677 7941 16711
rect 7975 16708 7987 16711
rect 8202 16708 8208 16720
rect 7975 16680 8208 16708
rect 7975 16677 7987 16680
rect 7929 16671 7987 16677
rect 8202 16668 8208 16680
rect 8260 16668 8266 16720
rect 5810 16640 5816 16652
rect 5771 16612 5816 16640
rect 5810 16600 5816 16612
rect 5868 16600 5874 16652
rect 8018 16600 8024 16652
rect 8076 16640 8082 16652
rect 8389 16643 8447 16649
rect 8389 16640 8401 16643
rect 8076 16612 8401 16640
rect 8076 16600 8082 16612
rect 8389 16609 8401 16612
rect 8435 16609 8447 16643
rect 9858 16640 9864 16652
rect 8389 16603 8447 16609
rect 9600 16612 9864 16640
rect 2222 16572 2228 16584
rect 2183 16544 2228 16572
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 4522 16572 4528 16584
rect 4483 16544 4528 16572
rect 4522 16532 4528 16544
rect 4580 16532 4586 16584
rect 4617 16575 4675 16581
rect 4617 16541 4629 16575
rect 4663 16541 4675 16575
rect 4617 16535 4675 16541
rect 3697 16507 3755 16513
rect 3697 16473 3709 16507
rect 3743 16504 3755 16507
rect 3970 16504 3976 16516
rect 3743 16476 3976 16504
rect 3743 16473 3755 16476
rect 3697 16467 3755 16473
rect 3970 16464 3976 16476
rect 4028 16464 4034 16516
rect 4154 16464 4160 16516
rect 4212 16504 4218 16516
rect 4632 16504 4660 16535
rect 5534 16532 5540 16584
rect 5592 16532 5598 16584
rect 8481 16575 8539 16581
rect 8481 16541 8493 16575
rect 8527 16541 8539 16575
rect 8662 16572 8668 16584
rect 8623 16544 8668 16572
rect 8481 16535 8539 16541
rect 4212 16476 4660 16504
rect 5169 16507 5227 16513
rect 4212 16464 4218 16476
rect 5169 16473 5181 16507
rect 5215 16504 5227 16507
rect 5350 16504 5356 16516
rect 5215 16476 5356 16504
rect 5215 16473 5227 16476
rect 5169 16467 5227 16473
rect 5350 16464 5356 16476
rect 5408 16464 5414 16516
rect 8386 16464 8392 16516
rect 8444 16504 8450 16516
rect 8496 16504 8524 16535
rect 8662 16532 8668 16544
rect 8720 16572 8726 16584
rect 9600 16572 9628 16612
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 10042 16600 10048 16652
rect 10100 16640 10106 16652
rect 10209 16643 10267 16649
rect 10209 16640 10221 16643
rect 10100 16612 10221 16640
rect 10100 16600 10106 16612
rect 10209 16609 10221 16612
rect 10255 16640 10267 16643
rect 10686 16640 10692 16652
rect 10255 16612 10692 16640
rect 10255 16609 10267 16612
rect 10209 16603 10267 16609
rect 10686 16600 10692 16612
rect 10744 16600 10750 16652
rect 8720 16544 9628 16572
rect 8720 16532 8726 16544
rect 9766 16532 9772 16584
rect 9824 16572 9830 16584
rect 9950 16572 9956 16584
rect 9824 16544 9956 16572
rect 9824 16532 9830 16544
rect 9950 16532 9956 16544
rect 10008 16532 10014 16584
rect 8444 16476 8524 16504
rect 8444 16464 8450 16476
rect 1486 16396 1492 16448
rect 1544 16436 1550 16448
rect 1673 16439 1731 16445
rect 1673 16436 1685 16439
rect 1544 16408 1685 16436
rect 1544 16396 1550 16408
rect 1673 16405 1685 16408
rect 1719 16405 1731 16439
rect 5442 16436 5448 16448
rect 5403 16408 5448 16436
rect 1673 16399 1731 16405
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 9125 16439 9183 16445
rect 9125 16405 9137 16439
rect 9171 16436 9183 16439
rect 9214 16436 9220 16448
rect 9171 16408 9220 16436
rect 9171 16405 9183 16408
rect 9125 16399 9183 16405
rect 9214 16396 9220 16408
rect 9272 16396 9278 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2222 16232 2228 16244
rect 2183 16204 2228 16232
rect 2222 16192 2228 16204
rect 2280 16232 2286 16244
rect 2682 16232 2688 16244
rect 2280 16204 2688 16232
rect 2280 16192 2286 16204
rect 2682 16192 2688 16204
rect 2740 16192 2746 16244
rect 4154 16232 4160 16244
rect 4115 16204 4160 16232
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 5074 16232 5080 16244
rect 5035 16204 5080 16232
rect 5074 16192 5080 16204
rect 5132 16192 5138 16244
rect 6086 16232 6092 16244
rect 6047 16204 6092 16232
rect 6086 16192 6092 16204
rect 6144 16192 6150 16244
rect 10134 16192 10140 16244
rect 10192 16232 10198 16244
rect 10229 16235 10287 16241
rect 10229 16232 10241 16235
rect 10192 16204 10241 16232
rect 10192 16192 10198 16204
rect 10229 16201 10241 16204
rect 10275 16201 10287 16235
rect 10229 16195 10287 16201
rect 1670 16096 1676 16108
rect 1631 16068 1676 16096
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 5442 16056 5448 16108
rect 5500 16096 5506 16108
rect 5721 16099 5779 16105
rect 5721 16096 5733 16099
rect 5500 16068 5733 16096
rect 5500 16056 5506 16068
rect 5721 16065 5733 16068
rect 5767 16096 5779 16099
rect 6086 16096 6092 16108
rect 5767 16068 6092 16096
rect 5767 16065 5779 16068
rect 5721 16059 5779 16065
rect 6086 16056 6092 16068
rect 6144 16056 6150 16108
rect 9401 16099 9459 16105
rect 9401 16065 9413 16099
rect 9447 16096 9459 16099
rect 10686 16096 10692 16108
rect 9447 16068 10692 16096
rect 9447 16065 9459 16068
rect 9401 16059 9459 16065
rect 10686 16056 10692 16068
rect 10744 16096 10750 16108
rect 10781 16099 10839 16105
rect 10781 16096 10793 16099
rect 10744 16068 10793 16096
rect 10744 16056 10750 16068
rect 10781 16065 10793 16068
rect 10827 16065 10839 16099
rect 10781 16059 10839 16065
rect 12434 16056 12440 16108
rect 12492 16096 12498 16108
rect 12492 16068 12537 16096
rect 12492 16056 12498 16068
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1486 16028 1492 16040
rect 1443 16000 1492 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1486 15988 1492 16000
rect 1544 15988 1550 16040
rect 2777 16031 2835 16037
rect 2777 15997 2789 16031
rect 2823 16028 2835 16031
rect 3970 16028 3976 16040
rect 2823 16000 3976 16028
rect 2823 15997 2835 16000
rect 2777 15991 2835 15997
rect 3970 15988 3976 16000
rect 4028 15988 4034 16040
rect 4430 15988 4436 16040
rect 4488 16028 4494 16040
rect 4893 16031 4951 16037
rect 4893 16028 4905 16031
rect 4488 16000 4905 16028
rect 4488 15988 4494 16000
rect 4893 15997 4905 16000
rect 4939 16028 4951 16031
rect 7377 16031 7435 16037
rect 4939 16000 7328 16028
rect 4939 15997 4951 16000
rect 4893 15991 4951 15997
rect 2685 15963 2743 15969
rect 2685 15929 2697 15963
rect 2731 15960 2743 15963
rect 2958 15960 2964 15972
rect 2731 15932 2964 15960
rect 2731 15929 2743 15932
rect 2685 15923 2743 15929
rect 2958 15920 2964 15932
rect 3016 15969 3022 15972
rect 3016 15963 3080 15969
rect 3016 15929 3034 15963
rect 3068 15929 3080 15963
rect 3016 15923 3080 15929
rect 5537 15963 5595 15969
rect 5537 15929 5549 15963
rect 5583 15960 5595 15963
rect 5583 15932 6592 15960
rect 5583 15929 5595 15932
rect 5537 15923 5595 15929
rect 3016 15920 3022 15923
rect 4522 15892 4528 15904
rect 4435 15864 4528 15892
rect 4522 15852 4528 15864
rect 4580 15892 4586 15904
rect 4982 15892 4988 15904
rect 4580 15864 4988 15892
rect 4580 15852 4586 15864
rect 4982 15852 4988 15864
rect 5040 15852 5046 15904
rect 5350 15852 5356 15904
rect 5408 15892 5414 15904
rect 6564 15901 6592 15932
rect 5445 15895 5503 15901
rect 5445 15892 5457 15895
rect 5408 15864 5457 15892
rect 5408 15852 5414 15864
rect 5445 15861 5457 15864
rect 5491 15861 5503 15895
rect 5445 15855 5503 15861
rect 6549 15895 6607 15901
rect 6549 15861 6561 15895
rect 6595 15892 6607 15895
rect 6822 15892 6828 15904
rect 6595 15864 6828 15892
rect 6595 15861 6607 15864
rect 6549 15855 6607 15861
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 7300 15901 7328 16000
rect 7377 15997 7389 16031
rect 7423 15997 7435 16031
rect 7377 15991 7435 15997
rect 7392 15960 7420 15991
rect 7466 15988 7472 16040
rect 7524 16028 7530 16040
rect 7633 16031 7691 16037
rect 7633 16028 7645 16031
rect 7524 16000 7645 16028
rect 7524 15988 7530 16000
rect 7633 15997 7645 16000
rect 7679 15997 7691 16031
rect 7633 15991 7691 15997
rect 8202 15960 8208 15972
rect 7392 15932 8208 15960
rect 8202 15920 8208 15932
rect 8260 15920 8266 15972
rect 10137 15963 10195 15969
rect 10137 15929 10149 15963
rect 10183 15960 10195 15963
rect 10689 15963 10747 15969
rect 10689 15960 10701 15963
rect 10183 15932 10701 15960
rect 10183 15929 10195 15932
rect 10137 15923 10195 15929
rect 10689 15929 10701 15932
rect 10735 15960 10747 15963
rect 11330 15960 11336 15972
rect 10735 15932 11336 15960
rect 10735 15929 10747 15932
rect 10689 15923 10747 15929
rect 11330 15920 11336 15932
rect 11388 15920 11394 15972
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 8018 15892 8024 15904
rect 7331 15864 8024 15892
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 8018 15852 8024 15864
rect 8076 15852 8082 15904
rect 8754 15892 8760 15904
rect 8715 15864 8760 15892
rect 8754 15852 8760 15864
rect 8812 15852 8818 15904
rect 9766 15892 9772 15904
rect 9679 15864 9772 15892
rect 9766 15852 9772 15864
rect 9824 15892 9830 15904
rect 10597 15895 10655 15901
rect 10597 15892 10609 15895
rect 9824 15864 10609 15892
rect 9824 15852 9830 15864
rect 10597 15861 10609 15864
rect 10643 15861 10655 15895
rect 11238 15892 11244 15904
rect 11151 15864 11244 15892
rect 10597 15855 10655 15861
rect 11238 15852 11244 15864
rect 11296 15892 11302 15904
rect 11701 15895 11759 15901
rect 11701 15892 11713 15895
rect 11296 15864 11713 15892
rect 11296 15852 11302 15864
rect 11701 15861 11713 15864
rect 11747 15892 11759 15895
rect 11790 15892 11796 15904
rect 11747 15864 11796 15892
rect 11747 15861 11759 15864
rect 11701 15855 11759 15861
rect 11790 15852 11796 15864
rect 11848 15852 11854 15904
rect 12066 15892 12072 15904
rect 12027 15864 12072 15892
rect 12066 15852 12072 15864
rect 12124 15852 12130 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1762 15648 1768 15700
rect 1820 15688 1826 15700
rect 2409 15691 2467 15697
rect 2409 15688 2421 15691
rect 1820 15660 2421 15688
rect 1820 15648 1826 15660
rect 2409 15657 2421 15660
rect 2455 15657 2467 15691
rect 2409 15651 2467 15657
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 3789 15691 3847 15697
rect 3789 15688 3801 15691
rect 2832 15660 3801 15688
rect 2832 15648 2838 15660
rect 3789 15657 3801 15660
rect 3835 15657 3847 15691
rect 4062 15688 4068 15700
rect 4023 15660 4068 15688
rect 3789 15651 3847 15657
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 4154 15648 4160 15700
rect 4212 15688 4218 15700
rect 4525 15691 4583 15697
rect 4525 15688 4537 15691
rect 4212 15660 4537 15688
rect 4212 15648 4218 15660
rect 4525 15657 4537 15660
rect 4571 15657 4583 15691
rect 4525 15651 4583 15657
rect 5626 15648 5632 15700
rect 5684 15688 5690 15700
rect 6730 15688 6736 15700
rect 5684 15660 6736 15688
rect 5684 15648 5690 15660
rect 6730 15648 6736 15660
rect 6788 15648 6794 15700
rect 7282 15688 7288 15700
rect 7243 15660 7288 15688
rect 7282 15648 7288 15660
rect 7340 15648 7346 15700
rect 8662 15688 8668 15700
rect 8623 15660 8668 15688
rect 8662 15648 8668 15660
rect 8720 15648 8726 15700
rect 10042 15688 10048 15700
rect 9955 15660 10048 15688
rect 10042 15648 10048 15660
rect 10100 15688 10106 15700
rect 11701 15691 11759 15697
rect 11701 15688 11713 15691
rect 10100 15660 11713 15688
rect 10100 15648 10106 15660
rect 11701 15657 11713 15660
rect 11747 15657 11759 15691
rect 11701 15651 11759 15657
rect 2317 15623 2375 15629
rect 2317 15589 2329 15623
rect 2363 15620 2375 15623
rect 2958 15620 2964 15632
rect 2363 15592 2964 15620
rect 2363 15589 2375 15592
rect 2317 15583 2375 15589
rect 2958 15580 2964 15592
rect 3016 15580 3022 15632
rect 4985 15623 5043 15629
rect 4985 15589 4997 15623
rect 5031 15620 5043 15623
rect 5322 15623 5380 15629
rect 5322 15620 5334 15623
rect 5031 15592 5334 15620
rect 5031 15589 5043 15592
rect 4985 15583 5043 15589
rect 5322 15589 5334 15592
rect 5368 15620 5380 15623
rect 5534 15620 5540 15632
rect 5368 15592 5540 15620
rect 5368 15589 5380 15592
rect 5322 15583 5380 15589
rect 5534 15580 5540 15592
rect 5592 15580 5598 15632
rect 10588 15623 10646 15629
rect 10588 15589 10600 15623
rect 10634 15620 10646 15623
rect 10686 15620 10692 15632
rect 10634 15592 10692 15620
rect 10634 15589 10646 15592
rect 10588 15583 10646 15589
rect 10686 15580 10692 15592
rect 10744 15620 10750 15632
rect 11054 15620 11060 15632
rect 10744 15592 11060 15620
rect 10744 15580 10750 15592
rect 11054 15580 11060 15592
rect 11112 15580 11118 15632
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 2777 15555 2835 15561
rect 2777 15552 2789 15555
rect 1443 15524 2789 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 2777 15521 2789 15524
rect 2823 15552 2835 15555
rect 3050 15552 3056 15564
rect 2823 15524 3056 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 3050 15512 3056 15524
rect 3108 15512 3114 15564
rect 5077 15555 5135 15561
rect 5077 15521 5089 15555
rect 5123 15552 5135 15555
rect 5166 15552 5172 15564
rect 5123 15524 5172 15552
rect 5123 15521 5135 15524
rect 5077 15515 5135 15521
rect 5166 15512 5172 15524
rect 5224 15512 5230 15564
rect 7650 15552 7656 15564
rect 7611 15524 7656 15552
rect 7650 15512 7656 15524
rect 7708 15512 7714 15564
rect 9306 15552 9312 15564
rect 9267 15524 9312 15552
rect 9306 15512 9312 15524
rect 9364 15512 9370 15564
rect 9950 15512 9956 15564
rect 10008 15552 10014 15564
rect 10321 15555 10379 15561
rect 10321 15552 10333 15555
rect 10008 15524 10333 15552
rect 10008 15512 10014 15524
rect 10321 15521 10333 15524
rect 10367 15552 10379 15555
rect 12066 15552 12072 15564
rect 10367 15524 12072 15552
rect 10367 15521 10379 15524
rect 10321 15515 10379 15521
rect 12066 15512 12072 15524
rect 12124 15512 12130 15564
rect 2869 15487 2927 15493
rect 2869 15453 2881 15487
rect 2915 15453 2927 15487
rect 2869 15447 2927 15453
rect 2884 15416 2912 15447
rect 2958 15444 2964 15496
rect 3016 15484 3022 15496
rect 3016 15456 4200 15484
rect 3016 15444 3022 15456
rect 3513 15419 3571 15425
rect 3513 15416 3525 15419
rect 2884 15388 3525 15416
rect 3513 15385 3525 15388
rect 3559 15416 3571 15419
rect 3559 15388 4108 15416
rect 3559 15385 3571 15388
rect 3513 15379 3571 15385
rect 4080 15360 4108 15388
rect 1946 15348 1952 15360
rect 1907 15320 1952 15348
rect 1946 15308 1952 15320
rect 2004 15308 2010 15360
rect 4062 15308 4068 15360
rect 4120 15308 4126 15360
rect 4172 15348 4200 15456
rect 7282 15444 7288 15496
rect 7340 15484 7346 15496
rect 7745 15487 7803 15493
rect 7745 15484 7757 15487
rect 7340 15456 7757 15484
rect 7340 15444 7346 15456
rect 7745 15453 7757 15456
rect 7791 15453 7803 15487
rect 7745 15447 7803 15453
rect 7837 15487 7895 15493
rect 7837 15453 7849 15487
rect 7883 15453 7895 15487
rect 7837 15447 7895 15453
rect 7852 15416 7880 15447
rect 7116 15388 7880 15416
rect 6457 15351 6515 15357
rect 6457 15348 6469 15351
rect 4172 15320 6469 15348
rect 6457 15317 6469 15320
rect 6503 15317 6515 15351
rect 6457 15311 6515 15317
rect 7006 15308 7012 15360
rect 7064 15348 7070 15360
rect 7116 15357 7144 15388
rect 7101 15351 7159 15357
rect 7101 15348 7113 15351
rect 7064 15320 7113 15348
rect 7064 15308 7070 15320
rect 7101 15317 7113 15320
rect 7147 15317 7159 15351
rect 8386 15348 8392 15360
rect 8347 15320 8392 15348
rect 7101 15311 7159 15317
rect 8386 15308 8392 15320
rect 8444 15308 8450 15360
rect 9125 15351 9183 15357
rect 9125 15317 9137 15351
rect 9171 15348 9183 15351
rect 9214 15348 9220 15360
rect 9171 15320 9220 15348
rect 9171 15317 9183 15320
rect 9125 15311 9183 15317
rect 9214 15308 9220 15320
rect 9272 15308 9278 15360
rect 12066 15348 12072 15360
rect 12027 15320 12072 15348
rect 12066 15308 12072 15320
rect 12124 15308 12130 15360
rect 12529 15351 12587 15357
rect 12529 15317 12541 15351
rect 12575 15348 12587 15351
rect 12802 15348 12808 15360
rect 12575 15320 12808 15348
rect 12575 15317 12587 15320
rect 12529 15311 12587 15317
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2038 15144 2044 15156
rect 1999 15116 2044 15144
rect 2038 15104 2044 15116
rect 2096 15104 2102 15156
rect 3050 15144 3056 15156
rect 3011 15116 3056 15144
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 3510 15104 3516 15156
rect 3568 15144 3574 15156
rect 3605 15147 3663 15153
rect 3605 15144 3617 15147
rect 3568 15116 3617 15144
rect 3568 15104 3574 15116
rect 3605 15113 3617 15116
rect 3651 15113 3663 15147
rect 3605 15107 3663 15113
rect 4154 15104 4160 15156
rect 4212 15144 4218 15156
rect 5169 15147 5227 15153
rect 5169 15144 5181 15147
rect 4212 15116 5181 15144
rect 4212 15104 4218 15116
rect 5169 15113 5181 15116
rect 5215 15113 5227 15147
rect 8110 15144 8116 15156
rect 5169 15107 5227 15113
rect 7760 15116 8116 15144
rect 1946 14968 1952 15020
rect 2004 15008 2010 15020
rect 2593 15011 2651 15017
rect 2593 15008 2605 15011
rect 2004 14980 2605 15008
rect 2004 14968 2010 14980
rect 2593 14977 2605 14980
rect 2639 14977 2651 15011
rect 2593 14971 2651 14977
rect 3510 14968 3516 15020
rect 3568 15008 3574 15020
rect 4157 15011 4215 15017
rect 4157 15008 4169 15011
rect 3568 14980 4169 15008
rect 3568 14968 3574 14980
rect 4157 14977 4169 14980
rect 4203 14977 4215 15011
rect 4157 14971 4215 14977
rect 5534 14968 5540 15020
rect 5592 15008 5598 15020
rect 5721 15011 5779 15017
rect 5721 15008 5733 15011
rect 5592 14980 5733 15008
rect 5592 14968 5598 14980
rect 5721 14977 5733 14980
rect 5767 15008 5779 15011
rect 6181 15011 6239 15017
rect 6181 15008 6193 15011
rect 5767 14980 6193 15008
rect 5767 14977 5779 14980
rect 5721 14971 5779 14977
rect 6181 14977 6193 14980
rect 6227 15008 6239 15011
rect 6362 15008 6368 15020
rect 6227 14980 6368 15008
rect 6227 14977 6239 14980
rect 6181 14971 6239 14977
rect 6362 14968 6368 14980
rect 6420 14968 6426 15020
rect 7760 15017 7788 15116
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 9674 15104 9680 15156
rect 9732 15144 9738 15156
rect 9953 15147 10011 15153
rect 9953 15144 9965 15147
rect 9732 15116 9965 15144
rect 9732 15104 9738 15116
rect 9953 15113 9965 15116
rect 9999 15113 10011 15147
rect 11054 15144 11060 15156
rect 11015 15116 11060 15144
rect 9953 15107 10011 15113
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 7745 15011 7803 15017
rect 7745 14977 7757 15011
rect 7791 14977 7803 15011
rect 7745 14971 7803 14977
rect 10597 15011 10655 15017
rect 10597 14977 10609 15011
rect 10643 15008 10655 15011
rect 10686 15008 10692 15020
rect 10643 14980 10692 15008
rect 10643 14977 10655 14980
rect 10597 14971 10655 14977
rect 10686 14968 10692 14980
rect 10744 14968 10750 15020
rect 11882 15008 11888 15020
rect 11795 14980 11888 15008
rect 11882 14968 11888 14980
rect 11940 15008 11946 15020
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 11940 14980 13001 15008
rect 11940 14968 11946 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 2409 14943 2467 14949
rect 2409 14909 2421 14943
rect 2455 14940 2467 14943
rect 2682 14940 2688 14952
rect 2455 14912 2688 14940
rect 2455 14909 2467 14912
rect 2409 14903 2467 14909
rect 2682 14900 2688 14912
rect 2740 14900 2746 14952
rect 12802 14940 12808 14952
rect 3160 14912 4844 14940
rect 12763 14912 12808 14940
rect 1949 14875 2007 14881
rect 1949 14841 1961 14875
rect 1995 14872 2007 14875
rect 2501 14875 2559 14881
rect 2501 14872 2513 14875
rect 1995 14844 2513 14872
rect 1995 14841 2007 14844
rect 1949 14835 2007 14841
rect 2501 14841 2513 14844
rect 2547 14872 2559 14875
rect 3160 14872 3188 14912
rect 2547 14844 3188 14872
rect 4065 14875 4123 14881
rect 2547 14841 2559 14844
rect 2501 14835 2559 14841
rect 4065 14841 4077 14875
rect 4111 14872 4123 14875
rect 4706 14872 4712 14884
rect 4111 14844 4712 14872
rect 4111 14841 4123 14844
rect 4065 14835 4123 14841
rect 4706 14832 4712 14844
rect 4764 14832 4770 14884
rect 3510 14804 3516 14816
rect 3471 14776 3516 14804
rect 3510 14764 3516 14776
rect 3568 14764 3574 14816
rect 3602 14764 3608 14816
rect 3660 14804 3666 14816
rect 3973 14807 4031 14813
rect 3973 14804 3985 14807
rect 3660 14776 3985 14804
rect 3660 14764 3666 14776
rect 3973 14773 3985 14776
rect 4019 14773 4031 14807
rect 3973 14767 4031 14773
rect 4617 14807 4675 14813
rect 4617 14773 4629 14807
rect 4663 14804 4675 14807
rect 4816 14804 4844 14912
rect 12802 14900 12808 14912
rect 12860 14900 12866 14952
rect 5077 14875 5135 14881
rect 5077 14841 5089 14875
rect 5123 14872 5135 14875
rect 6641 14875 6699 14881
rect 5123 14844 5672 14872
rect 5123 14841 5135 14844
rect 5077 14835 5135 14841
rect 5644 14816 5672 14844
rect 6641 14841 6653 14875
rect 6687 14872 6699 14875
rect 7650 14872 7656 14884
rect 6687 14844 7656 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 7650 14832 7656 14844
rect 7708 14832 7714 14884
rect 8012 14875 8070 14881
rect 8012 14841 8024 14875
rect 8058 14872 8070 14875
rect 8662 14872 8668 14884
rect 8058 14844 8668 14872
rect 8058 14841 8070 14844
rect 8012 14835 8070 14841
rect 8662 14832 8668 14844
rect 8720 14832 8726 14884
rect 9493 14875 9551 14881
rect 9493 14841 9505 14875
rect 9539 14872 9551 14875
rect 10042 14872 10048 14884
rect 9539 14844 10048 14872
rect 9539 14841 9551 14844
rect 9493 14835 9551 14841
rect 10042 14832 10048 14844
rect 10100 14872 10106 14884
rect 10413 14875 10471 14881
rect 10413 14872 10425 14875
rect 10100 14844 10425 14872
rect 10100 14832 10106 14844
rect 10413 14841 10425 14844
rect 10459 14841 10471 14875
rect 10413 14835 10471 14841
rect 10870 14832 10876 14884
rect 10928 14872 10934 14884
rect 12161 14875 12219 14881
rect 12161 14872 12173 14875
rect 10928 14844 12173 14872
rect 10928 14832 10934 14844
rect 12161 14841 12173 14844
rect 12207 14872 12219 14875
rect 12897 14875 12955 14881
rect 12897 14872 12909 14875
rect 12207 14844 12909 14872
rect 12207 14841 12219 14844
rect 12161 14835 12219 14841
rect 12897 14841 12909 14844
rect 12943 14841 12955 14875
rect 12897 14835 12955 14841
rect 4890 14804 4896 14816
rect 4663 14776 4896 14804
rect 4663 14773 4675 14776
rect 4617 14767 4675 14773
rect 4890 14764 4896 14776
rect 4948 14804 4954 14816
rect 5534 14804 5540 14816
rect 4948 14776 5540 14804
rect 4948 14764 4954 14776
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 5626 14764 5632 14816
rect 5684 14804 5690 14816
rect 7282 14804 7288 14816
rect 5684 14776 5729 14804
rect 7243 14776 7288 14804
rect 5684 14764 5690 14776
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 9122 14804 9128 14816
rect 9083 14776 9128 14804
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 9861 14807 9919 14813
rect 9861 14773 9873 14807
rect 9907 14804 9919 14807
rect 10321 14807 10379 14813
rect 10321 14804 10333 14807
rect 9907 14776 10333 14804
rect 9907 14773 9919 14776
rect 9861 14767 9919 14773
rect 10321 14773 10333 14776
rect 10367 14804 10379 14807
rect 10778 14804 10784 14816
rect 10367 14776 10784 14804
rect 10367 14773 10379 14776
rect 10321 14767 10379 14773
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 11425 14807 11483 14813
rect 11425 14773 11437 14807
rect 11471 14804 11483 14807
rect 11882 14804 11888 14816
rect 11471 14776 11888 14804
rect 11471 14773 11483 14776
rect 11425 14767 11483 14773
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 12250 14764 12256 14816
rect 12308 14804 12314 14816
rect 12437 14807 12495 14813
rect 12437 14804 12449 14807
rect 12308 14776 12449 14804
rect 12308 14764 12314 14776
rect 12437 14773 12449 14776
rect 12483 14773 12495 14807
rect 12437 14767 12495 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1394 14600 1400 14612
rect 1355 14572 1400 14600
rect 1394 14560 1400 14572
rect 1452 14560 1458 14612
rect 2409 14603 2467 14609
rect 2409 14569 2421 14603
rect 2455 14600 2467 14603
rect 2590 14600 2596 14612
rect 2455 14572 2596 14600
rect 2455 14569 2467 14572
rect 2409 14563 2467 14569
rect 2590 14560 2596 14572
rect 2648 14560 2654 14612
rect 3142 14560 3148 14612
rect 3200 14600 3206 14612
rect 3789 14603 3847 14609
rect 3789 14600 3801 14603
rect 3200 14572 3801 14600
rect 3200 14560 3206 14572
rect 3789 14569 3801 14572
rect 3835 14569 3847 14603
rect 4246 14600 4252 14612
rect 4207 14572 4252 14600
rect 3789 14563 3847 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 6362 14600 6368 14612
rect 6323 14572 6368 14600
rect 6362 14560 6368 14572
rect 6420 14560 6426 14612
rect 6914 14560 6920 14612
rect 6972 14600 6978 14612
rect 7193 14603 7251 14609
rect 7193 14600 7205 14603
rect 6972 14572 7205 14600
rect 6972 14560 6978 14572
rect 7193 14569 7205 14572
rect 7239 14569 7251 14603
rect 8662 14600 8668 14612
rect 8623 14572 8668 14600
rect 7193 14563 7251 14569
rect 8662 14560 8668 14572
rect 8720 14560 8726 14612
rect 8754 14560 8760 14612
rect 8812 14600 8818 14612
rect 9306 14600 9312 14612
rect 8812 14572 8857 14600
rect 9267 14572 9312 14600
rect 8812 14560 8818 14572
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 11054 14560 11060 14612
rect 11112 14600 11118 14612
rect 11609 14603 11667 14609
rect 11609 14600 11621 14603
rect 11112 14572 11621 14600
rect 11112 14560 11118 14572
rect 11609 14569 11621 14572
rect 11655 14569 11667 14603
rect 11882 14600 11888 14612
rect 11843 14572 11888 14600
rect 11609 14563 11667 14569
rect 11882 14560 11888 14572
rect 11940 14560 11946 14612
rect 12066 14560 12072 14612
rect 12124 14600 12130 14612
rect 12253 14603 12311 14609
rect 12253 14600 12265 14603
rect 12124 14572 12265 14600
rect 12124 14560 12130 14572
rect 12253 14569 12265 14572
rect 12299 14569 12311 14603
rect 12253 14563 12311 14569
rect 12437 14603 12495 14609
rect 12437 14569 12449 14603
rect 12483 14600 12495 14603
rect 12618 14600 12624 14612
rect 12483 14572 12624 14600
rect 12483 14569 12495 14572
rect 12437 14563 12495 14569
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 2133 14535 2191 14541
rect 2133 14501 2145 14535
rect 2179 14532 2191 14535
rect 2682 14532 2688 14544
rect 2179 14504 2688 14532
rect 2179 14501 2191 14504
rect 2133 14495 2191 14501
rect 2682 14492 2688 14504
rect 2740 14492 2746 14544
rect 2869 14535 2927 14541
rect 2869 14501 2881 14535
rect 2915 14532 2927 14535
rect 3970 14532 3976 14544
rect 2915 14504 3976 14532
rect 2915 14501 2927 14504
rect 2869 14495 2927 14501
rect 3970 14492 3976 14504
rect 4028 14492 4034 14544
rect 7561 14535 7619 14541
rect 7561 14501 7573 14535
rect 7607 14532 7619 14535
rect 7742 14532 7748 14544
rect 7607 14504 7748 14532
rect 7607 14501 7619 14504
rect 7561 14495 7619 14501
rect 7742 14492 7748 14504
rect 7800 14492 7806 14544
rect 8110 14492 8116 14544
rect 8168 14532 8174 14544
rect 8297 14535 8355 14541
rect 8297 14532 8309 14535
rect 8168 14504 8309 14532
rect 8168 14492 8174 14504
rect 8297 14501 8309 14504
rect 8343 14532 8355 14535
rect 9122 14532 9128 14544
rect 8343 14504 9128 14532
rect 8343 14501 8355 14504
rect 8297 14495 8355 14501
rect 9122 14492 9128 14504
rect 9180 14492 9186 14544
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 2832 14436 2877 14464
rect 2832 14424 2838 14436
rect 3326 14424 3332 14476
rect 3384 14464 3390 14476
rect 3421 14467 3479 14473
rect 3421 14464 3433 14467
rect 3384 14436 3433 14464
rect 3384 14424 3390 14436
rect 3421 14433 3433 14436
rect 3467 14433 3479 14467
rect 3421 14427 3479 14433
rect 4985 14467 5043 14473
rect 4985 14433 4997 14467
rect 5031 14464 5043 14467
rect 5074 14464 5080 14476
rect 5031 14436 5080 14464
rect 5031 14433 5043 14436
rect 4985 14427 5043 14433
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 5258 14473 5264 14476
rect 5252 14464 5264 14473
rect 5219 14436 5264 14464
rect 5252 14427 5264 14436
rect 5258 14424 5264 14427
rect 5316 14424 5322 14476
rect 8941 14467 8999 14473
rect 8941 14433 8953 14467
rect 8987 14464 8999 14467
rect 9324 14464 9352 14560
rect 10045 14535 10103 14541
rect 10045 14501 10057 14535
rect 10091 14532 10103 14535
rect 10496 14535 10554 14541
rect 10496 14532 10508 14535
rect 10091 14504 10508 14532
rect 10091 14501 10103 14504
rect 10045 14495 10103 14501
rect 10496 14501 10508 14504
rect 10542 14532 10554 14535
rect 10686 14532 10692 14544
rect 10542 14504 10692 14532
rect 10542 14501 10554 14504
rect 10496 14495 10554 14501
rect 10686 14492 10692 14504
rect 10744 14532 10750 14544
rect 11146 14532 11152 14544
rect 10744 14504 11152 14532
rect 10744 14492 10750 14504
rect 11146 14492 11152 14504
rect 11204 14492 11210 14544
rect 8987 14436 9352 14464
rect 8987 14433 8999 14436
rect 8941 14427 8999 14433
rect 10134 14424 10140 14476
rect 10192 14464 10198 14476
rect 10229 14467 10287 14473
rect 10229 14464 10241 14467
rect 10192 14436 10241 14464
rect 10192 14424 10198 14436
rect 10229 14433 10241 14436
rect 10275 14464 10287 14467
rect 11900 14464 11928 14560
rect 12805 14535 12863 14541
rect 12805 14501 12817 14535
rect 12851 14532 12863 14535
rect 12894 14532 12900 14544
rect 12851 14504 12900 14532
rect 12851 14501 12863 14504
rect 12805 14495 12863 14501
rect 12894 14492 12900 14504
rect 12952 14492 12958 14544
rect 23474 14464 23480 14476
rect 10275 14436 11928 14464
rect 23435 14436 23480 14464
rect 10275 14433 10287 14436
rect 10229 14427 10287 14433
rect 23474 14424 23480 14436
rect 23532 14424 23538 14476
rect 3050 14396 3056 14408
rect 3011 14368 3056 14396
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 4706 14396 4712 14408
rect 4667 14368 4712 14396
rect 4706 14356 4712 14368
rect 4764 14356 4770 14408
rect 6914 14356 6920 14408
rect 6972 14396 6978 14408
rect 7653 14399 7711 14405
rect 7653 14396 7665 14399
rect 6972 14368 7665 14396
rect 6972 14356 6978 14368
rect 7653 14365 7665 14368
rect 7699 14365 7711 14399
rect 7834 14396 7840 14408
rect 7795 14368 7840 14396
rect 7653 14359 7711 14365
rect 7834 14356 7840 14368
rect 7892 14356 7898 14408
rect 12250 14356 12256 14408
rect 12308 14396 12314 14408
rect 12897 14399 12955 14405
rect 12897 14396 12909 14399
rect 12308 14368 12909 14396
rect 12308 14356 12314 14368
rect 12897 14365 12909 14368
rect 12943 14365 12955 14399
rect 12897 14359 12955 14365
rect 12986 14356 12992 14408
rect 13044 14396 13050 14408
rect 13044 14368 13089 14396
rect 13044 14356 13050 14368
rect 5994 14288 6000 14340
rect 6052 14328 6058 14340
rect 8938 14328 8944 14340
rect 6052 14300 8944 14328
rect 6052 14288 6058 14300
rect 8938 14288 8944 14300
rect 8996 14288 9002 14340
rect 6362 14220 6368 14272
rect 6420 14260 6426 14272
rect 6641 14263 6699 14269
rect 6641 14260 6653 14263
rect 6420 14232 6653 14260
rect 6420 14220 6426 14232
rect 6641 14229 6653 14232
rect 6687 14260 6699 14263
rect 7009 14263 7067 14269
rect 7009 14260 7021 14263
rect 6687 14232 7021 14260
rect 6687 14229 6699 14232
rect 6641 14223 6699 14229
rect 7009 14229 7021 14232
rect 7055 14229 7067 14263
rect 7009 14223 7067 14229
rect 23661 14263 23719 14269
rect 23661 14229 23673 14263
rect 23707 14260 23719 14263
rect 24946 14260 24952 14272
rect 23707 14232 24952 14260
rect 23707 14229 23719 14232
rect 23661 14223 23719 14229
rect 24946 14220 24952 14232
rect 25004 14220 25010 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2866 14016 2872 14068
rect 2924 14056 2930 14068
rect 3326 14056 3332 14068
rect 2924 14028 3332 14056
rect 2924 14016 2930 14028
rect 3326 14016 3332 14028
rect 3384 14016 3390 14068
rect 4062 14056 4068 14068
rect 4023 14028 4068 14056
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 6638 14056 6644 14068
rect 6551 14028 6644 14056
rect 6638 14016 6644 14028
rect 6696 14056 6702 14068
rect 7834 14056 7840 14068
rect 6696 14028 7840 14056
rect 6696 14016 6702 14028
rect 7834 14016 7840 14028
rect 7892 14016 7898 14068
rect 10042 14056 10048 14068
rect 10003 14028 10048 14056
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 11790 14056 11796 14068
rect 11751 14028 11796 14056
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 12250 14056 12256 14068
rect 12211 14028 12256 14056
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 12986 14016 12992 14068
rect 13044 14056 13050 14068
rect 13265 14059 13323 14065
rect 13265 14056 13277 14059
rect 13044 14028 13277 14056
rect 13044 14016 13050 14028
rect 13265 14025 13277 14028
rect 13311 14025 13323 14059
rect 23474 14056 23480 14068
rect 23435 14028 23480 14056
rect 13265 14019 13323 14025
rect 23474 14016 23480 14028
rect 23532 14016 23538 14068
rect 3970 13948 3976 14000
rect 4028 13988 4034 14000
rect 5169 13991 5227 13997
rect 5169 13988 5181 13991
rect 4028 13960 5181 13988
rect 4028 13948 4034 13960
rect 5169 13957 5181 13960
rect 5215 13957 5227 13991
rect 5169 13951 5227 13957
rect 23845 13991 23903 13997
rect 23845 13957 23857 13991
rect 23891 13988 23903 13991
rect 24854 13988 24860 14000
rect 23891 13960 24860 13988
rect 23891 13957 23903 13960
rect 23845 13951 23903 13957
rect 24854 13948 24860 13960
rect 24912 13948 24918 14000
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13920 1915 13923
rect 1903 13892 2084 13920
rect 1903 13889 1915 13892
rect 1857 13883 1915 13889
rect 1949 13855 2007 13861
rect 1949 13821 1961 13855
rect 1995 13821 2007 13855
rect 2056 13852 2084 13892
rect 3050 13880 3056 13932
rect 3108 13920 3114 13932
rect 3697 13923 3755 13929
rect 3697 13920 3709 13923
rect 3108 13892 3709 13920
rect 3108 13880 3114 13892
rect 3697 13889 3709 13892
rect 3743 13920 3755 13923
rect 5077 13923 5135 13929
rect 3743 13892 4752 13920
rect 3743 13889 3755 13892
rect 3697 13883 3755 13889
rect 2774 13852 2780 13864
rect 2056 13824 2780 13852
rect 1949 13815 2007 13821
rect 1964 13784 1992 13815
rect 2774 13812 2780 13824
rect 2832 13852 2838 13864
rect 4724 13861 4752 13892
rect 5077 13889 5089 13923
rect 5123 13920 5135 13923
rect 5813 13923 5871 13929
rect 5813 13920 5825 13923
rect 5123 13892 5825 13920
rect 5123 13889 5135 13892
rect 5077 13883 5135 13889
rect 5813 13889 5825 13892
rect 5859 13920 5871 13923
rect 6546 13920 6552 13932
rect 5859 13892 6552 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 6546 13880 6552 13892
rect 6604 13880 6610 13932
rect 9585 13923 9643 13929
rect 9585 13889 9597 13923
rect 9631 13920 9643 13923
rect 10597 13923 10655 13929
rect 10597 13920 10609 13923
rect 9631 13892 10609 13920
rect 9631 13889 9643 13892
rect 9585 13883 9643 13889
rect 10597 13889 10609 13892
rect 10643 13920 10655 13923
rect 10686 13920 10692 13932
rect 10643 13892 10692 13920
rect 10643 13889 10655 13892
rect 10597 13883 10655 13889
rect 10686 13880 10692 13892
rect 10744 13880 10750 13932
rect 4709 13855 4767 13861
rect 2832 13824 4108 13852
rect 2832 13812 2838 13824
rect 2216 13787 2274 13793
rect 1964 13756 2053 13784
rect 1762 13676 1768 13728
rect 1820 13716 1826 13728
rect 2025 13716 2053 13756
rect 2216 13753 2228 13787
rect 2262 13784 2274 13787
rect 3050 13784 3056 13796
rect 2262 13756 3056 13784
rect 2262 13753 2274 13756
rect 2216 13747 2274 13753
rect 3050 13744 3056 13756
rect 3108 13784 3114 13796
rect 3234 13784 3240 13796
rect 3108 13756 3240 13784
rect 3108 13744 3114 13756
rect 3234 13744 3240 13756
rect 3292 13744 3298 13796
rect 4080 13784 4108 13824
rect 4709 13821 4721 13855
rect 4755 13852 4767 13855
rect 5258 13852 5264 13864
rect 4755 13824 5264 13852
rect 4755 13821 4767 13824
rect 4709 13815 4767 13821
rect 5258 13812 5264 13824
rect 5316 13852 5322 13864
rect 5316 13824 5764 13852
rect 5316 13812 5322 13824
rect 4157 13787 4215 13793
rect 4157 13784 4169 13787
rect 4080 13756 4169 13784
rect 4157 13753 4169 13756
rect 4203 13753 4215 13787
rect 4157 13747 4215 13753
rect 5442 13744 5448 13796
rect 5500 13784 5506 13796
rect 5629 13787 5687 13793
rect 5629 13784 5641 13787
rect 5500 13756 5641 13784
rect 5500 13744 5506 13756
rect 5629 13753 5641 13756
rect 5675 13753 5687 13787
rect 5736 13784 5764 13824
rect 6914 13812 6920 13864
rect 6972 13852 6978 13864
rect 7285 13855 7343 13861
rect 7285 13852 7297 13855
rect 6972 13824 7297 13852
rect 6972 13812 6978 13824
rect 7285 13821 7297 13824
rect 7331 13821 7343 13855
rect 7742 13852 7748 13864
rect 7703 13824 7748 13852
rect 7285 13815 7343 13821
rect 7742 13812 7748 13824
rect 7800 13812 7806 13864
rect 7834 13812 7840 13864
rect 7892 13852 7898 13864
rect 8110 13861 8116 13864
rect 8104 13852 8116 13861
rect 7892 13824 7937 13852
rect 8071 13824 8116 13852
rect 7892 13812 7898 13824
rect 8104 13815 8116 13824
rect 8110 13812 8116 13815
rect 8168 13812 8174 13864
rect 12894 13852 12900 13864
rect 12855 13824 12900 13852
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 23658 13852 23664 13864
rect 23619 13824 23664 13852
rect 23658 13812 23664 13824
rect 23716 13852 23722 13864
rect 24213 13855 24271 13861
rect 24213 13852 24225 13855
rect 23716 13824 24225 13852
rect 23716 13812 23722 13824
rect 24213 13821 24225 13824
rect 24259 13821 24271 13855
rect 24213 13815 24271 13821
rect 6730 13784 6736 13796
rect 5736 13756 6736 13784
rect 5629 13747 5687 13753
rect 6730 13744 6736 13756
rect 6788 13744 6794 13796
rect 9861 13787 9919 13793
rect 9861 13753 9873 13787
rect 9907 13784 9919 13787
rect 10505 13787 10563 13793
rect 10505 13784 10517 13787
rect 9907 13756 10517 13784
rect 9907 13753 9919 13756
rect 9861 13747 9919 13753
rect 10505 13753 10517 13756
rect 10551 13784 10563 13787
rect 11698 13784 11704 13796
rect 10551 13756 11704 13784
rect 10551 13753 10563 13756
rect 10505 13747 10563 13753
rect 11698 13744 11704 13756
rect 11756 13744 11762 13796
rect 2590 13716 2596 13728
rect 1820 13688 2596 13716
rect 1820 13676 1826 13688
rect 2590 13676 2596 13688
rect 2648 13676 2654 13728
rect 5537 13719 5595 13725
rect 5537 13685 5549 13719
rect 5583 13716 5595 13719
rect 6270 13716 6276 13728
rect 5583 13688 6276 13716
rect 5583 13685 5595 13688
rect 5537 13679 5595 13685
rect 6270 13676 6276 13688
rect 6328 13676 6334 13728
rect 6822 13716 6828 13728
rect 6783 13688 6828 13716
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 8110 13676 8116 13728
rect 8168 13716 8174 13728
rect 9217 13719 9275 13725
rect 9217 13716 9229 13719
rect 8168 13688 9229 13716
rect 8168 13676 8174 13688
rect 9217 13685 9229 13688
rect 9263 13685 9275 13719
rect 9217 13679 9275 13685
rect 9950 13676 9956 13728
rect 10008 13716 10014 13728
rect 10413 13719 10471 13725
rect 10413 13716 10425 13719
rect 10008 13688 10425 13716
rect 10008 13676 10014 13688
rect 10413 13685 10425 13688
rect 10459 13685 10471 13719
rect 11146 13716 11152 13728
rect 11107 13688 11152 13716
rect 10413 13679 10471 13685
rect 11146 13676 11152 13688
rect 11204 13676 11210 13728
rect 11517 13719 11575 13725
rect 11517 13685 11529 13719
rect 11563 13716 11575 13719
rect 11882 13716 11888 13728
rect 11563 13688 11888 13716
rect 11563 13685 11575 13688
rect 11517 13679 11575 13685
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 12492 13688 12537 13716
rect 12492 13676 12498 13688
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 3050 13472 3056 13524
rect 3108 13512 3114 13524
rect 3145 13515 3203 13521
rect 3145 13512 3157 13515
rect 3108 13484 3157 13512
rect 3108 13472 3114 13484
rect 3145 13481 3157 13484
rect 3191 13481 3203 13515
rect 3145 13475 3203 13481
rect 3878 13472 3884 13524
rect 3936 13512 3942 13524
rect 4249 13515 4307 13521
rect 4249 13512 4261 13515
rect 3936 13484 4261 13512
rect 3936 13472 3942 13484
rect 4249 13481 4261 13484
rect 4295 13481 4307 13515
rect 4249 13475 4307 13481
rect 5261 13515 5319 13521
rect 5261 13481 5273 13515
rect 5307 13512 5319 13515
rect 5442 13512 5448 13524
rect 5307 13484 5448 13512
rect 5307 13481 5319 13484
rect 5261 13475 5319 13481
rect 5442 13472 5448 13484
rect 5500 13512 5506 13524
rect 7561 13515 7619 13521
rect 7561 13512 7573 13515
rect 5500 13484 7573 13512
rect 5500 13472 5506 13484
rect 7561 13481 7573 13484
rect 7607 13481 7619 13515
rect 7561 13475 7619 13481
rect 8849 13515 8907 13521
rect 8849 13481 8861 13515
rect 8895 13512 8907 13515
rect 9125 13515 9183 13521
rect 9125 13512 9137 13515
rect 8895 13484 9137 13512
rect 8895 13481 8907 13484
rect 8849 13475 8907 13481
rect 9125 13481 9137 13484
rect 9171 13512 9183 13515
rect 9306 13512 9312 13524
rect 9171 13484 9312 13512
rect 9171 13481 9183 13484
rect 9125 13475 9183 13481
rect 9306 13472 9312 13484
rect 9364 13472 9370 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10045 13515 10103 13521
rect 10045 13512 10057 13515
rect 10008 13484 10057 13512
rect 10008 13472 10014 13484
rect 10045 13481 10057 13484
rect 10091 13481 10103 13515
rect 10045 13475 10103 13481
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 11609 13515 11667 13521
rect 11609 13512 11621 13515
rect 11204 13484 11621 13512
rect 11204 13472 11210 13484
rect 11609 13481 11621 13484
rect 11655 13481 11667 13515
rect 11882 13512 11888 13524
rect 11843 13484 11888 13512
rect 11609 13475 11667 13481
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 1946 13404 1952 13456
rect 2004 13453 2010 13456
rect 2004 13447 2068 13453
rect 2004 13413 2022 13447
rect 2056 13444 2068 13447
rect 3234 13444 3240 13456
rect 2056 13416 3240 13444
rect 2056 13413 2068 13416
rect 2004 13407 2068 13413
rect 2004 13404 2010 13407
rect 3234 13404 3240 13416
rect 3292 13444 3298 13456
rect 3421 13447 3479 13453
rect 3421 13444 3433 13447
rect 3292 13416 3433 13444
rect 3292 13404 3298 13416
rect 3421 13413 3433 13416
rect 3467 13413 3479 13447
rect 6362 13444 6368 13456
rect 3421 13407 3479 13413
rect 5368 13416 6368 13444
rect 1762 13376 1768 13388
rect 1723 13348 1768 13376
rect 1762 13336 1768 13348
rect 1820 13336 1826 13388
rect 2498 13336 2504 13388
rect 2556 13376 2562 13388
rect 4062 13376 4068 13388
rect 2556 13348 4068 13376
rect 2556 13336 2562 13348
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 3602 13268 3608 13320
rect 3660 13308 3666 13320
rect 3878 13308 3884 13320
rect 3660 13280 3884 13308
rect 3660 13268 3666 13280
rect 3878 13268 3884 13280
rect 3936 13268 3942 13320
rect 5258 13268 5264 13320
rect 5316 13308 5322 13320
rect 5368 13317 5396 13416
rect 6362 13404 6368 13416
rect 6420 13404 6426 13456
rect 10496 13447 10554 13453
rect 10496 13413 10508 13447
rect 10542 13444 10554 13447
rect 10686 13444 10692 13456
rect 10542 13416 10692 13444
rect 10542 13413 10554 13416
rect 10496 13407 10554 13413
rect 10686 13404 10692 13416
rect 10744 13404 10750 13456
rect 5620 13379 5678 13385
rect 5620 13345 5632 13379
rect 5666 13376 5678 13379
rect 5994 13376 6000 13388
rect 5666 13348 6000 13376
rect 5666 13345 5678 13348
rect 5620 13339 5678 13345
rect 5994 13336 6000 13348
rect 6052 13336 6058 13388
rect 7929 13379 7987 13385
rect 7929 13345 7941 13379
rect 7975 13376 7987 13379
rect 8570 13376 8576 13388
rect 7975 13348 8576 13376
rect 7975 13345 7987 13348
rect 7929 13339 7987 13345
rect 8570 13336 8576 13348
rect 8628 13336 8634 13388
rect 9306 13376 9312 13388
rect 9267 13348 9312 13376
rect 9306 13336 9312 13348
rect 9364 13336 9370 13388
rect 10134 13336 10140 13388
rect 10192 13376 10198 13388
rect 10229 13379 10287 13385
rect 10229 13376 10241 13379
rect 10192 13348 10241 13376
rect 10192 13336 10198 13348
rect 10229 13345 10241 13348
rect 10275 13345 10287 13379
rect 22278 13376 22284 13388
rect 22239 13348 22284 13376
rect 10229 13339 10287 13345
rect 22278 13336 22284 13348
rect 22336 13336 22342 13388
rect 5353 13311 5411 13317
rect 5353 13308 5365 13311
rect 5316 13280 5365 13308
rect 5316 13268 5322 13280
rect 5353 13277 5365 13280
rect 5399 13277 5411 13311
rect 5353 13271 5411 13277
rect 7650 13268 7656 13320
rect 7708 13308 7714 13320
rect 8021 13311 8079 13317
rect 8021 13308 8033 13311
rect 7708 13280 8033 13308
rect 7708 13268 7714 13280
rect 8021 13277 8033 13280
rect 8067 13277 8079 13311
rect 8202 13308 8208 13320
rect 8163 13280 8208 13308
rect 8021 13271 8079 13277
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 6730 13240 6736 13252
rect 6691 13212 6736 13240
rect 6730 13200 6736 13212
rect 6788 13200 6794 13252
rect 1673 13175 1731 13181
rect 1673 13141 1685 13175
rect 1719 13172 1731 13175
rect 1762 13172 1768 13184
rect 1719 13144 1768 13172
rect 1719 13141 1731 13144
rect 1673 13135 1731 13141
rect 1762 13132 1768 13144
rect 1820 13132 1826 13184
rect 4709 13175 4767 13181
rect 4709 13141 4721 13175
rect 4755 13172 4767 13175
rect 4798 13172 4804 13184
rect 4755 13144 4804 13172
rect 4755 13141 4767 13144
rect 4709 13135 4767 13141
rect 4798 13132 4804 13144
rect 4856 13132 4862 13184
rect 7193 13175 7251 13181
rect 7193 13141 7205 13175
rect 7239 13172 7251 13175
rect 7374 13172 7380 13184
rect 7239 13144 7380 13172
rect 7239 13141 7251 13144
rect 7193 13135 7251 13141
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 11974 13132 11980 13184
rect 12032 13172 12038 13184
rect 12345 13175 12403 13181
rect 12345 13172 12357 13175
rect 12032 13144 12357 13172
rect 12032 13132 12038 13144
rect 12345 13141 12357 13144
rect 12391 13172 12403 13175
rect 12621 13175 12679 13181
rect 12621 13172 12633 13175
rect 12391 13144 12633 13172
rect 12391 13141 12403 13144
rect 12345 13135 12403 13141
rect 12621 13141 12633 13144
rect 12667 13141 12679 13175
rect 12621 13135 12679 13141
rect 22465 13175 22523 13181
rect 22465 13141 22477 13175
rect 22511 13172 22523 13175
rect 23474 13172 23480 13184
rect 22511 13144 23480 13172
rect 22511 13141 22523 13144
rect 22465 13135 22523 13141
rect 23474 13132 23480 13144
rect 23532 13132 23538 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 2314 12928 2320 12980
rect 2372 12968 2378 12980
rect 2501 12971 2559 12977
rect 2501 12968 2513 12971
rect 2372 12940 2513 12968
rect 2372 12928 2378 12940
rect 2501 12937 2513 12940
rect 2547 12937 2559 12971
rect 2501 12931 2559 12937
rect 3694 12928 3700 12980
rect 3752 12968 3758 12980
rect 3752 12940 4016 12968
rect 3752 12928 3758 12940
rect 3988 12900 4016 12940
rect 4062 12928 4068 12980
rect 4120 12968 4126 12980
rect 4709 12971 4767 12977
rect 4709 12968 4721 12971
rect 4120 12940 4721 12968
rect 4120 12928 4126 12940
rect 4709 12937 4721 12940
rect 4755 12937 4767 12971
rect 10134 12968 10140 12980
rect 4709 12931 4767 12937
rect 9784 12940 10140 12968
rect 5445 12903 5503 12909
rect 5445 12900 5457 12903
rect 3988 12872 5457 12900
rect 5445 12869 5457 12872
rect 5491 12869 5503 12903
rect 8570 12900 8576 12912
rect 8531 12872 8576 12900
rect 5445 12863 5503 12869
rect 8570 12860 8576 12872
rect 8628 12860 8634 12912
rect 9784 12844 9812 12940
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 10686 12928 10692 12980
rect 10744 12968 10750 12980
rect 11149 12971 11207 12977
rect 11149 12968 11161 12971
rect 10744 12940 11161 12968
rect 10744 12928 10750 12940
rect 11149 12937 11161 12940
rect 11195 12968 11207 12971
rect 11425 12971 11483 12977
rect 11425 12968 11437 12971
rect 11195 12940 11437 12968
rect 11195 12937 11207 12940
rect 11149 12931 11207 12937
rect 11425 12937 11437 12940
rect 11471 12937 11483 12971
rect 11974 12968 11980 12980
rect 11935 12940 11980 12968
rect 11425 12931 11483 12937
rect 11974 12928 11980 12940
rect 12032 12928 12038 12980
rect 11882 12900 11888 12912
rect 11843 12872 11888 12900
rect 11882 12860 11888 12872
rect 11940 12860 11946 12912
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12832 2191 12835
rect 2866 12832 2872 12844
rect 2179 12804 2872 12832
rect 2179 12801 2191 12804
rect 2133 12795 2191 12801
rect 2866 12792 2872 12804
rect 2924 12792 2930 12844
rect 7466 12792 7472 12844
rect 7524 12832 7530 12844
rect 7653 12835 7711 12841
rect 7653 12832 7665 12835
rect 7524 12804 7665 12832
rect 7524 12792 7530 12804
rect 7653 12801 7665 12804
rect 7699 12801 7711 12835
rect 9766 12832 9772 12844
rect 9679 12804 9772 12832
rect 7653 12795 7711 12801
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 1854 12724 1860 12776
rect 1912 12764 1918 12776
rect 1949 12767 2007 12773
rect 1949 12764 1961 12767
rect 1912 12736 1961 12764
rect 1912 12724 1918 12736
rect 1949 12733 1961 12736
rect 1995 12733 2007 12767
rect 1949 12727 2007 12733
rect 2590 12724 2596 12776
rect 2648 12764 2654 12776
rect 3326 12773 3332 12776
rect 3053 12767 3111 12773
rect 3053 12764 3065 12767
rect 2648 12736 3065 12764
rect 2648 12724 2654 12736
rect 3053 12733 3065 12736
rect 3099 12733 3111 12767
rect 3320 12764 3332 12773
rect 3287 12736 3332 12764
rect 3053 12727 3111 12733
rect 3320 12727 3332 12736
rect 3068 12696 3096 12727
rect 3326 12724 3332 12727
rect 3384 12724 3390 12776
rect 5261 12767 5319 12773
rect 5261 12764 5273 12767
rect 5092 12736 5273 12764
rect 4338 12696 4344 12708
rect 3068 12668 4344 12696
rect 4338 12656 4344 12668
rect 4396 12656 4402 12708
rect 5092 12640 5120 12736
rect 5261 12733 5273 12736
rect 5307 12733 5319 12767
rect 12158 12764 12164 12776
rect 12071 12736 12164 12764
rect 5261 12727 5319 12733
rect 12158 12724 12164 12736
rect 12216 12764 12222 12776
rect 12621 12767 12679 12773
rect 12621 12764 12633 12767
rect 12216 12736 12633 12764
rect 12216 12724 12222 12736
rect 12621 12733 12633 12736
rect 12667 12733 12679 12767
rect 12986 12764 12992 12776
rect 12947 12736 12992 12764
rect 12621 12727 12679 12733
rect 12986 12724 12992 12736
rect 13044 12724 13050 12776
rect 22278 12764 22284 12776
rect 22239 12736 22284 12764
rect 22278 12724 22284 12736
rect 22336 12724 22342 12776
rect 5534 12656 5540 12708
rect 5592 12696 5598 12708
rect 6181 12699 6239 12705
rect 6181 12696 6193 12699
rect 5592 12668 6193 12696
rect 5592 12656 5598 12668
rect 6181 12665 6193 12668
rect 6227 12665 6239 12699
rect 6181 12659 6239 12665
rect 6641 12699 6699 12705
rect 6641 12665 6653 12699
rect 6687 12696 6699 12699
rect 7469 12699 7527 12705
rect 7469 12696 7481 12699
rect 6687 12668 7481 12696
rect 6687 12665 6699 12668
rect 6641 12659 6699 12665
rect 7469 12665 7481 12668
rect 7515 12696 7527 12699
rect 8386 12696 8392 12708
rect 7515 12668 8392 12696
rect 7515 12665 7527 12668
rect 7469 12659 7527 12665
rect 8386 12656 8392 12668
rect 8444 12656 8450 12708
rect 8662 12656 8668 12708
rect 8720 12696 8726 12708
rect 9217 12699 9275 12705
rect 9217 12696 9229 12699
rect 8720 12668 9229 12696
rect 8720 12656 8726 12668
rect 9217 12665 9229 12668
rect 9263 12696 9275 12699
rect 9306 12696 9312 12708
rect 9263 12668 9312 12696
rect 9263 12665 9275 12668
rect 9217 12659 9275 12665
rect 9306 12656 9312 12668
rect 9364 12656 9370 12708
rect 9674 12656 9680 12708
rect 9732 12696 9738 12708
rect 10042 12705 10048 12708
rect 10036 12696 10048 12705
rect 9732 12668 10048 12696
rect 9732 12656 9738 12668
rect 10036 12659 10048 12668
rect 10042 12656 10048 12659
rect 10100 12656 10106 12708
rect 11882 12656 11888 12708
rect 11940 12696 11946 12708
rect 13004 12696 13032 12724
rect 11940 12668 13032 12696
rect 11940 12656 11946 12668
rect 1486 12628 1492 12640
rect 1447 12600 1492 12628
rect 1486 12588 1492 12600
rect 1544 12588 1550 12640
rect 1857 12631 1915 12637
rect 1857 12597 1869 12631
rect 1903 12628 1915 12631
rect 2314 12628 2320 12640
rect 1903 12600 2320 12628
rect 1903 12597 1915 12600
rect 1857 12591 1915 12597
rect 2314 12588 2320 12600
rect 2372 12628 2378 12640
rect 3418 12628 3424 12640
rect 2372 12600 3424 12628
rect 2372 12588 2378 12600
rect 3418 12588 3424 12600
rect 3476 12588 3482 12640
rect 4433 12631 4491 12637
rect 4433 12597 4445 12631
rect 4479 12628 4491 12631
rect 4706 12628 4712 12640
rect 4479 12600 4712 12628
rect 4479 12597 4491 12600
rect 4433 12591 4491 12597
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 5074 12628 5080 12640
rect 5035 12600 5080 12628
rect 5074 12588 5080 12600
rect 5132 12588 5138 12640
rect 5905 12631 5963 12637
rect 5905 12597 5917 12631
rect 5951 12628 5963 12631
rect 5994 12628 6000 12640
rect 5951 12600 6000 12628
rect 5951 12597 5963 12600
rect 5905 12591 5963 12597
rect 5994 12588 6000 12600
rect 6052 12628 6058 12640
rect 6730 12628 6736 12640
rect 6052 12600 6736 12628
rect 6052 12588 6058 12600
rect 6730 12588 6736 12600
rect 6788 12588 6794 12640
rect 7098 12628 7104 12640
rect 7059 12600 7104 12628
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 7374 12588 7380 12640
rect 7432 12628 7438 12640
rect 7561 12631 7619 12637
rect 7561 12628 7573 12631
rect 7432 12600 7573 12628
rect 7432 12588 7438 12600
rect 7561 12597 7573 12600
rect 7607 12597 7619 12631
rect 8202 12628 8208 12640
rect 8163 12600 8208 12628
rect 7561 12591 7619 12597
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 8754 12628 8760 12640
rect 8715 12600 8760 12628
rect 8754 12588 8760 12600
rect 8812 12588 8818 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 3326 12384 3332 12436
rect 3384 12424 3390 12436
rect 3421 12427 3479 12433
rect 3421 12424 3433 12427
rect 3384 12396 3433 12424
rect 3384 12384 3390 12396
rect 3421 12393 3433 12396
rect 3467 12393 3479 12427
rect 3421 12387 3479 12393
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4249 12427 4307 12433
rect 4249 12424 4261 12427
rect 4212 12396 4261 12424
rect 4212 12384 4218 12396
rect 4249 12393 4261 12396
rect 4295 12393 4307 12427
rect 4249 12387 4307 12393
rect 4338 12384 4344 12436
rect 4396 12424 4402 12436
rect 5169 12427 5227 12433
rect 5169 12424 5181 12427
rect 4396 12396 5181 12424
rect 4396 12384 4402 12396
rect 5169 12393 5181 12396
rect 5215 12424 5227 12427
rect 5258 12424 5264 12436
rect 5215 12396 5264 12424
rect 5215 12393 5227 12396
rect 5169 12387 5227 12393
rect 5258 12384 5264 12396
rect 5316 12424 5322 12436
rect 5316 12396 5580 12424
rect 5316 12384 5322 12396
rect 1857 12291 1915 12297
rect 1857 12257 1869 12291
rect 1903 12288 1915 12291
rect 2314 12288 2320 12300
rect 1903 12260 2320 12288
rect 1903 12257 1915 12260
rect 1857 12251 1915 12257
rect 2314 12248 2320 12260
rect 2372 12248 2378 12300
rect 4065 12291 4123 12297
rect 4065 12257 4077 12291
rect 4111 12288 4123 12291
rect 4338 12288 4344 12300
rect 4111 12260 4344 12288
rect 4111 12257 4123 12260
rect 4065 12251 4123 12257
rect 4338 12248 4344 12260
rect 4396 12248 4402 12300
rect 5258 12248 5264 12300
rect 5316 12288 5322 12300
rect 5353 12291 5411 12297
rect 5353 12288 5365 12291
rect 5316 12260 5365 12288
rect 5316 12248 5322 12260
rect 5353 12257 5365 12260
rect 5399 12257 5411 12291
rect 5353 12251 5411 12257
rect 5552 12232 5580 12396
rect 6822 12384 6828 12436
rect 6880 12424 6886 12436
rect 6917 12427 6975 12433
rect 6917 12424 6929 12427
rect 6880 12396 6929 12424
rect 6880 12384 6886 12396
rect 6917 12393 6929 12396
rect 6963 12424 6975 12427
rect 7006 12424 7012 12436
rect 6963 12396 7012 12424
rect 6963 12393 6975 12396
rect 6917 12387 6975 12393
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 7285 12427 7343 12433
rect 7285 12393 7297 12427
rect 7331 12424 7343 12427
rect 7466 12424 7472 12436
rect 7331 12396 7472 12424
rect 7331 12393 7343 12396
rect 7285 12387 7343 12393
rect 7466 12384 7472 12396
rect 7524 12384 7530 12436
rect 7926 12384 7932 12436
rect 7984 12424 7990 12436
rect 8021 12427 8079 12433
rect 8021 12424 8033 12427
rect 7984 12396 8033 12424
rect 7984 12384 7990 12396
rect 8021 12393 8033 12396
rect 8067 12393 8079 12427
rect 8021 12387 8079 12393
rect 8389 12427 8447 12433
rect 8389 12393 8401 12427
rect 8435 12424 8447 12427
rect 8754 12424 8760 12436
rect 8435 12396 8760 12424
rect 8435 12393 8447 12396
rect 8389 12387 8447 12393
rect 8754 12384 8760 12396
rect 8812 12384 8818 12436
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 11057 12427 11115 12433
rect 11057 12424 11069 12427
rect 10100 12396 11069 12424
rect 10100 12384 10106 12396
rect 11057 12393 11069 12396
rect 11103 12393 11115 12427
rect 11057 12387 11115 12393
rect 9493 12359 9551 12365
rect 9493 12325 9505 12359
rect 9539 12356 9551 12359
rect 9944 12359 10002 12365
rect 9944 12356 9956 12359
rect 9539 12328 9956 12356
rect 9539 12325 9551 12328
rect 9493 12319 9551 12325
rect 9944 12325 9956 12328
rect 9990 12356 10002 12359
rect 10594 12356 10600 12368
rect 9990 12328 10600 12356
rect 9990 12325 10002 12328
rect 9944 12319 10002 12325
rect 10594 12316 10600 12328
rect 10652 12316 10658 12368
rect 5804 12291 5862 12297
rect 5804 12257 5816 12291
rect 5850 12288 5862 12291
rect 6086 12288 6092 12300
rect 5850 12260 6092 12288
rect 5850 12257 5862 12260
rect 5804 12251 5862 12257
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 9677 12291 9735 12297
rect 9677 12257 9689 12291
rect 9723 12288 9735 12291
rect 9766 12288 9772 12300
rect 9723 12260 9772 12288
rect 9723 12257 9735 12260
rect 9677 12251 9735 12257
rect 9766 12248 9772 12260
rect 9824 12248 9830 12300
rect 11606 12248 11612 12300
rect 11664 12288 11670 12300
rect 11701 12291 11759 12297
rect 11701 12288 11713 12291
rect 11664 12260 11713 12288
rect 11664 12248 11670 12260
rect 11701 12257 11713 12260
rect 11747 12257 11759 12291
rect 11701 12251 11759 12257
rect 12244 12291 12302 12297
rect 12244 12257 12256 12291
rect 12290 12288 12302 12291
rect 12710 12288 12716 12300
rect 12290 12260 12716 12288
rect 12290 12257 12302 12260
rect 12244 12251 12302 12257
rect 12710 12248 12716 12260
rect 12768 12248 12774 12300
rect 21726 12288 21732 12300
rect 21687 12260 21732 12288
rect 21726 12248 21732 12260
rect 21784 12248 21790 12300
rect 1949 12223 2007 12229
rect 1949 12189 1961 12223
rect 1995 12189 2007 12223
rect 1949 12183 2007 12189
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 3050 12220 3056 12232
rect 2179 12192 3056 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 1964 12152 1992 12183
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 5534 12220 5540 12232
rect 5495 12192 5540 12220
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 8478 12220 8484 12232
rect 8439 12192 8484 12220
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 8665 12223 8723 12229
rect 8665 12189 8677 12223
rect 8711 12189 8723 12223
rect 9122 12220 9128 12232
rect 9083 12192 9128 12220
rect 8665 12183 8723 12189
rect 1964 12124 3924 12152
rect 3896 12096 3924 12124
rect 7742 12112 7748 12164
rect 7800 12152 7806 12164
rect 8680 12152 8708 12183
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 10686 12180 10692 12232
rect 10744 12220 10750 12232
rect 11974 12220 11980 12232
rect 10744 12192 11980 12220
rect 10744 12180 10750 12192
rect 11974 12180 11980 12192
rect 12032 12180 12038 12232
rect 7800 12124 9720 12152
rect 7800 12112 7806 12124
rect 9692 12096 9720 12124
rect 1489 12087 1547 12093
rect 1489 12053 1501 12087
rect 1535 12084 1547 12087
rect 1946 12084 1952 12096
rect 1535 12056 1952 12084
rect 1535 12053 1547 12056
rect 1489 12047 1547 12053
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 2777 12087 2835 12093
rect 2777 12053 2789 12087
rect 2823 12084 2835 12087
rect 2958 12084 2964 12096
rect 2823 12056 2964 12084
rect 2823 12053 2835 12056
rect 2777 12047 2835 12053
rect 2958 12044 2964 12056
rect 3016 12044 3022 12096
rect 3878 12084 3884 12096
rect 3839 12056 3884 12084
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 4338 12044 4344 12096
rect 4396 12084 4402 12096
rect 4617 12087 4675 12093
rect 4617 12084 4629 12087
rect 4396 12056 4629 12084
rect 4396 12044 4402 12056
rect 4617 12053 4629 12056
rect 4663 12053 4675 12087
rect 4617 12047 4675 12053
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 5077 12087 5135 12093
rect 5077 12084 5089 12087
rect 4856 12056 5089 12084
rect 4856 12044 4862 12056
rect 5077 12053 5089 12056
rect 5123 12084 5135 12087
rect 5166 12084 5172 12096
rect 5123 12056 5172 12084
rect 5123 12053 5135 12056
rect 5077 12047 5135 12053
rect 5166 12044 5172 12056
rect 5224 12044 5230 12096
rect 7650 12084 7656 12096
rect 7611 12056 7656 12084
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 9674 12044 9680 12096
rect 9732 12044 9738 12096
rect 11146 12044 11152 12096
rect 11204 12084 11210 12096
rect 11333 12087 11391 12093
rect 11333 12084 11345 12087
rect 11204 12056 11345 12084
rect 11204 12044 11210 12056
rect 11333 12053 11345 12056
rect 11379 12053 11391 12087
rect 11333 12047 11391 12053
rect 13262 12044 13268 12096
rect 13320 12084 13326 12096
rect 13357 12087 13415 12093
rect 13357 12084 13369 12087
rect 13320 12056 13369 12084
rect 13320 12044 13326 12056
rect 13357 12053 13369 12056
rect 13403 12053 13415 12087
rect 21910 12084 21916 12096
rect 21871 12056 21916 12084
rect 13357 12047 13415 12053
rect 21910 12044 21916 12056
rect 21968 12044 21974 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 2685 11883 2743 11889
rect 2685 11880 2697 11883
rect 2464 11852 2697 11880
rect 2464 11840 2470 11852
rect 2685 11849 2697 11852
rect 2731 11849 2743 11883
rect 2685 11843 2743 11849
rect 3510 11840 3516 11892
rect 3568 11880 3574 11892
rect 4341 11883 4399 11889
rect 4341 11880 4353 11883
rect 3568 11852 4353 11880
rect 3568 11840 3574 11852
rect 4341 11849 4353 11852
rect 4387 11849 4399 11883
rect 4341 11843 4399 11849
rect 5905 11883 5963 11889
rect 5905 11849 5917 11883
rect 5951 11880 5963 11883
rect 5994 11880 6000 11892
rect 5951 11852 6000 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 1670 11744 1676 11756
rect 1631 11716 1676 11744
rect 1670 11704 1676 11716
rect 1728 11704 1734 11756
rect 3234 11744 3240 11756
rect 3195 11716 3240 11744
rect 3234 11704 3240 11716
rect 3292 11744 3298 11756
rect 3697 11747 3755 11753
rect 3697 11744 3709 11747
rect 3292 11716 3709 11744
rect 3292 11704 3298 11716
rect 3697 11713 3709 11716
rect 3743 11713 3755 11747
rect 4356 11744 4384 11843
rect 5994 11840 6000 11852
rect 6052 11880 6058 11892
rect 6638 11880 6644 11892
rect 6052 11852 6644 11880
rect 6052 11840 6058 11852
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 7742 11880 7748 11892
rect 7703 11852 7748 11880
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 8113 11883 8171 11889
rect 8113 11849 8125 11883
rect 8159 11880 8171 11883
rect 8754 11880 8760 11892
rect 8159 11852 8760 11880
rect 8159 11849 8171 11852
rect 8113 11843 8171 11849
rect 8754 11840 8760 11852
rect 8812 11840 8818 11892
rect 11974 11840 11980 11892
rect 12032 11880 12038 11892
rect 13357 11883 13415 11889
rect 13357 11880 13369 11883
rect 12032 11852 13369 11880
rect 12032 11840 12038 11852
rect 13357 11849 13369 11852
rect 13403 11880 13415 11883
rect 13725 11883 13783 11889
rect 13725 11880 13737 11883
rect 13403 11852 13737 11880
rect 13403 11849 13415 11852
rect 13357 11843 13415 11849
rect 13725 11849 13737 11852
rect 13771 11880 13783 11883
rect 14093 11883 14151 11889
rect 14093 11880 14105 11883
rect 13771 11852 14105 11880
rect 13771 11849 13783 11852
rect 13725 11843 13783 11849
rect 14093 11849 14105 11852
rect 14139 11849 14151 11883
rect 14093 11843 14151 11849
rect 21726 11812 21732 11824
rect 21687 11784 21732 11812
rect 21726 11772 21732 11784
rect 21784 11772 21790 11824
rect 4356 11716 4660 11744
rect 3697 11707 3755 11713
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 3326 11676 3332 11688
rect 1443 11648 3332 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 3326 11636 3332 11648
rect 3384 11636 3390 11688
rect 4525 11679 4583 11685
rect 4525 11645 4537 11679
rect 4571 11645 4583 11679
rect 4632 11676 4660 11716
rect 9766 11704 9772 11756
rect 9824 11744 9830 11756
rect 10686 11744 10692 11756
rect 9824 11716 10692 11744
rect 9824 11704 9830 11716
rect 10686 11704 10692 11716
rect 10744 11704 10750 11756
rect 4781 11679 4839 11685
rect 4781 11676 4793 11679
rect 4632 11648 4793 11676
rect 4525 11639 4583 11645
rect 4781 11645 4793 11648
rect 4827 11676 4839 11679
rect 5534 11676 5540 11688
rect 4827 11648 5540 11676
rect 4827 11645 4839 11648
rect 4781 11639 4839 11645
rect 2590 11608 2596 11620
rect 2503 11580 2596 11608
rect 2590 11568 2596 11580
rect 2648 11608 2654 11620
rect 3145 11611 3203 11617
rect 3145 11608 3157 11611
rect 2648 11580 3157 11608
rect 2648 11568 2654 11580
rect 3145 11577 3157 11580
rect 3191 11577 3203 11611
rect 4540 11608 4568 11639
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 12710 11676 12716 11688
rect 12671 11648 12716 11676
rect 12710 11636 12716 11648
rect 12768 11636 12774 11688
rect 5626 11608 5632 11620
rect 4540 11580 5632 11608
rect 3145 11571 3203 11577
rect 5626 11568 5632 11580
rect 5684 11568 5690 11620
rect 6549 11611 6607 11617
rect 6549 11608 6561 11611
rect 5736 11580 6561 11608
rect 2225 11543 2283 11549
rect 2225 11509 2237 11543
rect 2271 11540 2283 11543
rect 2314 11540 2320 11552
rect 2271 11512 2320 11540
rect 2271 11509 2283 11512
rect 2225 11503 2283 11509
rect 2314 11500 2320 11512
rect 2372 11500 2378 11552
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3053 11543 3111 11549
rect 3053 11540 3065 11543
rect 3016 11512 3065 11540
rect 3016 11500 3022 11512
rect 3053 11509 3065 11512
rect 3099 11509 3111 11543
rect 3053 11503 3111 11509
rect 5166 11500 5172 11552
rect 5224 11540 5230 11552
rect 5736 11540 5764 11580
rect 6549 11577 6561 11580
rect 6595 11577 6607 11611
rect 6549 11571 6607 11577
rect 7377 11611 7435 11617
rect 7377 11577 7389 11611
rect 7423 11608 7435 11611
rect 8478 11608 8484 11620
rect 7423 11580 8484 11608
rect 7423 11577 7435 11580
rect 7377 11571 7435 11577
rect 8478 11568 8484 11580
rect 8536 11568 8542 11620
rect 8757 11611 8815 11617
rect 8757 11577 8769 11611
rect 8803 11608 8815 11611
rect 8846 11608 8852 11620
rect 8803 11580 8852 11608
rect 8803 11577 8815 11580
rect 8757 11571 8815 11577
rect 8846 11568 8852 11580
rect 8904 11568 8910 11620
rect 9214 11568 9220 11620
rect 9272 11608 9278 11620
rect 10934 11611 10992 11617
rect 10934 11608 10946 11611
rect 9272 11580 10946 11608
rect 9272 11568 9278 11580
rect 10934 11577 10946 11580
rect 10980 11608 10992 11611
rect 11146 11608 11152 11620
rect 10980 11580 11152 11608
rect 10980 11577 10992 11580
rect 10934 11571 10992 11577
rect 11146 11568 11152 11580
rect 11204 11568 11210 11620
rect 5224 11512 5764 11540
rect 5224 11500 5230 11512
rect 6086 11500 6092 11552
rect 6144 11540 6150 11552
rect 6270 11540 6276 11552
rect 6144 11512 6276 11540
rect 6144 11500 6150 11512
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 6825 11543 6883 11549
rect 6825 11509 6837 11543
rect 6871 11540 6883 11543
rect 6914 11540 6920 11552
rect 6871 11512 6920 11540
rect 6871 11509 6883 11512
rect 6825 11503 6883 11509
rect 6914 11500 6920 11512
rect 6972 11500 6978 11552
rect 10134 11540 10140 11552
rect 10095 11512 10140 11540
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 10686 11500 10692 11552
rect 10744 11540 10750 11552
rect 12069 11543 12127 11549
rect 12069 11540 12081 11543
rect 10744 11512 12081 11540
rect 10744 11500 10750 11512
rect 12069 11509 12081 11512
rect 12115 11509 12127 11543
rect 12069 11503 12127 11509
rect 12986 11500 12992 11552
rect 13044 11540 13050 11552
rect 13081 11543 13139 11549
rect 13081 11540 13093 11543
rect 13044 11512 13093 11540
rect 13044 11500 13050 11512
rect 13081 11509 13093 11512
rect 13127 11540 13139 11543
rect 13722 11540 13728 11552
rect 13127 11512 13728 11540
rect 13127 11509 13139 11512
rect 13081 11503 13139 11509
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 3053 11339 3111 11345
rect 3053 11305 3065 11339
rect 3099 11336 3111 11339
rect 3142 11336 3148 11348
rect 3099 11308 3148 11336
rect 3099 11305 3111 11308
rect 3053 11299 3111 11305
rect 3142 11296 3148 11308
rect 3200 11296 3206 11348
rect 3326 11336 3332 11348
rect 3287 11308 3332 11336
rect 3326 11296 3332 11308
rect 3384 11336 3390 11348
rect 4065 11339 4123 11345
rect 4065 11336 4077 11339
rect 3384 11308 4077 11336
rect 3384 11296 3390 11308
rect 4065 11305 4077 11308
rect 4111 11305 4123 11339
rect 5258 11336 5264 11348
rect 5219 11308 5264 11336
rect 4065 11299 4123 11305
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 6270 11296 6276 11348
rect 6328 11336 6334 11348
rect 7009 11339 7067 11345
rect 7009 11336 7021 11339
rect 6328 11308 7021 11336
rect 6328 11296 6334 11308
rect 7009 11305 7021 11308
rect 7055 11305 7067 11339
rect 7009 11299 7067 11305
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 8294 11336 8300 11348
rect 7156 11308 8300 11336
rect 7156 11296 7162 11308
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 8478 11296 8484 11348
rect 8536 11336 8542 11348
rect 9677 11339 9735 11345
rect 9677 11336 9689 11339
rect 8536 11308 9689 11336
rect 8536 11296 8542 11308
rect 9677 11305 9689 11308
rect 9723 11305 9735 11339
rect 11238 11336 11244 11348
rect 11199 11308 11244 11336
rect 9677 11299 9735 11305
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 11606 11296 11612 11348
rect 11664 11336 11670 11348
rect 11701 11339 11759 11345
rect 11701 11336 11713 11339
rect 11664 11308 11713 11336
rect 11664 11296 11670 11308
rect 11701 11305 11713 11308
rect 11747 11305 11759 11339
rect 12802 11336 12808 11348
rect 12763 11308 12808 11336
rect 11701 11299 11759 11305
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 2498 11268 2504 11280
rect 1688 11240 2504 11268
rect 1688 11209 1716 11240
rect 2498 11228 2504 11240
rect 2556 11228 2562 11280
rect 5896 11271 5954 11277
rect 5896 11237 5908 11271
rect 5942 11268 5954 11271
rect 5994 11268 6000 11280
rect 5942 11240 6000 11268
rect 5942 11237 5954 11240
rect 5896 11231 5954 11237
rect 5994 11228 6000 11240
rect 6052 11228 6058 11280
rect 8110 11277 8116 11280
rect 7745 11271 7803 11277
rect 7745 11237 7757 11271
rect 7791 11268 7803 11271
rect 8104 11268 8116 11277
rect 7791 11240 8116 11268
rect 7791 11237 7803 11240
rect 7745 11231 7803 11237
rect 8104 11231 8116 11240
rect 8110 11228 8116 11231
rect 8168 11228 8174 11280
rect 1673 11203 1731 11209
rect 1673 11169 1685 11203
rect 1719 11169 1731 11203
rect 1673 11163 1731 11169
rect 1762 11160 1768 11212
rect 1820 11200 1826 11212
rect 1929 11203 1987 11209
rect 1929 11200 1941 11203
rect 1820 11172 1941 11200
rect 1820 11160 1826 11172
rect 1929 11169 1941 11172
rect 1975 11169 1987 11203
rect 1929 11163 1987 11169
rect 2958 11160 2964 11212
rect 3016 11200 3022 11212
rect 3142 11200 3148 11212
rect 3016 11172 3148 11200
rect 3016 11160 3022 11172
rect 3142 11160 3148 11172
rect 3200 11160 3206 11212
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4212 11172 4445 11200
rect 4212 11160 4218 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 5626 11200 5632 11212
rect 5539 11172 5632 11200
rect 4433 11163 4491 11169
rect 5626 11160 5632 11172
rect 5684 11200 5690 11212
rect 7837 11203 7895 11209
rect 5684 11172 6684 11200
rect 5684 11160 5690 11172
rect 3881 11135 3939 11141
rect 3881 11101 3893 11135
rect 3927 11132 3939 11135
rect 4062 11132 4068 11144
rect 3927 11104 4068 11132
rect 3927 11101 3939 11104
rect 3881 11095 3939 11101
rect 4062 11092 4068 11104
rect 4120 11132 4126 11144
rect 4525 11135 4583 11141
rect 4525 11132 4537 11135
rect 4120 11104 4537 11132
rect 4120 11092 4126 11104
rect 4525 11101 4537 11104
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 4614 11092 4620 11144
rect 4672 11132 4678 11144
rect 6656 11132 6684 11172
rect 7837 11169 7849 11203
rect 7883 11200 7895 11203
rect 9122 11200 9128 11212
rect 7883 11172 9128 11200
rect 7883 11169 7895 11172
rect 7837 11163 7895 11169
rect 7852 11132 7880 11163
rect 9122 11160 9128 11172
rect 9180 11160 9186 11212
rect 10042 11200 10048 11212
rect 10003 11172 10048 11200
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 11054 11200 11060 11212
rect 11015 11172 11060 11200
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 11606 11200 11612 11212
rect 11567 11172 11612 11200
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 13170 11200 13176 11212
rect 13131 11172 13176 11200
rect 13170 11160 13176 11172
rect 13228 11160 13234 11212
rect 13265 11203 13323 11209
rect 13265 11169 13277 11203
rect 13311 11200 13323 11203
rect 13446 11200 13452 11212
rect 13311 11172 13452 11200
rect 13311 11169 13323 11172
rect 13265 11163 13323 11169
rect 13446 11160 13452 11172
rect 13504 11160 13510 11212
rect 4672 11104 4717 11132
rect 6656 11104 7880 11132
rect 4672 11092 4678 11104
rect 9950 11092 9956 11144
rect 10008 11132 10014 11144
rect 10137 11135 10195 11141
rect 10137 11132 10149 11135
rect 10008 11104 10149 11132
rect 10008 11092 10014 11104
rect 10137 11101 10149 11104
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11132 10379 11135
rect 10686 11132 10692 11144
rect 10367 11104 10692 11132
rect 10367 11101 10379 11104
rect 10321 11095 10379 11101
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 11072 11132 11100 11160
rect 11793 11135 11851 11141
rect 11793 11132 11805 11135
rect 11072 11104 11805 11132
rect 11793 11101 11805 11104
rect 11839 11101 11851 11135
rect 11793 11095 11851 11101
rect 13078 11092 13084 11144
rect 13136 11132 13142 11144
rect 13357 11135 13415 11141
rect 13357 11132 13369 11135
rect 13136 11104 13369 11132
rect 13136 11092 13142 11104
rect 13357 11101 13369 11104
rect 13403 11101 13415 11135
rect 13357 11095 13415 11101
rect 9214 11064 9220 11076
rect 8772 11036 9220 11064
rect 1302 10956 1308 11008
rect 1360 10996 1366 11008
rect 3326 10996 3332 11008
rect 1360 10968 3332 10996
rect 1360 10956 1366 10968
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 7374 10996 7380 11008
rect 7335 10968 7380 10996
rect 7374 10956 7380 10968
rect 7432 10956 7438 11008
rect 8202 10956 8208 11008
rect 8260 10996 8266 11008
rect 8772 10996 8800 11036
rect 9214 11024 9220 11036
rect 9272 11024 9278 11076
rect 9766 11024 9772 11076
rect 9824 11064 9830 11076
rect 10781 11067 10839 11073
rect 10781 11064 10793 11067
rect 9824 11036 10793 11064
rect 9824 11024 9830 11036
rect 10781 11033 10793 11036
rect 10827 11064 10839 11067
rect 10962 11064 10968 11076
rect 10827 11036 10968 11064
rect 10827 11033 10839 11036
rect 10781 11027 10839 11033
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 8260 10968 8800 10996
rect 12529 10999 12587 11005
rect 8260 10956 8266 10968
rect 12529 10965 12541 10999
rect 12575 10996 12587 10999
rect 12802 10996 12808 11008
rect 12575 10968 12808 10996
rect 12575 10965 12587 10968
rect 12529 10959 12587 10965
rect 12802 10956 12808 10968
rect 12860 10956 12866 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 3050 10792 3056 10804
rect 3011 10764 3056 10792
rect 3050 10752 3056 10764
rect 3108 10752 3114 10804
rect 4157 10795 4215 10801
rect 4157 10761 4169 10795
rect 4203 10792 4215 10795
rect 4246 10792 4252 10804
rect 4203 10764 4252 10792
rect 4203 10761 4215 10764
rect 4157 10755 4215 10761
rect 4246 10752 4252 10764
rect 4304 10792 4310 10804
rect 4614 10792 4620 10804
rect 4304 10764 4620 10792
rect 4304 10752 4310 10764
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 5592 10764 5641 10792
rect 5592 10752 5598 10764
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 5994 10792 6000 10804
rect 5955 10764 6000 10792
rect 5629 10755 5687 10761
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7285 10795 7343 10801
rect 7285 10792 7297 10795
rect 6972 10764 7297 10792
rect 6972 10752 6978 10764
rect 7285 10761 7297 10764
rect 7331 10761 7343 10795
rect 7285 10755 7343 10761
rect 1394 10588 1400 10600
rect 1355 10560 1400 10588
rect 1394 10548 1400 10560
rect 1452 10548 1458 10600
rect 1664 10591 1722 10597
rect 1664 10557 1676 10591
rect 1710 10588 1722 10591
rect 2590 10588 2596 10600
rect 1710 10560 2596 10588
rect 1710 10557 1722 10560
rect 1664 10551 1722 10557
rect 2590 10548 2596 10560
rect 2648 10588 2654 10600
rect 3050 10588 3056 10600
rect 2648 10560 3056 10588
rect 2648 10548 2654 10560
rect 3050 10548 3056 10560
rect 3108 10548 3114 10600
rect 4249 10591 4307 10597
rect 4249 10557 4261 10591
rect 4295 10588 4307 10591
rect 4295 10560 5212 10588
rect 4295 10557 4307 10560
rect 4249 10551 4307 10557
rect 5184 10532 5212 10560
rect 5994 10548 6000 10600
rect 6052 10588 6058 10600
rect 6178 10588 6184 10600
rect 6052 10560 6184 10588
rect 6052 10548 6058 10560
rect 6178 10548 6184 10560
rect 6236 10548 6242 10600
rect 7300 10588 7328 10755
rect 7374 10752 7380 10804
rect 7432 10792 7438 10804
rect 7837 10795 7895 10801
rect 7837 10792 7849 10795
rect 7432 10764 7849 10792
rect 7432 10752 7438 10764
rect 7837 10761 7849 10764
rect 7883 10792 7895 10795
rect 7926 10792 7932 10804
rect 7883 10764 7932 10792
rect 7883 10761 7895 10764
rect 7837 10755 7895 10761
rect 7926 10752 7932 10764
rect 7984 10752 7990 10804
rect 8386 10752 8392 10804
rect 8444 10752 8450 10804
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 10689 10795 10747 10801
rect 10689 10792 10701 10795
rect 9732 10764 10701 10792
rect 9732 10752 9738 10764
rect 10689 10761 10701 10764
rect 10735 10761 10747 10795
rect 10689 10755 10747 10761
rect 12437 10795 12495 10801
rect 12437 10761 12449 10795
rect 12483 10792 12495 10795
rect 12526 10792 12532 10804
rect 12483 10764 12532 10792
rect 12483 10761 12495 10764
rect 12437 10755 12495 10761
rect 12526 10752 12532 10764
rect 12584 10752 12590 10804
rect 13814 10752 13820 10804
rect 13872 10792 13878 10804
rect 14185 10795 14243 10801
rect 14185 10792 14197 10795
rect 13872 10764 14197 10792
rect 13872 10752 13878 10764
rect 14185 10761 14197 10764
rect 14231 10761 14243 10795
rect 14185 10755 14243 10761
rect 7742 10724 7748 10736
rect 7655 10696 7748 10724
rect 7742 10684 7748 10696
rect 7800 10724 7806 10736
rect 8404 10724 8432 10752
rect 7800 10696 8432 10724
rect 7800 10684 7806 10696
rect 12250 10684 12256 10736
rect 12308 10724 12314 10736
rect 12308 10696 12940 10724
rect 12308 10684 12314 10696
rect 8110 10616 8116 10668
rect 8168 10656 8174 10668
rect 8389 10659 8447 10665
rect 8389 10656 8401 10659
rect 8168 10628 8401 10656
rect 8168 10616 8174 10628
rect 8389 10625 8401 10628
rect 8435 10656 8447 10659
rect 9490 10656 9496 10668
rect 8435 10628 9496 10656
rect 8435 10625 8447 10628
rect 8389 10619 8447 10625
rect 9490 10616 9496 10628
rect 9548 10656 9554 10668
rect 9677 10659 9735 10665
rect 9677 10656 9689 10659
rect 9548 10628 9689 10656
rect 9548 10616 9554 10628
rect 9677 10625 9689 10628
rect 9723 10625 9735 10659
rect 9677 10619 9735 10625
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 11241 10659 11299 10665
rect 11241 10656 11253 10659
rect 11112 10628 11253 10656
rect 11112 10616 11118 10628
rect 11241 10625 11253 10628
rect 11287 10656 11299 10659
rect 12342 10656 12348 10668
rect 11287 10628 12348 10656
rect 11287 10625 11299 10628
rect 11241 10619 11299 10625
rect 12342 10616 12348 10628
rect 12400 10616 12406 10668
rect 12912 10665 12940 10696
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10625 12955 10659
rect 13078 10656 13084 10668
rect 13039 10628 13084 10656
rect 12897 10619 12955 10625
rect 13078 10616 13084 10628
rect 13136 10656 13142 10668
rect 13817 10659 13875 10665
rect 13817 10656 13829 10659
rect 13136 10628 13829 10656
rect 13136 10616 13142 10628
rect 13817 10625 13829 10628
rect 13863 10625 13875 10659
rect 13817 10619 13875 10625
rect 8205 10591 8263 10597
rect 8205 10588 8217 10591
rect 7300 10560 8217 10588
rect 8205 10557 8217 10560
rect 8251 10557 8263 10591
rect 12161 10591 12219 10597
rect 12161 10588 12173 10591
rect 8205 10551 8263 10557
rect 8404 10560 12173 10588
rect 8404 10532 8432 10560
rect 12161 10557 12173 10560
rect 12207 10588 12219 10591
rect 12250 10588 12256 10600
rect 12207 10560 12256 10588
rect 12207 10557 12219 10560
rect 12161 10551 12219 10557
rect 12250 10548 12256 10560
rect 12308 10548 12314 10600
rect 12802 10588 12808 10600
rect 12763 10560 12808 10588
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 3789 10523 3847 10529
rect 3789 10489 3801 10523
rect 3835 10520 3847 10523
rect 4516 10523 4574 10529
rect 4516 10520 4528 10523
rect 3835 10492 4528 10520
rect 3835 10489 3847 10492
rect 3789 10483 3847 10489
rect 4516 10489 4528 10492
rect 4562 10489 4574 10523
rect 4516 10483 4574 10489
rect 1762 10412 1768 10464
rect 1820 10452 1826 10464
rect 2777 10455 2835 10461
rect 2777 10452 2789 10455
rect 1820 10424 2789 10452
rect 1820 10412 1826 10424
rect 2777 10421 2789 10424
rect 2823 10421 2835 10455
rect 4531 10452 4559 10483
rect 5166 10480 5172 10532
rect 5224 10480 5230 10532
rect 6914 10520 6920 10532
rect 5267 10492 6920 10520
rect 4706 10452 4712 10464
rect 4531 10424 4712 10452
rect 2777 10415 2835 10421
rect 4706 10412 4712 10424
rect 4764 10452 4770 10464
rect 5267 10452 5295 10492
rect 6914 10480 6920 10492
rect 6972 10480 6978 10532
rect 8297 10523 8355 10529
rect 8297 10489 8309 10523
rect 8343 10520 8355 10523
rect 8386 10520 8392 10532
rect 8343 10492 8392 10520
rect 8343 10489 8355 10492
rect 8297 10483 8355 10489
rect 8386 10480 8392 10492
rect 8444 10480 8450 10532
rect 9033 10523 9091 10529
rect 9033 10489 9045 10523
rect 9079 10520 9091 10523
rect 10597 10523 10655 10529
rect 9079 10492 9628 10520
rect 9079 10489 9091 10492
rect 9033 10483 9091 10489
rect 4764 10424 5295 10452
rect 4764 10412 4770 10424
rect 6178 10412 6184 10464
rect 6236 10452 6242 10464
rect 6549 10455 6607 10461
rect 6549 10452 6561 10455
rect 6236 10424 6561 10452
rect 6236 10412 6242 10424
rect 6549 10421 6561 10424
rect 6595 10421 6607 10455
rect 9122 10452 9128 10464
rect 9083 10424 9128 10452
rect 6549 10415 6607 10421
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 9398 10412 9404 10464
rect 9456 10452 9462 10464
rect 9600 10461 9628 10492
rect 10597 10489 10609 10523
rect 10643 10520 10655 10523
rect 10643 10492 11192 10520
rect 10643 10489 10655 10492
rect 10597 10483 10655 10489
rect 11164 10464 11192 10492
rect 9493 10455 9551 10461
rect 9493 10452 9505 10455
rect 9456 10424 9505 10452
rect 9456 10412 9462 10424
rect 9493 10421 9505 10424
rect 9539 10421 9551 10455
rect 9493 10415 9551 10421
rect 9585 10455 9643 10461
rect 9585 10421 9597 10455
rect 9631 10452 9643 10455
rect 9858 10452 9864 10464
rect 9631 10424 9864 10452
rect 9631 10421 9643 10424
rect 9585 10415 9643 10421
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 9950 10412 9956 10464
rect 10008 10452 10014 10464
rect 10137 10455 10195 10461
rect 10137 10452 10149 10455
rect 10008 10424 10149 10452
rect 10008 10412 10014 10424
rect 10137 10421 10149 10424
rect 10183 10421 10195 10455
rect 11054 10452 11060 10464
rect 11015 10424 11060 10452
rect 10137 10415 10195 10421
rect 11054 10412 11060 10424
rect 11112 10412 11118 10464
rect 11146 10412 11152 10464
rect 11204 10452 11210 10464
rect 11204 10424 11249 10452
rect 11204 10412 11210 10424
rect 11606 10412 11612 10464
rect 11664 10452 11670 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 11664 10424 11713 10452
rect 11664 10412 11670 10424
rect 11701 10421 11713 10424
rect 11747 10421 11759 10455
rect 13446 10452 13452 10464
rect 13407 10424 13452 10452
rect 11701 10415 11759 10421
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1762 10248 1768 10260
rect 1723 10220 1768 10248
rect 1762 10208 1768 10220
rect 1820 10208 1826 10260
rect 4062 10248 4068 10260
rect 4023 10220 4068 10248
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 5629 10251 5687 10257
rect 5629 10217 5641 10251
rect 5675 10248 5687 10251
rect 6086 10248 6092 10260
rect 5675 10220 6092 10248
rect 5675 10217 5687 10220
rect 5629 10211 5687 10217
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 7561 10251 7619 10257
rect 7561 10248 7573 10251
rect 7248 10220 7573 10248
rect 7248 10208 7254 10220
rect 7561 10217 7573 10220
rect 7607 10217 7619 10251
rect 7926 10248 7932 10260
rect 7887 10220 7932 10248
rect 7561 10211 7619 10217
rect 7926 10208 7932 10220
rect 7984 10208 7990 10260
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 8665 10251 8723 10257
rect 8665 10248 8677 10251
rect 8168 10220 8677 10248
rect 8168 10208 8174 10220
rect 8665 10217 8677 10220
rect 8711 10217 8723 10251
rect 8665 10211 8723 10217
rect 9953 10251 10011 10257
rect 9953 10217 9965 10251
rect 9999 10248 10011 10251
rect 10042 10248 10048 10260
rect 9999 10220 10048 10248
rect 9999 10217 10011 10220
rect 9953 10211 10011 10217
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10321 10251 10379 10257
rect 10321 10217 10333 10251
rect 10367 10248 10379 10251
rect 10686 10248 10692 10260
rect 10367 10220 10692 10248
rect 10367 10217 10379 10220
rect 10321 10211 10379 10217
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 12342 10248 12348 10260
rect 12303 10220 12348 10248
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 12897 10251 12955 10257
rect 12897 10217 12909 10251
rect 12943 10248 12955 10251
rect 13170 10248 13176 10260
rect 12943 10220 13176 10248
rect 12943 10217 12955 10220
rect 12897 10211 12955 10217
rect 1486 10140 1492 10192
rect 1544 10180 1550 10192
rect 2501 10183 2559 10189
rect 2501 10180 2513 10183
rect 1544 10152 2513 10180
rect 1544 10140 1550 10152
rect 2501 10149 2513 10152
rect 2547 10180 2559 10183
rect 3053 10183 3111 10189
rect 3053 10180 3065 10183
rect 2547 10152 3065 10180
rect 2547 10149 2559 10152
rect 2501 10143 2559 10149
rect 3053 10149 3065 10152
rect 3099 10149 3111 10183
rect 3053 10143 3111 10149
rect 3329 10183 3387 10189
rect 3329 10149 3341 10183
rect 3375 10180 3387 10183
rect 3513 10183 3571 10189
rect 3513 10180 3525 10183
rect 3375 10152 3525 10180
rect 3375 10149 3387 10152
rect 3329 10143 3387 10149
rect 3513 10149 3525 10152
rect 3559 10180 3571 10183
rect 4154 10180 4160 10192
rect 3559 10152 4160 10180
rect 3559 10149 3571 10152
rect 3513 10143 3571 10149
rect 4154 10140 4160 10152
rect 4212 10140 4218 10192
rect 5997 10183 6055 10189
rect 5997 10149 6009 10183
rect 6043 10180 6055 10183
rect 6362 10180 6368 10192
rect 6043 10152 6368 10180
rect 6043 10149 6055 10152
rect 5997 10143 6055 10149
rect 6362 10140 6368 10152
rect 6420 10180 6426 10192
rect 7742 10180 7748 10192
rect 6420 10152 7748 10180
rect 6420 10140 6426 10152
rect 7742 10140 7748 10152
rect 7800 10140 7806 10192
rect 9398 10140 9404 10192
rect 9456 10180 9462 10192
rect 10781 10183 10839 10189
rect 10781 10180 10793 10183
rect 9456 10152 10793 10180
rect 9456 10140 9462 10152
rect 10781 10149 10793 10152
rect 10827 10180 10839 10183
rect 11054 10180 11060 10192
rect 10827 10152 11060 10180
rect 10827 10149 10839 10152
rect 10781 10143 10839 10149
rect 11054 10140 11060 10152
rect 11112 10180 11118 10192
rect 12912 10180 12940 10211
rect 13170 10208 13176 10220
rect 13228 10208 13234 10260
rect 11112 10152 12940 10180
rect 11112 10140 11118 10152
rect 2406 10112 2412 10124
rect 2367 10084 2412 10112
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 4062 10072 4068 10124
rect 4120 10112 4126 10124
rect 4433 10115 4491 10121
rect 4433 10112 4445 10115
rect 4120 10084 4445 10112
rect 4120 10072 4126 10084
rect 4433 10081 4445 10084
rect 4479 10081 4491 10115
rect 4433 10075 4491 10081
rect 7101 10115 7159 10121
rect 7101 10081 7113 10115
rect 7147 10112 7159 10115
rect 7374 10112 7380 10124
rect 7147 10084 7380 10112
rect 7147 10081 7159 10084
rect 7101 10075 7159 10081
rect 7374 10072 7380 10084
rect 7432 10112 7438 10124
rect 7834 10112 7840 10124
rect 7432 10084 7840 10112
rect 7432 10072 7438 10084
rect 7834 10072 7840 10084
rect 7892 10072 7898 10124
rect 8021 10115 8079 10121
rect 8021 10081 8033 10115
rect 8067 10112 8079 10115
rect 9122 10112 9128 10124
rect 8067 10084 9128 10112
rect 8067 10081 8079 10084
rect 8021 10075 8079 10081
rect 9122 10072 9128 10084
rect 9180 10072 9186 10124
rect 11238 10121 11244 10124
rect 11232 10075 11244 10121
rect 11296 10112 11302 10124
rect 11296 10084 11332 10112
rect 11238 10072 11244 10075
rect 11296 10072 11302 10084
rect 2590 10044 2596 10056
rect 2551 10016 2596 10044
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 4709 10047 4767 10053
rect 4709 10013 4721 10047
rect 4755 10044 4767 10047
rect 4798 10044 4804 10056
rect 4755 10016 4804 10044
rect 4755 10013 4767 10016
rect 4709 10007 4767 10013
rect 2958 9936 2964 9988
rect 3016 9976 3022 9988
rect 3789 9979 3847 9985
rect 3789 9976 3801 9979
rect 3016 9948 3801 9976
rect 3016 9936 3022 9948
rect 3789 9945 3801 9948
rect 3835 9976 3847 9979
rect 4540 9976 4568 10007
rect 4798 10004 4804 10016
rect 4856 10004 4862 10056
rect 6086 10044 6092 10056
rect 6047 10016 6092 10044
rect 6086 10004 6092 10016
rect 6144 10004 6150 10056
rect 6178 10004 6184 10056
rect 6236 10044 6242 10056
rect 7190 10044 7196 10056
rect 6236 10016 7052 10044
rect 7151 10016 7196 10044
rect 6236 10004 6242 10016
rect 6730 9976 6736 9988
rect 3835 9948 4568 9976
rect 5000 9948 5939 9976
rect 6691 9948 6736 9976
rect 3835 9945 3847 9948
rect 3789 9939 3847 9945
rect 2038 9908 2044 9920
rect 1999 9880 2044 9908
rect 2038 9868 2044 9880
rect 2096 9868 2102 9920
rect 2498 9868 2504 9920
rect 2556 9908 2562 9920
rect 3329 9911 3387 9917
rect 3329 9908 3341 9911
rect 2556 9880 3341 9908
rect 2556 9868 2562 9880
rect 3329 9877 3341 9880
rect 3375 9877 3387 9911
rect 3329 9871 3387 9877
rect 3418 9868 3424 9920
rect 3476 9908 3482 9920
rect 5000 9908 5028 9948
rect 5166 9908 5172 9920
rect 3476 9880 5028 9908
rect 5127 9880 5172 9908
rect 3476 9868 3482 9880
rect 5166 9868 5172 9880
rect 5224 9908 5230 9920
rect 5445 9911 5503 9917
rect 5445 9908 5457 9911
rect 5224 9880 5457 9908
rect 5224 9868 5230 9880
rect 5445 9877 5457 9880
rect 5491 9877 5503 9911
rect 5911 9908 5939 9948
rect 6730 9936 6736 9948
rect 6788 9936 6794 9988
rect 7024 9976 7052 10016
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 7285 10047 7343 10053
rect 7285 10013 7297 10047
rect 7331 10013 7343 10047
rect 8110 10044 8116 10056
rect 8071 10016 8116 10044
rect 7285 10007 7343 10013
rect 7300 9976 7328 10007
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 10962 10044 10968 10056
rect 10923 10016 10968 10044
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 13170 10044 13176 10056
rect 13131 10016 13176 10044
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 7024 9948 7328 9976
rect 9125 9911 9183 9917
rect 9125 9908 9137 9911
rect 5911 9880 9137 9908
rect 5445 9871 5503 9877
rect 9125 9877 9137 9880
rect 9171 9908 9183 9911
rect 9398 9908 9404 9920
rect 9171 9880 9404 9908
rect 9171 9877 9183 9880
rect 9125 9871 9183 9877
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 13633 9911 13691 9917
rect 13633 9877 13645 9911
rect 13679 9908 13691 9911
rect 13722 9908 13728 9920
rect 13679 9880 13728 9908
rect 13679 9877 13691 9880
rect 13633 9871 13691 9877
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1673 9707 1731 9713
rect 1673 9673 1685 9707
rect 1719 9704 1731 9707
rect 1762 9704 1768 9716
rect 1719 9676 1768 9704
rect 1719 9673 1731 9676
rect 1673 9667 1731 9673
rect 1762 9664 1768 9676
rect 1820 9664 1826 9716
rect 2590 9664 2596 9716
rect 2648 9704 2654 9716
rect 2958 9704 2964 9716
rect 2648 9676 2964 9704
rect 2648 9664 2654 9676
rect 2958 9664 2964 9676
rect 3016 9664 3022 9716
rect 3050 9664 3056 9716
rect 3108 9704 3114 9716
rect 3237 9707 3295 9713
rect 3237 9704 3249 9707
rect 3108 9676 3249 9704
rect 3108 9664 3114 9676
rect 3237 9673 3249 9676
rect 3283 9673 3295 9707
rect 3237 9667 3295 9673
rect 9490 9664 9496 9716
rect 9548 9704 9554 9716
rect 9585 9707 9643 9713
rect 9585 9704 9597 9707
rect 9548 9676 9597 9704
rect 9548 9664 9554 9676
rect 9585 9673 9597 9676
rect 9631 9673 9643 9707
rect 9585 9667 9643 9673
rect 11238 9664 11244 9716
rect 11296 9704 11302 9716
rect 11517 9707 11575 9713
rect 11517 9704 11529 9707
rect 11296 9676 11529 9704
rect 11296 9664 11302 9676
rect 11517 9673 11529 9676
rect 11563 9704 11575 9707
rect 11793 9707 11851 9713
rect 11793 9704 11805 9707
rect 11563 9676 11805 9704
rect 11563 9673 11575 9676
rect 11517 9667 11575 9673
rect 11793 9673 11805 9676
rect 11839 9673 11851 9707
rect 11793 9667 11851 9673
rect 4062 9636 4068 9648
rect 4023 9608 4068 9636
rect 4062 9596 4068 9608
rect 4120 9596 4126 9648
rect 5445 9639 5503 9645
rect 5445 9636 5457 9639
rect 4172 9608 5457 9636
rect 1394 9528 1400 9580
rect 1452 9568 1458 9580
rect 1854 9568 1860 9580
rect 1452 9540 1860 9568
rect 1452 9528 1458 9540
rect 1854 9528 1860 9540
rect 1912 9528 1918 9580
rect 2866 9528 2872 9580
rect 2924 9568 2930 9580
rect 4172 9568 4200 9608
rect 5445 9605 5457 9608
rect 5491 9636 5503 9639
rect 6178 9636 6184 9648
rect 5491 9608 6184 9636
rect 5491 9605 5503 9608
rect 5445 9599 5503 9605
rect 6178 9596 6184 9608
rect 6236 9596 6242 9648
rect 4522 9568 4528 9580
rect 2924 9540 4200 9568
rect 4448 9540 4528 9568
rect 2924 9528 2930 9540
rect 2124 9503 2182 9509
rect 2124 9469 2136 9503
rect 2170 9500 2182 9503
rect 2884 9500 2912 9528
rect 4448 9509 4476 9540
rect 4522 9528 4528 9540
rect 4580 9528 4586 9580
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 5077 9571 5135 9577
rect 5077 9568 5089 9571
rect 4755 9540 5089 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 5077 9537 5089 9540
rect 5123 9568 5135 9571
rect 5258 9568 5264 9580
rect 5123 9540 5264 9568
rect 5123 9537 5135 9540
rect 5077 9531 5135 9537
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 5534 9528 5540 9580
rect 5592 9568 5598 9580
rect 5629 9571 5687 9577
rect 5629 9568 5641 9571
rect 5592 9540 5641 9568
rect 5592 9528 5598 9540
rect 5629 9537 5641 9540
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 2170 9472 2912 9500
rect 3528 9472 4445 9500
rect 2170 9469 2182 9472
rect 2124 9463 2182 9469
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 3528 9373 3556 9472
rect 4433 9469 4445 9472
rect 4479 9469 4491 9503
rect 4433 9463 4491 9469
rect 7190 9460 7196 9512
rect 7248 9500 7254 9512
rect 7561 9503 7619 9509
rect 7561 9500 7573 9503
rect 7248 9472 7573 9500
rect 7248 9460 7254 9472
rect 7561 9469 7573 9472
rect 7607 9469 7619 9503
rect 7561 9463 7619 9469
rect 10137 9503 10195 9509
rect 10137 9469 10149 9503
rect 10183 9500 10195 9503
rect 10686 9500 10692 9512
rect 10183 9472 10692 9500
rect 10183 9469 10195 9472
rect 10137 9463 10195 9469
rect 10686 9460 10692 9472
rect 10744 9500 10750 9512
rect 10962 9500 10968 9512
rect 10744 9472 10968 9500
rect 10744 9460 10750 9472
rect 10962 9460 10968 9472
rect 11020 9460 11026 9512
rect 4525 9435 4583 9441
rect 4525 9432 4537 9435
rect 3896 9404 4537 9432
rect 3513 9367 3571 9373
rect 3513 9364 3525 9367
rect 3476 9336 3525 9364
rect 3476 9324 3482 9336
rect 3513 9333 3525 9336
rect 3559 9333 3571 9367
rect 3513 9327 3571 9333
rect 3786 9324 3792 9376
rect 3844 9364 3850 9376
rect 3896 9373 3924 9404
rect 4525 9401 4537 9404
rect 4571 9432 4583 9435
rect 4890 9432 4896 9444
rect 4571 9404 4896 9432
rect 4571 9401 4583 9404
rect 4525 9395 4583 9401
rect 4890 9392 4896 9404
rect 4948 9392 4954 9444
rect 6362 9392 6368 9444
rect 6420 9392 6426 9444
rect 7466 9392 7472 9444
rect 7524 9432 7530 9444
rect 7806 9435 7864 9441
rect 7806 9432 7818 9435
rect 7524 9404 7818 9432
rect 7524 9392 7530 9404
rect 7806 9401 7818 9404
rect 7852 9432 7864 9435
rect 9217 9435 9275 9441
rect 9217 9432 9229 9435
rect 7852 9404 9229 9432
rect 7852 9401 7864 9404
rect 7806 9395 7864 9401
rect 9217 9401 9229 9404
rect 9263 9432 9275 9435
rect 9766 9432 9772 9444
rect 9263 9404 9772 9432
rect 9263 9401 9275 9404
rect 9217 9395 9275 9401
rect 9766 9392 9772 9404
rect 9824 9392 9830 9444
rect 10382 9435 10440 9441
rect 10382 9432 10394 9435
rect 10060 9404 10394 9432
rect 3881 9367 3939 9373
rect 3881 9364 3893 9367
rect 3844 9336 3893 9364
rect 3844 9324 3850 9336
rect 3881 9333 3893 9336
rect 3927 9333 3939 9367
rect 3881 9327 3939 9333
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 6086 9364 6092 9376
rect 4212 9336 6092 9364
rect 4212 9324 4218 9336
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 6380 9364 6408 9392
rect 10060 9376 10088 9404
rect 10382 9401 10394 9404
rect 10428 9401 10440 9435
rect 11808 9432 11836 9667
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 12492 9608 12537 9636
rect 12492 9596 12498 9608
rect 13722 9596 13728 9648
rect 13780 9636 13786 9648
rect 13780 9608 13825 9636
rect 13780 9596 13786 9608
rect 12342 9528 12348 9580
rect 12400 9568 12406 9580
rect 12802 9568 12808 9580
rect 12400 9540 12808 9568
rect 12400 9528 12406 9540
rect 12802 9528 12808 9540
rect 12860 9568 12866 9580
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12860 9540 13001 9568
rect 12860 9528 12866 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 12158 9500 12164 9512
rect 12119 9472 12164 9500
rect 12158 9460 12164 9472
rect 12216 9500 12222 9512
rect 12897 9503 12955 9509
rect 12897 9500 12909 9503
rect 12216 9472 12909 9500
rect 12216 9460 12222 9472
rect 12897 9469 12909 9472
rect 12943 9469 12955 9503
rect 12897 9463 12955 9469
rect 12986 9432 12992 9444
rect 11808 9404 12992 9432
rect 10382 9395 10440 9401
rect 12986 9392 12992 9404
rect 13044 9392 13050 9444
rect 13725 9435 13783 9441
rect 13725 9432 13737 9435
rect 13188 9404 13737 9432
rect 13188 9376 13216 9404
rect 13725 9401 13737 9404
rect 13771 9432 13783 9435
rect 13817 9435 13875 9441
rect 13817 9432 13829 9435
rect 13771 9404 13829 9432
rect 13771 9401 13783 9404
rect 13725 9395 13783 9401
rect 13817 9401 13829 9404
rect 13863 9401 13875 9435
rect 13817 9395 13875 9401
rect 6457 9367 6515 9373
rect 6457 9364 6469 9367
rect 6236 9336 6469 9364
rect 6236 9324 6242 9336
rect 6457 9333 6469 9336
rect 6503 9333 6515 9367
rect 7098 9364 7104 9376
rect 7059 9336 7104 9364
rect 6457 9327 6515 9333
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 7374 9364 7380 9376
rect 7335 9336 7380 9364
rect 7374 9324 7380 9336
rect 7432 9324 7438 9376
rect 8846 9324 8852 9376
rect 8904 9364 8910 9376
rect 8941 9367 8999 9373
rect 8941 9364 8953 9367
rect 8904 9336 8953 9364
rect 8904 9324 8910 9336
rect 8941 9333 8953 9336
rect 8987 9333 8999 9367
rect 10042 9364 10048 9376
rect 10003 9336 10048 9364
rect 8941 9327 8999 9333
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 12434 9324 12440 9376
rect 12492 9364 12498 9376
rect 12805 9367 12863 9373
rect 12805 9364 12817 9367
rect 12492 9336 12817 9364
rect 12492 9324 12498 9336
rect 12805 9333 12817 9336
rect 12851 9333 12863 9367
rect 12805 9327 12863 9333
rect 13170 9324 13176 9376
rect 13228 9324 13234 9376
rect 13262 9324 13268 9376
rect 13320 9364 13326 9376
rect 13449 9367 13507 9373
rect 13449 9364 13461 9367
rect 13320 9336 13461 9364
rect 13320 9324 13326 9336
rect 13449 9333 13461 9336
rect 13495 9333 13507 9367
rect 13449 9327 13507 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1489 9163 1547 9169
rect 1489 9129 1501 9163
rect 1535 9160 1547 9163
rect 1578 9160 1584 9172
rect 1535 9132 1584 9160
rect 1535 9129 1547 9132
rect 1489 9123 1547 9129
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9160 2007 9163
rect 2038 9160 2044 9172
rect 1995 9132 2044 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 2038 9120 2044 9132
rect 2096 9120 2102 9172
rect 2593 9163 2651 9169
rect 2593 9129 2605 9163
rect 2639 9160 2651 9163
rect 2866 9160 2872 9172
rect 2639 9132 2872 9160
rect 2639 9129 2651 9132
rect 2593 9123 2651 9129
rect 2866 9120 2872 9132
rect 2924 9120 2930 9172
rect 2961 9163 3019 9169
rect 2961 9129 2973 9163
rect 3007 9160 3019 9163
rect 3050 9160 3056 9172
rect 3007 9132 3056 9160
rect 3007 9129 3019 9132
rect 2961 9123 3019 9129
rect 3050 9120 3056 9132
rect 3108 9120 3114 9172
rect 3605 9163 3663 9169
rect 3605 9129 3617 9163
rect 3651 9160 3663 9163
rect 4062 9160 4068 9172
rect 3651 9132 4068 9160
rect 3651 9129 3663 9132
rect 3605 9123 3663 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 6546 9120 6552 9172
rect 6604 9160 6610 9172
rect 6733 9163 6791 9169
rect 6733 9160 6745 9163
rect 6604 9132 6745 9160
rect 6604 9120 6610 9132
rect 6733 9129 6745 9132
rect 6779 9129 6791 9163
rect 6733 9123 6791 9129
rect 7285 9163 7343 9169
rect 7285 9129 7297 9163
rect 7331 9160 7343 9163
rect 8110 9160 8116 9172
rect 7331 9132 8116 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 8110 9120 8116 9132
rect 8168 9120 8174 9172
rect 9122 9120 9128 9172
rect 9180 9160 9186 9172
rect 9401 9163 9459 9169
rect 9401 9160 9413 9163
rect 9180 9132 9413 9160
rect 9180 9120 9186 9132
rect 9401 9129 9413 9132
rect 9447 9129 9459 9163
rect 9401 9123 9459 9129
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10413 9163 10471 9169
rect 10413 9160 10425 9163
rect 10192 9132 10425 9160
rect 10192 9120 10198 9132
rect 10413 9129 10425 9132
rect 10459 9129 10471 9163
rect 12802 9160 12808 9172
rect 12763 9132 12808 9160
rect 10413 9123 10471 9129
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 14001 9163 14059 9169
rect 14001 9160 14013 9163
rect 13780 9132 14013 9160
rect 13780 9120 13786 9132
rect 14001 9129 14013 9132
rect 14047 9129 14059 9163
rect 14001 9123 14059 9129
rect 2056 9092 2084 9120
rect 2682 9092 2688 9104
rect 2056 9064 2688 9092
rect 2682 9052 2688 9064
rect 2740 9052 2746 9104
rect 4338 9092 4344 9104
rect 4299 9064 4344 9092
rect 4338 9052 4344 9064
rect 4396 9052 4402 9104
rect 4890 9052 4896 9104
rect 4948 9092 4954 9104
rect 7374 9092 7380 9104
rect 4948 9064 7380 9092
rect 4948 9052 4954 9064
rect 7374 9052 7380 9064
rect 7432 9052 7438 9104
rect 8389 9095 8447 9101
rect 8389 9061 8401 9095
rect 8435 9092 8447 9095
rect 8478 9092 8484 9104
rect 8435 9064 8484 9092
rect 8435 9061 8447 9064
rect 8389 9055 8447 9061
rect 8478 9052 8484 9064
rect 8536 9052 8542 9104
rect 12434 9092 12440 9104
rect 12395 9064 12440 9092
rect 12434 9052 12440 9064
rect 12492 9052 12498 9104
rect 13357 9095 13415 9101
rect 13357 9061 13369 9095
rect 13403 9092 13415 9095
rect 13446 9092 13452 9104
rect 13403 9064 13452 9092
rect 13403 9061 13415 9064
rect 13357 9055 13415 9061
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 9024 1915 9027
rect 1946 9024 1952 9036
rect 1903 8996 1952 9024
rect 1903 8993 1915 8996
rect 1857 8987 1915 8993
rect 1946 8984 1952 8996
rect 2004 9024 2010 9036
rect 2498 9024 2504 9036
rect 2004 8996 2504 9024
rect 2004 8984 2010 8996
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 3881 9027 3939 9033
rect 3881 8993 3893 9027
rect 3927 8993 3939 9027
rect 3881 8987 3939 8993
rect 1762 8916 1768 8968
rect 1820 8956 1826 8968
rect 2041 8959 2099 8965
rect 2041 8956 2053 8959
rect 1820 8928 2053 8956
rect 1820 8916 1826 8928
rect 2041 8925 2053 8928
rect 2087 8925 2099 8959
rect 3896 8956 3924 8987
rect 3970 8984 3976 9036
rect 4028 9024 4034 9036
rect 4065 9027 4123 9033
rect 4065 9024 4077 9027
rect 4028 8996 4077 9024
rect 4028 8984 4034 8996
rect 4065 8993 4077 8996
rect 4111 8993 4123 9027
rect 4065 8987 4123 8993
rect 4706 8984 4712 9036
rect 4764 9024 4770 9036
rect 5609 9027 5667 9033
rect 5609 9024 5621 9027
rect 4764 8996 5621 9024
rect 4764 8984 4770 8996
rect 5609 8993 5621 8996
rect 5655 9024 5667 9027
rect 6362 9024 6368 9036
rect 5655 8996 6368 9024
rect 5655 8993 5667 8996
rect 5609 8987 5667 8993
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 6730 8984 6736 9036
rect 6788 9024 6794 9036
rect 7929 9027 7987 9033
rect 7929 9024 7941 9027
rect 6788 8996 7941 9024
rect 6788 8984 6794 8996
rect 7929 8993 7941 8996
rect 7975 9024 7987 9027
rect 8018 9024 8024 9036
rect 7975 8996 8024 9024
rect 7975 8993 7987 8996
rect 7929 8987 7987 8993
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 9674 9024 9680 9036
rect 8404 8996 9680 9024
rect 4338 8956 4344 8968
rect 3896 8928 4344 8956
rect 2041 8919 2099 8925
rect 4338 8916 4344 8928
rect 4396 8916 4402 8968
rect 5353 8959 5411 8965
rect 5353 8925 5365 8959
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8956 7711 8959
rect 8404 8956 8432 8996
rect 8588 8965 8616 8996
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 10686 8984 10692 9036
rect 10744 9024 10750 9036
rect 10781 9027 10839 9033
rect 10781 9024 10793 9027
rect 10744 8996 10793 9024
rect 10744 8984 10750 8996
rect 10781 8993 10793 8996
rect 10827 8993 10839 9027
rect 10781 8987 10839 8993
rect 11048 9027 11106 9033
rect 11048 8993 11060 9027
rect 11094 9024 11106 9027
rect 11514 9024 11520 9036
rect 11094 8996 11520 9024
rect 11094 8993 11106 8996
rect 11048 8987 11106 8993
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 7699 8928 8432 8956
rect 8481 8959 8539 8965
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 8481 8925 8493 8959
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8925 8631 8959
rect 9766 8956 9772 8968
rect 9727 8928 9772 8956
rect 8573 8919 8631 8925
rect 5166 8888 5172 8900
rect 3712 8860 5172 8888
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 3712 8829 3740 8860
rect 5166 8848 5172 8860
rect 5224 8888 5230 8900
rect 5368 8888 5396 8919
rect 5224 8860 5396 8888
rect 8496 8888 8524 8919
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 13262 8916 13268 8968
rect 13320 8956 13326 8968
rect 13449 8959 13507 8965
rect 13449 8956 13461 8959
rect 13320 8928 13461 8956
rect 13320 8916 13326 8928
rect 13449 8925 13461 8928
rect 13495 8925 13507 8959
rect 13630 8956 13636 8968
rect 13591 8928 13636 8956
rect 13449 8919 13507 8925
rect 13630 8916 13636 8928
rect 13688 8916 13694 8968
rect 9306 8888 9312 8900
rect 8496 8860 9312 8888
rect 5224 8848 5230 8860
rect 9306 8848 9312 8860
rect 9364 8848 9370 8900
rect 3697 8823 3755 8829
rect 3697 8820 3709 8823
rect 3108 8792 3709 8820
rect 3108 8780 3114 8792
rect 3697 8789 3709 8792
rect 3743 8789 3755 8823
rect 4798 8820 4804 8832
rect 4759 8792 4804 8820
rect 3697 8783 3755 8789
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 5261 8823 5319 8829
rect 5261 8789 5273 8823
rect 5307 8820 5319 8823
rect 5350 8820 5356 8832
rect 5307 8792 5356 8820
rect 5307 8789 5319 8792
rect 5261 8783 5319 8789
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 7742 8820 7748 8832
rect 7703 8792 7748 8820
rect 7742 8780 7748 8792
rect 7800 8780 7806 8832
rect 8018 8820 8024 8832
rect 7979 8792 8024 8820
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 9125 8823 9183 8829
rect 9125 8789 9137 8823
rect 9171 8820 9183 8823
rect 9490 8820 9496 8832
rect 9171 8792 9496 8820
rect 9171 8789 9183 8792
rect 9125 8783 9183 8789
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 12158 8820 12164 8832
rect 12119 8792 12164 8820
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 12989 8823 13047 8829
rect 12989 8789 13001 8823
rect 13035 8820 13047 8823
rect 13722 8820 13728 8832
rect 13035 8792 13728 8820
rect 13035 8789 13047 8792
rect 12989 8783 13047 8789
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 3329 8619 3387 8625
rect 3329 8616 3341 8619
rect 2924 8588 3341 8616
rect 2924 8576 2930 8588
rect 3329 8585 3341 8588
rect 3375 8585 3387 8619
rect 3694 8616 3700 8628
rect 3655 8588 3700 8616
rect 3329 8579 3387 8585
rect 3694 8576 3700 8588
rect 3752 8576 3758 8628
rect 3970 8616 3976 8628
rect 3931 8588 3976 8616
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 4706 8616 4712 8628
rect 4667 8588 4712 8616
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 6454 8576 6460 8628
rect 6512 8616 6518 8628
rect 7098 8616 7104 8628
rect 6512 8588 7104 8616
rect 6512 8576 6518 8588
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 8294 8616 8300 8628
rect 8255 8588 8300 8616
rect 8294 8576 8300 8588
rect 8352 8616 8358 8628
rect 8665 8619 8723 8625
rect 8665 8616 8677 8619
rect 8352 8588 8677 8616
rect 8352 8576 8358 8588
rect 8665 8585 8677 8588
rect 8711 8585 8723 8619
rect 8846 8616 8852 8628
rect 8807 8588 8852 8616
rect 8665 8579 8723 8585
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 9766 8576 9772 8628
rect 9824 8616 9830 8628
rect 11885 8619 11943 8625
rect 11885 8616 11897 8619
rect 9824 8588 11897 8616
rect 9824 8576 9830 8588
rect 11885 8585 11897 8588
rect 11931 8616 11943 8619
rect 11931 8588 12848 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 5166 8548 5172 8560
rect 5127 8520 5172 8548
rect 5166 8508 5172 8520
rect 5224 8508 5230 8560
rect 6825 8551 6883 8557
rect 6825 8548 6837 8551
rect 6104 8520 6837 8548
rect 1854 8440 1860 8492
rect 1912 8480 1918 8492
rect 1949 8483 2007 8489
rect 1949 8480 1961 8483
rect 1912 8452 1961 8480
rect 1912 8440 1918 8452
rect 1949 8449 1961 8452
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 4430 8480 4436 8492
rect 4203 8452 4436 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 1964 8412 1992 8443
rect 4430 8440 4436 8452
rect 4488 8440 4494 8492
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8480 5135 8483
rect 5721 8483 5779 8489
rect 5721 8480 5733 8483
rect 5123 8452 5733 8480
rect 5123 8449 5135 8452
rect 5077 8443 5135 8449
rect 5721 8449 5733 8452
rect 5767 8480 5779 8483
rect 5994 8480 6000 8492
rect 5767 8452 6000 8480
rect 5767 8449 5779 8452
rect 5721 8443 5779 8449
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 3050 8412 3056 8424
rect 1964 8384 3056 8412
rect 3050 8372 3056 8384
rect 3108 8372 3114 8424
rect 5534 8412 5540 8424
rect 5447 8384 5540 8412
rect 5534 8372 5540 8384
rect 5592 8412 5598 8424
rect 6104 8412 6132 8520
rect 6825 8517 6837 8520
rect 6871 8517 6883 8551
rect 6825 8511 6883 8517
rect 8389 8551 8447 8557
rect 8389 8517 8401 8551
rect 8435 8517 8447 8551
rect 8389 8511 8447 8517
rect 10413 8551 10471 8557
rect 10413 8517 10425 8551
rect 10459 8548 10471 8551
rect 12437 8551 12495 8557
rect 10459 8520 11928 8548
rect 10459 8517 10471 8520
rect 10413 8511 10471 8517
rect 6273 8483 6331 8489
rect 6273 8449 6285 8483
rect 6319 8480 6331 8483
rect 6914 8480 6920 8492
rect 6319 8452 6920 8480
rect 6319 8449 6331 8452
rect 6273 8443 6331 8449
rect 6914 8440 6920 8452
rect 6972 8480 6978 8492
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 6972 8452 7389 8480
rect 6972 8440 6978 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 8294 8440 8300 8492
rect 8352 8480 8358 8492
rect 8404 8480 8432 8511
rect 9490 8480 9496 8492
rect 8352 8452 8432 8480
rect 9451 8452 9496 8480
rect 8352 8440 8358 8452
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 9953 8483 10011 8489
rect 9953 8449 9965 8483
rect 9999 8480 10011 8483
rect 10042 8480 10048 8492
rect 9999 8452 10048 8480
rect 9999 8449 10011 8452
rect 9953 8443 10011 8449
rect 10042 8440 10048 8452
rect 10100 8480 10106 8492
rect 10962 8480 10968 8492
rect 10100 8452 10968 8480
rect 10100 8440 10106 8452
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 11900 8480 11928 8520
rect 12437 8517 12449 8551
rect 12483 8548 12495 8551
rect 12618 8548 12624 8560
rect 12483 8520 12624 8548
rect 12483 8517 12495 8520
rect 12437 8511 12495 8517
rect 12618 8508 12624 8520
rect 12676 8508 12682 8560
rect 11900 8452 12756 8480
rect 5592 8384 6132 8412
rect 5592 8372 5598 8384
rect 7742 8372 7748 8424
rect 7800 8412 7806 8424
rect 8573 8415 8631 8421
rect 8573 8412 8585 8415
rect 7800 8384 8585 8412
rect 7800 8372 7806 8384
rect 8573 8381 8585 8384
rect 8619 8412 8631 8415
rect 9674 8412 9680 8424
rect 8619 8384 9680 8412
rect 8619 8381 8631 8384
rect 8573 8375 8631 8381
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 10134 8372 10140 8424
rect 10192 8412 10198 8424
rect 10781 8415 10839 8421
rect 10781 8412 10793 8415
rect 10192 8384 10793 8412
rect 10192 8372 10198 8384
rect 10781 8381 10793 8384
rect 10827 8381 10839 8415
rect 11514 8412 11520 8424
rect 11475 8384 11520 8412
rect 10781 8375 10839 8381
rect 11514 8372 11520 8384
rect 11572 8372 11578 8424
rect 12250 8412 12256 8424
rect 12211 8384 12256 8412
rect 12250 8372 12256 8384
rect 12308 8372 12314 8424
rect 2216 8347 2274 8353
rect 2216 8313 2228 8347
rect 2262 8313 2274 8347
rect 2216 8307 2274 8313
rect 1857 8279 1915 8285
rect 1857 8245 1869 8279
rect 1903 8276 1915 8279
rect 2231 8276 2259 8307
rect 5350 8304 5356 8356
rect 5408 8344 5414 8356
rect 5629 8347 5687 8353
rect 5629 8344 5641 8347
rect 5408 8316 5641 8344
rect 5408 8304 5414 8316
rect 5629 8313 5641 8316
rect 5675 8313 5687 8347
rect 7285 8347 7343 8353
rect 7285 8344 7297 8347
rect 5629 8307 5687 8313
rect 6564 8316 7297 8344
rect 2406 8276 2412 8288
rect 1903 8248 2412 8276
rect 1903 8245 1915 8248
rect 1857 8239 1915 8245
rect 2406 8236 2412 8248
rect 2464 8236 2470 8288
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 6564 8285 6592 8316
rect 7285 8313 7297 8316
rect 7331 8344 7343 8347
rect 7834 8344 7840 8356
rect 7331 8316 7840 8344
rect 7331 8313 7343 8316
rect 7285 8307 7343 8313
rect 7834 8304 7840 8316
rect 7892 8304 7898 8356
rect 7929 8347 7987 8353
rect 7929 8313 7941 8347
rect 7975 8344 7987 8347
rect 8478 8344 8484 8356
rect 7975 8316 8484 8344
rect 7975 8313 7987 8316
rect 7929 8307 7987 8313
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 8665 8347 8723 8353
rect 8665 8313 8677 8347
rect 8711 8344 8723 8347
rect 9217 8347 9275 8353
rect 9217 8344 9229 8347
rect 8711 8316 9229 8344
rect 8711 8313 8723 8316
rect 8665 8307 8723 8313
rect 9217 8313 9229 8316
rect 9263 8313 9275 8347
rect 10229 8347 10287 8353
rect 10229 8344 10241 8347
rect 9217 8307 9275 8313
rect 9324 8316 10241 8344
rect 6549 8279 6607 8285
rect 6549 8276 6561 8279
rect 3016 8248 6561 8276
rect 3016 8236 3022 8248
rect 6549 8245 6561 8248
rect 6595 8245 6607 8279
rect 6549 8239 6607 8245
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 7193 8279 7251 8285
rect 7193 8276 7205 8279
rect 7064 8248 7205 8276
rect 7064 8236 7070 8248
rect 7193 8245 7205 8248
rect 7239 8245 7251 8279
rect 7193 8239 7251 8245
rect 9030 8236 9036 8288
rect 9088 8276 9094 8288
rect 9324 8285 9352 8316
rect 10229 8313 10241 8316
rect 10275 8344 10287 8347
rect 10873 8347 10931 8353
rect 10873 8344 10885 8347
rect 10275 8316 10885 8344
rect 10275 8313 10287 8316
rect 10229 8307 10287 8313
rect 10873 8313 10885 8316
rect 10919 8313 10931 8347
rect 12728 8344 12756 8452
rect 12820 8421 12848 8588
rect 13630 8576 13636 8628
rect 13688 8616 13694 8628
rect 13817 8619 13875 8625
rect 13817 8616 13829 8619
rect 13688 8588 13829 8616
rect 13688 8576 13694 8588
rect 13817 8585 13829 8588
rect 13863 8585 13875 8619
rect 13817 8579 13875 8585
rect 13906 8576 13912 8628
rect 13964 8616 13970 8628
rect 14366 8616 14372 8628
rect 13964 8588 14372 8616
rect 13964 8576 13970 8588
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 17126 8548 17132 8560
rect 17087 8520 17132 8548
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 12986 8480 12992 8492
rect 12947 8452 12992 8480
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 14461 8483 14519 8489
rect 14461 8480 14473 8483
rect 13280 8452 14473 8480
rect 12805 8415 12863 8421
rect 12805 8381 12817 8415
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 12897 8415 12955 8421
rect 12897 8381 12909 8415
rect 12943 8412 12955 8415
rect 13280 8412 13308 8452
rect 14461 8449 14473 8452
rect 14507 8449 14519 8483
rect 14461 8443 14519 8449
rect 13998 8412 14004 8424
rect 12943 8384 13308 8412
rect 13959 8384 14004 8412
rect 12943 8381 12955 8384
rect 12897 8375 12955 8381
rect 12912 8344 12940 8375
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 15746 8412 15752 8424
rect 15707 8384 15752 8412
rect 15746 8372 15752 8384
rect 15804 8372 15810 8424
rect 13538 8344 13544 8356
rect 12728 8316 12940 8344
rect 13188 8316 13544 8344
rect 10873 8307 10931 8313
rect 13188 8288 13216 8316
rect 13538 8304 13544 8316
rect 13596 8304 13602 8356
rect 15994 8347 16052 8353
rect 15994 8344 16006 8347
rect 15672 8316 16006 8344
rect 15672 8288 15700 8316
rect 15994 8313 16006 8316
rect 16040 8313 16052 8347
rect 15994 8307 16052 8313
rect 9309 8279 9367 8285
rect 9309 8276 9321 8279
rect 9088 8248 9321 8276
rect 9088 8236 9094 8248
rect 9309 8245 9321 8248
rect 9355 8245 9367 8279
rect 9309 8239 9367 8245
rect 10686 8236 10692 8288
rect 10744 8276 10750 8288
rect 12069 8279 12127 8285
rect 12069 8276 12081 8279
rect 10744 8248 12081 8276
rect 10744 8236 10750 8248
rect 12069 8245 12081 8248
rect 12115 8276 12127 8279
rect 13170 8276 13176 8288
rect 12115 8248 13176 8276
rect 12115 8245 12127 8248
rect 12069 8239 12127 8245
rect 13170 8236 13176 8248
rect 13228 8236 13234 8288
rect 13446 8276 13452 8288
rect 13407 8248 13452 8276
rect 13446 8236 13452 8248
rect 13504 8236 13510 8288
rect 15654 8276 15660 8288
rect 15615 8248 15660 8276
rect 15654 8236 15660 8248
rect 15712 8236 15718 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 3421 8075 3479 8081
rect 3421 8072 3433 8075
rect 2832 8044 3433 8072
rect 2832 8032 2838 8044
rect 3421 8041 3433 8044
rect 3467 8041 3479 8075
rect 4338 8072 4344 8084
rect 4299 8044 4344 8072
rect 3421 8035 3479 8041
rect 4338 8032 4344 8044
rect 4396 8032 4402 8084
rect 4709 8075 4767 8081
rect 4709 8041 4721 8075
rect 4755 8072 4767 8075
rect 5442 8072 5448 8084
rect 4755 8044 5448 8072
rect 4755 8041 4767 8044
rect 4709 8035 4767 8041
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 6181 8075 6239 8081
rect 6181 8041 6193 8075
rect 6227 8041 6239 8075
rect 6181 8035 6239 8041
rect 6549 8075 6607 8081
rect 6549 8041 6561 8075
rect 6595 8072 6607 8075
rect 6730 8072 6736 8084
rect 6595 8044 6736 8072
rect 6595 8041 6607 8044
rect 6549 8035 6607 8041
rect 1854 8004 1860 8016
rect 1412 7976 1860 8004
rect 1412 7945 1440 7976
rect 1854 7964 1860 7976
rect 1912 7964 1918 8016
rect 2498 7964 2504 8016
rect 2556 8004 2562 8016
rect 5074 8013 5080 8016
rect 3789 8007 3847 8013
rect 3789 8004 3801 8007
rect 2556 7976 3801 8004
rect 2556 7964 2562 7976
rect 3789 7973 3801 7976
rect 3835 7973 3847 8007
rect 5068 8004 5080 8013
rect 5035 7976 5080 8004
rect 3789 7967 3847 7973
rect 5068 7967 5080 7976
rect 5074 7964 5080 7967
rect 5132 7964 5138 8016
rect 5258 7964 5264 8016
rect 5316 8004 5322 8016
rect 6196 8004 6224 8035
rect 6730 8032 6736 8044
rect 6788 8032 6794 8084
rect 7650 8032 7656 8084
rect 7708 8072 7714 8084
rect 9490 8072 9496 8084
rect 7708 8044 9496 8072
rect 7708 8032 7714 8044
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 9861 8075 9919 8081
rect 9861 8072 9873 8075
rect 9732 8044 9873 8072
rect 9732 8032 9738 8044
rect 9861 8041 9873 8044
rect 9907 8041 9919 8075
rect 9861 8035 9919 8041
rect 12897 8075 12955 8081
rect 12897 8041 12909 8075
rect 12943 8072 12955 8075
rect 12986 8072 12992 8084
rect 12943 8044 12992 8072
rect 12943 8041 12955 8044
rect 12897 8035 12955 8041
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 5316 7976 6224 8004
rect 11416 8007 11474 8013
rect 5316 7964 5322 7976
rect 11416 7973 11428 8007
rect 11462 8004 11474 8007
rect 12158 8004 12164 8016
rect 11462 7976 12164 8004
rect 11462 7973 11474 7976
rect 11416 7967 11474 7973
rect 12158 7964 12164 7976
rect 12216 7964 12222 8016
rect 13538 7964 13544 8016
rect 13596 8004 13602 8016
rect 14737 8007 14795 8013
rect 14737 8004 14749 8007
rect 13596 7976 14749 8004
rect 13596 7964 13602 7976
rect 14737 7973 14749 7976
rect 14783 8004 14795 8007
rect 15746 8004 15752 8016
rect 14783 7976 15752 8004
rect 14783 7973 14795 7976
rect 14737 7967 14795 7973
rect 15746 7964 15752 7976
rect 15804 7964 15810 8016
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7905 1455 7939
rect 1397 7899 1455 7905
rect 1664 7939 1722 7945
rect 1664 7905 1676 7939
rect 1710 7936 1722 7939
rect 2222 7936 2228 7948
rect 1710 7908 2228 7936
rect 1710 7905 1722 7908
rect 1664 7899 1722 7905
rect 2222 7896 2228 7908
rect 2280 7896 2286 7948
rect 2774 7896 2780 7948
rect 2832 7936 2838 7948
rect 3145 7939 3203 7945
rect 3145 7936 3157 7939
rect 2832 7908 3157 7936
rect 2832 7896 2838 7908
rect 3145 7905 3157 7908
rect 3191 7936 3203 7939
rect 5276 7936 5304 7964
rect 7466 7945 7472 7948
rect 7460 7936 7472 7945
rect 3191 7908 5304 7936
rect 7427 7908 7472 7936
rect 3191 7905 3203 7908
rect 3145 7899 3203 7905
rect 7460 7899 7472 7908
rect 7466 7896 7472 7899
rect 7524 7896 7530 7948
rect 10686 7896 10692 7948
rect 10744 7936 10750 7948
rect 11149 7939 11207 7945
rect 11149 7936 11161 7939
rect 10744 7908 11161 7936
rect 10744 7896 10750 7908
rect 11149 7905 11161 7908
rect 11195 7905 11207 7939
rect 11149 7899 11207 7905
rect 12986 7896 12992 7948
rect 13044 7936 13050 7948
rect 13725 7939 13783 7945
rect 13725 7936 13737 7939
rect 13044 7908 13737 7936
rect 13044 7896 13050 7908
rect 13725 7905 13737 7908
rect 13771 7905 13783 7939
rect 13725 7899 13783 7905
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 7190 7868 7196 7880
rect 7151 7840 7196 7868
rect 4801 7831 4859 7837
rect 2406 7760 2412 7812
rect 2464 7800 2470 7812
rect 2777 7803 2835 7809
rect 2777 7800 2789 7803
rect 2464 7772 2789 7800
rect 2464 7760 2470 7772
rect 2777 7769 2789 7772
rect 2823 7800 2835 7803
rect 4246 7800 4252 7812
rect 2823 7772 4252 7800
rect 2823 7769 2835 7772
rect 2777 7763 2835 7769
rect 4246 7760 4252 7772
rect 4304 7760 4310 7812
rect 4816 7732 4844 7831
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 10137 7871 10195 7877
rect 10137 7837 10149 7871
rect 10183 7868 10195 7871
rect 10778 7868 10784 7880
rect 10183 7840 10784 7868
rect 10183 7837 10195 7840
rect 10137 7831 10195 7837
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 13170 7828 13176 7880
rect 13228 7868 13234 7880
rect 13817 7871 13875 7877
rect 13817 7868 13829 7871
rect 13228 7840 13829 7868
rect 13228 7828 13234 7840
rect 13817 7837 13829 7840
rect 13863 7837 13875 7871
rect 13817 7831 13875 7837
rect 13909 7871 13967 7877
rect 13909 7837 13921 7871
rect 13955 7837 13967 7871
rect 13909 7831 13967 7837
rect 12526 7800 12532 7812
rect 12487 7772 12532 7800
rect 12526 7760 12532 7772
rect 12584 7760 12590 7812
rect 13924 7800 13952 7831
rect 15838 7828 15844 7880
rect 15896 7868 15902 7880
rect 16025 7871 16083 7877
rect 16025 7868 16037 7871
rect 15896 7840 16037 7868
rect 15896 7828 15902 7840
rect 16025 7837 16037 7840
rect 16071 7837 16083 7871
rect 16025 7831 16083 7837
rect 13188 7772 13952 7800
rect 5442 7732 5448 7744
rect 4816 7704 5448 7732
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 6917 7735 6975 7741
rect 6917 7701 6929 7735
rect 6963 7732 6975 7735
rect 7006 7732 7012 7744
rect 6963 7704 7012 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 8570 7732 8576 7744
rect 8531 7704 8576 7732
rect 8570 7692 8576 7704
rect 8628 7692 8634 7744
rect 8941 7735 8999 7741
rect 8941 7701 8953 7735
rect 8987 7732 8999 7735
rect 9030 7732 9036 7744
rect 8987 7704 9036 7732
rect 8987 7701 8999 7704
rect 8941 7695 8999 7701
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 9306 7732 9312 7744
rect 9267 7704 9312 7732
rect 9306 7692 9312 7704
rect 9364 7692 9370 7744
rect 12894 7692 12900 7744
rect 12952 7732 12958 7744
rect 13188 7741 13216 7772
rect 13173 7735 13231 7741
rect 13173 7732 13185 7735
rect 12952 7704 13185 7732
rect 12952 7692 12958 7704
rect 13173 7701 13185 7704
rect 13219 7701 13231 7735
rect 13173 7695 13231 7701
rect 13357 7735 13415 7741
rect 13357 7701 13369 7735
rect 13403 7732 13415 7735
rect 13814 7732 13820 7744
rect 13403 7704 13820 7732
rect 13403 7701 13415 7704
rect 13357 7695 13415 7701
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 14090 7692 14096 7744
rect 14148 7732 14154 7744
rect 14369 7735 14427 7741
rect 14369 7732 14381 7735
rect 14148 7704 14381 7732
rect 14148 7692 14154 7704
rect 14369 7701 14381 7704
rect 14415 7701 14427 7735
rect 14369 7695 14427 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1397 7531 1455 7537
rect 1397 7497 1409 7531
rect 1443 7528 1455 7531
rect 2590 7528 2596 7540
rect 1443 7500 2596 7528
rect 1443 7497 1455 7500
rect 1397 7491 1455 7497
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 3142 7528 3148 7540
rect 2832 7500 3148 7528
rect 2832 7488 2838 7500
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 4617 7531 4675 7537
rect 4617 7528 4629 7531
rect 4212 7500 4629 7528
rect 4212 7488 4218 7500
rect 4617 7497 4629 7500
rect 4663 7497 4675 7531
rect 4617 7491 4675 7497
rect 6273 7531 6331 7537
rect 6273 7497 6285 7531
rect 6319 7528 6331 7531
rect 7377 7531 7435 7537
rect 7377 7528 7389 7531
rect 6319 7500 7389 7528
rect 6319 7497 6331 7500
rect 6273 7491 6331 7497
rect 7377 7497 7389 7500
rect 7423 7528 7435 7531
rect 7466 7528 7472 7540
rect 7423 7500 7472 7528
rect 7423 7497 7435 7500
rect 7377 7491 7435 7497
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7392 2099 7395
rect 2866 7392 2872 7404
rect 2087 7364 2872 7392
rect 2087 7361 2099 7364
rect 2041 7355 2099 7361
rect 2866 7352 2872 7364
rect 2924 7392 2930 7404
rect 2924 7364 3096 7392
rect 2924 7352 2930 7364
rect 1765 7327 1823 7333
rect 1765 7293 1777 7327
rect 1811 7324 1823 7327
rect 2774 7324 2780 7336
rect 1811 7296 2780 7324
rect 1811 7293 1823 7296
rect 1765 7287 1823 7293
rect 2774 7284 2780 7296
rect 2832 7324 2838 7336
rect 2961 7327 3019 7333
rect 2832 7296 2925 7324
rect 2832 7284 2838 7296
rect 2961 7293 2973 7327
rect 3007 7293 3019 7327
rect 3068 7324 3096 7364
rect 3217 7327 3275 7333
rect 3217 7324 3229 7327
rect 3068 7296 3229 7324
rect 2961 7287 3019 7293
rect 3217 7293 3229 7296
rect 3263 7293 3275 7327
rect 4632 7324 4660 7491
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 6288 7392 6316 7491
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 8754 7528 8760 7540
rect 8036 7500 8760 7528
rect 6822 7392 6828 7404
rect 5859 7364 6316 7392
rect 6783 7364 6828 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 8036 7401 8064 7500
rect 8754 7488 8760 7500
rect 8812 7488 8818 7540
rect 9674 7528 9680 7540
rect 9635 7500 9680 7528
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 12158 7528 12164 7540
rect 11931 7500 12164 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 10137 7395 10195 7401
rect 10137 7361 10149 7395
rect 10183 7392 10195 7395
rect 11425 7395 11483 7401
rect 11425 7392 11437 7395
rect 10183 7364 11437 7392
rect 10183 7361 10195 7364
rect 10137 7355 10195 7361
rect 11425 7361 11437 7364
rect 11471 7392 11483 7395
rect 11900 7392 11928 7491
rect 12158 7488 12164 7500
rect 12216 7488 12222 7540
rect 12986 7528 12992 7540
rect 12947 7500 12992 7528
rect 12986 7488 12992 7500
rect 13044 7488 13050 7540
rect 14458 7488 14464 7540
rect 14516 7528 14522 7540
rect 15105 7531 15163 7537
rect 15105 7528 15117 7531
rect 14516 7500 15117 7528
rect 14516 7488 14522 7500
rect 15105 7497 15117 7500
rect 15151 7497 15163 7531
rect 15838 7528 15844 7540
rect 15799 7500 15844 7528
rect 15105 7491 15163 7497
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 11471 7364 11928 7392
rect 12529 7395 12587 7401
rect 11471 7361 11483 7364
rect 11425 7355 11483 7361
rect 12529 7361 12541 7395
rect 12575 7392 12587 7395
rect 13446 7392 13452 7404
rect 12575 7364 13452 7392
rect 12575 7361 12587 7364
rect 12529 7355 12587 7361
rect 13446 7352 13452 7364
rect 13504 7352 13510 7404
rect 13538 7352 13544 7404
rect 13596 7392 13602 7404
rect 13725 7395 13783 7401
rect 13725 7392 13737 7395
rect 13596 7364 13737 7392
rect 13596 7352 13602 7364
rect 13725 7361 13737 7364
rect 13771 7361 13783 7395
rect 13725 7355 13783 7361
rect 5537 7327 5595 7333
rect 5537 7324 5549 7327
rect 4632 7296 5549 7324
rect 3217 7287 3275 7293
rect 5537 7293 5549 7296
rect 5583 7293 5595 7327
rect 8288 7327 8346 7333
rect 8288 7324 8300 7327
rect 5537 7287 5595 7293
rect 8220 7296 8300 7324
rect 2976 7256 3004 7287
rect 3050 7256 3056 7268
rect 2963 7228 3056 7256
rect 3050 7216 3056 7228
rect 3108 7256 3114 7268
rect 3878 7256 3884 7268
rect 3108 7228 3884 7256
rect 3108 7216 3114 7228
rect 3878 7216 3884 7228
rect 3936 7216 3942 7268
rect 5077 7259 5135 7265
rect 5077 7225 5089 7259
rect 5123 7256 5135 7259
rect 5258 7256 5264 7268
rect 5123 7228 5264 7256
rect 5123 7225 5135 7228
rect 5077 7219 5135 7225
rect 5258 7216 5264 7228
rect 5316 7256 5322 7268
rect 5629 7259 5687 7265
rect 5629 7256 5641 7259
rect 5316 7228 5641 7256
rect 5316 7216 5322 7228
rect 5629 7225 5641 7228
rect 5675 7225 5687 7259
rect 5629 7219 5687 7225
rect 7929 7259 7987 7265
rect 7929 7225 7941 7259
rect 7975 7256 7987 7259
rect 8220 7256 8248 7296
rect 8288 7293 8300 7296
rect 8334 7324 8346 7327
rect 8570 7324 8576 7336
rect 8334 7296 8576 7324
rect 8334 7293 8346 7296
rect 8288 7287 8346 7293
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 9674 7284 9680 7336
rect 9732 7324 9738 7336
rect 10413 7327 10471 7333
rect 10413 7324 10425 7327
rect 9732 7296 10425 7324
rect 9732 7284 9738 7296
rect 10413 7293 10425 7296
rect 10459 7293 10471 7327
rect 10413 7287 10471 7293
rect 10778 7284 10784 7336
rect 10836 7324 10842 7336
rect 11149 7327 11207 7333
rect 11149 7324 11161 7327
rect 10836 7296 11161 7324
rect 10836 7284 10842 7296
rect 11149 7293 11161 7296
rect 11195 7293 11207 7327
rect 11149 7287 11207 7293
rect 11238 7284 11244 7336
rect 11296 7324 11302 7336
rect 12161 7327 12219 7333
rect 12161 7324 12173 7327
rect 11296 7296 12173 7324
rect 11296 7284 11302 7296
rect 12161 7293 12173 7296
rect 12207 7293 12219 7327
rect 15856 7324 15884 7488
rect 16482 7392 16488 7404
rect 16443 7364 16488 7392
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 16301 7327 16359 7333
rect 16301 7324 16313 7327
rect 15856 7296 16313 7324
rect 12161 7287 12219 7293
rect 16301 7293 16313 7296
rect 16347 7293 16359 7327
rect 16301 7287 16359 7293
rect 7975 7228 8248 7256
rect 13992 7259 14050 7265
rect 7975 7225 7987 7228
rect 7929 7219 7987 7225
rect 13992 7225 14004 7259
rect 14038 7256 14050 7259
rect 14090 7256 14096 7268
rect 14038 7228 14096 7256
rect 14038 7225 14050 7228
rect 13992 7219 14050 7225
rect 14090 7216 14096 7228
rect 14148 7216 14154 7268
rect 15473 7259 15531 7265
rect 15473 7225 15485 7259
rect 15519 7256 15531 7259
rect 15654 7256 15660 7268
rect 15519 7228 15660 7256
rect 15519 7225 15531 7228
rect 15473 7219 15531 7225
rect 15654 7216 15660 7228
rect 15712 7256 15718 7268
rect 16482 7256 16488 7268
rect 15712 7228 16488 7256
rect 15712 7216 15718 7228
rect 16482 7216 16488 7228
rect 16540 7216 16546 7268
rect 1857 7191 1915 7197
rect 1857 7157 1869 7191
rect 1903 7188 1915 7191
rect 2498 7188 2504 7200
rect 1903 7160 2504 7188
rect 1903 7157 1915 7160
rect 1857 7151 1915 7157
rect 2498 7148 2504 7160
rect 2556 7148 2562 7200
rect 3510 7148 3516 7200
rect 3568 7188 3574 7200
rect 4341 7191 4399 7197
rect 4341 7188 4353 7191
rect 3568 7160 4353 7188
rect 3568 7148 3574 7160
rect 4341 7157 4353 7160
rect 4387 7188 4399 7191
rect 4798 7188 4804 7200
rect 4387 7160 4804 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 5166 7188 5172 7200
rect 5127 7160 5172 7188
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 5442 7148 5448 7200
rect 5500 7188 5506 7200
rect 6641 7191 6699 7197
rect 6641 7188 6653 7191
rect 5500 7160 6653 7188
rect 5500 7148 5506 7160
rect 6641 7157 6653 7160
rect 6687 7188 6699 7191
rect 7190 7188 7196 7200
rect 6687 7160 7196 7188
rect 6687 7157 6699 7160
rect 6641 7151 6699 7157
rect 7190 7148 7196 7160
rect 7248 7188 7254 7200
rect 8202 7188 8208 7200
rect 7248 7160 8208 7188
rect 7248 7148 7254 7160
rect 8202 7148 8208 7160
rect 8260 7148 8266 7200
rect 9398 7188 9404 7200
rect 9359 7160 9404 7188
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 10229 7191 10287 7197
rect 10229 7188 10241 7191
rect 10192 7160 10241 7188
rect 10192 7148 10198 7160
rect 10229 7157 10241 7160
rect 10275 7157 10287 7191
rect 10778 7188 10784 7200
rect 10739 7160 10784 7188
rect 10229 7151 10287 7157
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 13357 7191 13415 7197
rect 13357 7188 13369 7191
rect 13228 7160 13369 7188
rect 13228 7148 13234 7160
rect 13357 7157 13369 7160
rect 13403 7157 13415 7191
rect 15930 7188 15936 7200
rect 15891 7160 15936 7188
rect 13357 7151 13415 7157
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 16390 7188 16396 7200
rect 16351 7160 16396 7188
rect 16390 7148 16396 7160
rect 16448 7188 16454 7200
rect 16945 7191 17003 7197
rect 16945 7188 16957 7191
rect 16448 7160 16957 7188
rect 16448 7148 16454 7160
rect 16945 7157 16957 7160
rect 16991 7157 17003 7191
rect 16945 7151 17003 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2866 6984 2872 6996
rect 2827 6956 2872 6984
rect 2866 6944 2872 6956
rect 2924 6944 2930 6996
rect 4065 6987 4123 6993
rect 4065 6984 4077 6987
rect 3232 6956 4077 6984
rect 2314 6876 2320 6928
rect 2372 6916 2378 6928
rect 3232 6916 3260 6956
rect 4065 6953 4077 6956
rect 4111 6953 4123 6987
rect 4065 6947 4123 6953
rect 4893 6987 4951 6993
rect 4893 6953 4905 6987
rect 4939 6984 4951 6987
rect 5074 6984 5080 6996
rect 4939 6956 5080 6984
rect 4939 6953 4951 6956
rect 4893 6947 4951 6953
rect 5074 6944 5080 6956
rect 5132 6944 5138 6996
rect 9030 6944 9036 6996
rect 9088 6984 9094 6996
rect 9674 6984 9680 6996
rect 9088 6956 9680 6984
rect 9088 6944 9094 6956
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 12897 6987 12955 6993
rect 12897 6953 12909 6987
rect 12943 6984 12955 6987
rect 13538 6984 13544 6996
rect 12943 6956 13544 6984
rect 12943 6953 12955 6956
rect 12897 6947 12955 6953
rect 3878 6916 3884 6928
rect 2372 6888 3260 6916
rect 3791 6888 3884 6916
rect 2372 6876 2378 6888
rect 3878 6876 3884 6888
rect 3936 6916 3942 6928
rect 3936 6888 5488 6916
rect 3936 6876 3942 6888
rect 5460 6860 5488 6888
rect 10134 6876 10140 6928
rect 10192 6916 10198 6928
rect 12912 6916 12940 6947
rect 13538 6944 13544 6956
rect 13596 6984 13602 6996
rect 14645 6987 14703 6993
rect 14645 6984 14657 6987
rect 13596 6956 14657 6984
rect 13596 6944 13602 6956
rect 14645 6953 14657 6956
rect 14691 6984 14703 6987
rect 15654 6984 15660 6996
rect 14691 6956 15660 6984
rect 14691 6953 14703 6956
rect 14645 6947 14703 6953
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 16390 6916 16396 6928
rect 10192 6888 11008 6916
rect 10192 6876 10198 6888
rect 1762 6848 1768 6860
rect 1723 6820 1768 6848
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 2222 6808 2228 6860
rect 2280 6848 2286 6860
rect 2280 6820 2636 6848
rect 2280 6808 2286 6820
rect 1578 6740 1584 6792
rect 1636 6780 1642 6792
rect 1857 6783 1915 6789
rect 1857 6780 1869 6783
rect 1636 6752 1869 6780
rect 1636 6740 1642 6752
rect 1857 6749 1869 6752
rect 1903 6749 1915 6783
rect 1857 6743 1915 6749
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6780 2099 6783
rect 2608 6780 2636 6820
rect 4338 6808 4344 6860
rect 4396 6848 4402 6860
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 4396 6820 5365 6848
rect 4396 6808 4402 6820
rect 5353 6817 5365 6820
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 5442 6808 5448 6860
rect 5500 6848 5506 6860
rect 5712 6851 5770 6857
rect 5500 6820 5545 6848
rect 5500 6808 5506 6820
rect 5712 6817 5724 6851
rect 5758 6848 5770 6851
rect 6730 6848 6736 6860
rect 5758 6820 6736 6848
rect 5758 6817 5770 6820
rect 5712 6811 5770 6817
rect 6730 6808 6736 6820
rect 6788 6808 6794 6860
rect 7098 6848 7104 6860
rect 7059 6820 7104 6848
rect 7098 6808 7104 6820
rect 7156 6808 7162 6860
rect 8110 6848 8116 6860
rect 8071 6820 8116 6848
rect 8110 6808 8116 6820
rect 8168 6808 8174 6860
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 10318 6857 10324 6860
rect 8260 6820 8305 6848
rect 8260 6808 8266 6820
rect 10312 6811 10324 6857
rect 10376 6848 10382 6860
rect 10980 6848 11008 6888
rect 12820 6888 12940 6916
rect 15120 6888 16396 6916
rect 12161 6851 12219 6857
rect 12161 6848 12173 6851
rect 10376 6820 10412 6848
rect 10980 6820 12173 6848
rect 10318 6808 10324 6811
rect 10376 6808 10382 6820
rect 12161 6817 12173 6820
rect 12207 6848 12219 6851
rect 12250 6848 12256 6860
rect 12207 6820 12256 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 12250 6808 12256 6820
rect 12308 6808 12314 6860
rect 12820 6792 12848 6888
rect 12894 6808 12900 6860
rect 12952 6848 12958 6860
rect 13245 6851 13303 6857
rect 13245 6848 13257 6851
rect 12952 6820 13257 6848
rect 12952 6808 12958 6820
rect 13245 6817 13257 6820
rect 13291 6817 13303 6851
rect 13245 6811 13303 6817
rect 14826 6808 14832 6860
rect 14884 6848 14890 6860
rect 15120 6848 15148 6888
rect 16390 6876 16396 6888
rect 16448 6876 16454 6928
rect 15746 6848 15752 6860
rect 14884 6820 15148 6848
rect 15580 6820 15752 6848
rect 14884 6808 14890 6820
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2087 6752 2452 6780
rect 2608 6752 2973 6780
rect 2087 6749 2099 6752
rect 2041 6743 2099 6749
rect 2424 6656 2452 6752
rect 2961 6749 2973 6752
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6780 8447 6783
rect 8570 6780 8576 6792
rect 8435 6752 8576 6780
rect 8435 6749 8447 6752
rect 8389 6743 8447 6749
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 10045 6783 10103 6789
rect 10045 6749 10057 6783
rect 10091 6749 10103 6783
rect 12802 6780 12808 6792
rect 12715 6752 12808 6780
rect 10045 6743 10103 6749
rect 7742 6712 7748 6724
rect 7703 6684 7748 6712
rect 7742 6672 7748 6684
rect 7800 6672 7806 6724
rect 8294 6672 8300 6724
rect 8352 6712 8358 6724
rect 8352 6684 9168 6712
rect 8352 6672 8358 6684
rect 9140 6656 9168 6684
rect 1394 6644 1400 6656
rect 1355 6616 1400 6644
rect 1394 6604 1400 6616
rect 1452 6604 1458 6656
rect 2406 6644 2412 6656
rect 2367 6616 2412 6644
rect 2406 6604 2412 6616
rect 2464 6604 2470 6656
rect 3510 6644 3516 6656
rect 3471 6616 3516 6644
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 5169 6647 5227 6653
rect 5169 6613 5181 6647
rect 5215 6644 5227 6647
rect 5442 6644 5448 6656
rect 5215 6616 5448 6644
rect 5215 6613 5227 6616
rect 5169 6607 5227 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 6086 6604 6092 6656
rect 6144 6644 6150 6656
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 6144 6616 6837 6644
rect 6144 6604 6150 6616
rect 6825 6613 6837 6616
rect 6871 6613 6883 6647
rect 7466 6644 7472 6656
rect 7427 6616 7472 6644
rect 6825 6607 6883 6613
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 8754 6644 8760 6656
rect 8715 6616 8760 6644
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 9122 6644 9128 6656
rect 9083 6616 9128 6644
rect 9122 6604 9128 6616
rect 9180 6644 9186 6656
rect 9861 6647 9919 6653
rect 9861 6644 9873 6647
rect 9180 6616 9873 6644
rect 9180 6604 9186 6616
rect 9861 6613 9873 6616
rect 9907 6613 9919 6647
rect 10060 6644 10088 6743
rect 12802 6740 12808 6752
rect 12860 6780 12866 6792
rect 12989 6783 13047 6789
rect 12989 6780 13001 6783
rect 12860 6752 13001 6780
rect 12860 6740 12866 6752
rect 12989 6749 13001 6752
rect 13035 6749 13047 6783
rect 12989 6743 13047 6749
rect 15105 6783 15163 6789
rect 15105 6749 15117 6783
rect 15151 6780 15163 6783
rect 15580 6780 15608 6820
rect 15746 6808 15752 6820
rect 15804 6848 15810 6860
rect 15913 6851 15971 6857
rect 15913 6848 15925 6851
rect 15804 6820 15925 6848
rect 15804 6808 15810 6820
rect 15913 6817 15925 6820
rect 15959 6817 15971 6851
rect 17862 6848 17868 6860
rect 17823 6820 17868 6848
rect 15913 6811 15971 6817
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 15151 6752 15608 6780
rect 15151 6749 15163 6752
rect 15105 6743 15163 6749
rect 15654 6740 15660 6792
rect 15712 6789 15718 6792
rect 15712 6780 15722 6789
rect 18138 6780 18144 6792
rect 15712 6752 15757 6780
rect 18099 6752 18144 6780
rect 15712 6743 15722 6752
rect 15712 6740 15718 6743
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 10778 6644 10784 6656
rect 10060 6616 10784 6644
rect 9861 6607 9919 6613
rect 10778 6604 10784 6616
rect 10836 6604 10842 6656
rect 11422 6644 11428 6656
rect 11383 6616 11428 6644
rect 11422 6604 11428 6616
rect 11480 6604 11486 6656
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 11701 6647 11759 6653
rect 11701 6644 11713 6647
rect 11664 6616 11713 6644
rect 11664 6604 11670 6616
rect 11701 6613 11713 6616
rect 11747 6644 11759 6647
rect 12437 6647 12495 6653
rect 12437 6644 12449 6647
rect 11747 6616 12449 6644
rect 11747 6613 11759 6616
rect 11701 6607 11759 6613
rect 12437 6613 12449 6616
rect 12483 6613 12495 6647
rect 12437 6607 12495 6613
rect 14090 6604 14096 6656
rect 14148 6644 14154 6656
rect 14369 6647 14427 6653
rect 14369 6644 14381 6647
rect 14148 6616 14381 6644
rect 14148 6604 14154 6616
rect 14369 6613 14381 6616
rect 14415 6613 14427 6647
rect 14369 6607 14427 6613
rect 16574 6604 16580 6656
rect 16632 6644 16638 6656
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 16632 6616 17049 6644
rect 16632 6604 16638 6616
rect 17037 6613 17049 6616
rect 17083 6613 17095 6647
rect 17037 6607 17095 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1762 6400 1768 6452
rect 1820 6440 1826 6452
rect 1949 6443 2007 6449
rect 1949 6440 1961 6443
rect 1820 6412 1961 6440
rect 1820 6400 1826 6412
rect 1949 6409 1961 6412
rect 1995 6409 2007 6443
rect 1949 6403 2007 6409
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 4985 6443 5043 6449
rect 4985 6440 4997 6443
rect 4212 6412 4997 6440
rect 4212 6400 4218 6412
rect 4985 6409 4997 6412
rect 5031 6440 5043 6443
rect 6822 6440 6828 6452
rect 5031 6412 5304 6440
rect 6783 6412 6828 6440
rect 5031 6409 5043 6412
rect 4985 6403 5043 6409
rect 4065 6375 4123 6381
rect 4065 6341 4077 6375
rect 4111 6372 4123 6375
rect 4338 6372 4344 6384
rect 4111 6344 4344 6372
rect 4111 6341 4123 6344
rect 4065 6335 4123 6341
rect 4338 6332 4344 6344
rect 4396 6332 4402 6384
rect 5169 6375 5227 6381
rect 5169 6341 5181 6375
rect 5215 6341 5227 6375
rect 5169 6335 5227 6341
rect 2038 6264 2044 6316
rect 2096 6304 2102 6316
rect 2406 6304 2412 6316
rect 2096 6276 2412 6304
rect 2096 6264 2102 6276
rect 2406 6264 2412 6276
rect 2464 6304 2470 6316
rect 2777 6307 2835 6313
rect 2777 6304 2789 6307
rect 2464 6276 2789 6304
rect 2464 6264 2470 6276
rect 2777 6273 2789 6276
rect 2823 6273 2835 6307
rect 2777 6267 2835 6273
rect 2682 6196 2688 6248
rect 2740 6196 2746 6248
rect 5184 6236 5212 6335
rect 5276 6304 5304 6412
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 7929 6443 7987 6449
rect 7929 6409 7941 6443
rect 7975 6440 7987 6443
rect 8110 6440 8116 6452
rect 7975 6412 8116 6440
rect 7975 6409 7987 6412
rect 7929 6403 7987 6409
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 8297 6443 8355 6449
rect 8297 6409 8309 6443
rect 8343 6440 8355 6443
rect 8570 6440 8576 6452
rect 8343 6412 8576 6440
rect 8343 6409 8355 6412
rect 8297 6403 8355 6409
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 9766 6400 9772 6452
rect 9824 6440 9830 6452
rect 10137 6443 10195 6449
rect 10137 6440 10149 6443
rect 9824 6412 10149 6440
rect 9824 6400 9830 6412
rect 10137 6409 10149 6412
rect 10183 6409 10195 6443
rect 10137 6403 10195 6409
rect 10318 6400 10324 6452
rect 10376 6440 10382 6452
rect 10413 6443 10471 6449
rect 10413 6440 10425 6443
rect 10376 6412 10425 6440
rect 10376 6400 10382 6412
rect 10413 6409 10425 6412
rect 10459 6409 10471 6443
rect 10413 6403 10471 6409
rect 11422 6400 11428 6452
rect 11480 6440 11486 6452
rect 11701 6443 11759 6449
rect 11701 6440 11713 6443
rect 11480 6412 11713 6440
rect 11480 6400 11486 6412
rect 11701 6409 11713 6412
rect 11747 6440 11759 6443
rect 11882 6440 11888 6452
rect 11747 6412 11888 6440
rect 11747 6409 11759 6412
rect 11701 6403 11759 6409
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 13078 6400 13084 6452
rect 13136 6440 13142 6452
rect 13446 6440 13452 6452
rect 13136 6412 13452 6440
rect 13136 6400 13142 6412
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 14826 6400 14832 6452
rect 14884 6440 14890 6452
rect 15013 6443 15071 6449
rect 15013 6440 15025 6443
rect 14884 6412 15025 6440
rect 14884 6400 14890 6412
rect 15013 6409 15025 6412
rect 15059 6409 15071 6443
rect 15013 6403 15071 6409
rect 15654 6400 15660 6452
rect 15712 6440 15718 6452
rect 16393 6443 16451 6449
rect 16393 6440 16405 6443
rect 15712 6412 16405 6440
rect 15712 6400 15718 6412
rect 16393 6409 16405 6412
rect 16439 6409 16451 6443
rect 16393 6403 16451 6409
rect 17862 6400 17868 6452
rect 17920 6440 17926 6452
rect 18509 6443 18567 6449
rect 18509 6440 18521 6443
rect 17920 6412 18521 6440
rect 17920 6400 17926 6412
rect 18509 6409 18521 6412
rect 18555 6409 18567 6443
rect 18509 6403 18567 6409
rect 5534 6332 5540 6384
rect 5592 6372 5598 6384
rect 6273 6375 6331 6381
rect 6273 6372 6285 6375
rect 5592 6344 6285 6372
rect 5592 6332 5598 6344
rect 6273 6341 6285 6344
rect 6319 6372 6331 6375
rect 6730 6372 6736 6384
rect 6319 6344 6736 6372
rect 6319 6341 6331 6344
rect 6273 6335 6331 6341
rect 6730 6332 6736 6344
rect 6788 6332 6794 6384
rect 5629 6307 5687 6313
rect 5629 6304 5641 6307
rect 5276 6276 5641 6304
rect 5629 6273 5641 6276
rect 5675 6273 5687 6307
rect 5629 6267 5687 6273
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 5994 6304 6000 6316
rect 5859 6276 6000 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 5994 6264 6000 6276
rect 6052 6264 6058 6316
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6304 6699 6307
rect 7374 6304 7380 6316
rect 6687 6276 7380 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6304 8723 6307
rect 12802 6304 12808 6316
rect 8711 6276 8892 6304
rect 12763 6276 12808 6304
rect 8711 6273 8723 6276
rect 8665 6267 8723 6273
rect 7193 6239 7251 6245
rect 7193 6236 7205 6239
rect 5184 6208 7205 6236
rect 7193 6205 7205 6208
rect 7239 6236 7251 6239
rect 7466 6236 7472 6248
rect 7239 6208 7472 6236
rect 7239 6205 7251 6208
rect 7193 6199 7251 6205
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 8757 6239 8815 6245
rect 8757 6205 8769 6239
rect 8803 6205 8815 6239
rect 8864 6236 8892 6276
rect 12802 6264 12808 6276
rect 12860 6264 12866 6316
rect 15657 6307 15715 6313
rect 15657 6273 15669 6307
rect 15703 6304 15715 6307
rect 15746 6304 15752 6316
rect 15703 6276 15752 6304
rect 15703 6273 15715 6276
rect 15657 6267 15715 6273
rect 15746 6264 15752 6276
rect 15804 6304 15810 6316
rect 16114 6304 16120 6316
rect 15804 6276 16120 6304
rect 15804 6264 15810 6276
rect 16114 6264 16120 6276
rect 16172 6264 16178 6316
rect 9024 6239 9082 6245
rect 9024 6236 9036 6239
rect 8864 6208 9036 6236
rect 8757 6199 8815 6205
rect 9024 6205 9036 6208
rect 9070 6236 9082 6239
rect 9398 6236 9404 6248
rect 9070 6208 9404 6236
rect 9070 6205 9082 6208
rect 9024 6199 9082 6205
rect 1670 6128 1676 6180
rect 1728 6168 1734 6180
rect 2593 6171 2651 6177
rect 1728 6140 2544 6168
rect 1728 6128 1734 6140
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 2225 6103 2283 6109
rect 2225 6069 2237 6103
rect 2271 6100 2283 6103
rect 2406 6100 2412 6112
rect 2271 6072 2412 6100
rect 2271 6069 2283 6072
rect 2225 6063 2283 6069
rect 2406 6060 2412 6072
rect 2464 6060 2470 6112
rect 2516 6100 2544 6140
rect 2593 6137 2605 6171
rect 2639 6168 2651 6171
rect 2700 6168 2728 6196
rect 3605 6171 3663 6177
rect 3605 6168 3617 6171
rect 2639 6140 3617 6168
rect 2639 6137 2651 6140
rect 2593 6131 2651 6137
rect 3605 6137 3617 6140
rect 3651 6137 3663 6171
rect 3605 6131 3663 6137
rect 4157 6171 4215 6177
rect 4157 6137 4169 6171
rect 4203 6168 4215 6171
rect 4709 6171 4767 6177
rect 4709 6168 4721 6171
rect 4203 6140 4721 6168
rect 4203 6137 4215 6140
rect 4157 6131 4215 6137
rect 4709 6137 4721 6140
rect 4755 6168 4767 6171
rect 5537 6171 5595 6177
rect 5537 6168 5549 6171
rect 4755 6140 5549 6168
rect 4755 6137 4767 6140
rect 4709 6131 4767 6137
rect 5537 6137 5549 6140
rect 5583 6137 5595 6171
rect 5537 6131 5595 6137
rect 7098 6128 7104 6180
rect 7156 6168 7162 6180
rect 7285 6171 7343 6177
rect 7285 6168 7297 6171
rect 7156 6140 7297 6168
rect 7156 6128 7162 6140
rect 7285 6137 7297 6140
rect 7331 6137 7343 6171
rect 7285 6131 7343 6137
rect 2685 6103 2743 6109
rect 2685 6100 2697 6103
rect 2516 6072 2697 6100
rect 2685 6069 2697 6072
rect 2731 6100 2743 6103
rect 3237 6103 3295 6109
rect 3237 6100 3249 6103
rect 2731 6072 3249 6100
rect 2731 6069 2743 6072
rect 2685 6063 2743 6069
rect 3237 6069 3249 6072
rect 3283 6069 3295 6103
rect 8772 6100 8800 6199
rect 9398 6196 9404 6208
rect 9456 6196 9462 6248
rect 13078 6245 13084 6248
rect 13072 6236 13084 6245
rect 12991 6208 13084 6236
rect 13072 6199 13084 6208
rect 13136 6236 13142 6248
rect 13630 6236 13636 6248
rect 13136 6208 13636 6236
rect 13078 6196 13084 6199
rect 13136 6196 13142 6208
rect 13630 6196 13636 6208
rect 13688 6196 13694 6248
rect 14550 6196 14556 6248
rect 14608 6236 14614 6248
rect 15381 6239 15439 6245
rect 15381 6236 15393 6239
rect 14608 6208 15393 6236
rect 14608 6196 14614 6208
rect 15381 6205 15393 6208
rect 15427 6205 15439 6239
rect 16574 6236 16580 6248
rect 16535 6208 16580 6236
rect 15381 6199 15439 6205
rect 16574 6196 16580 6208
rect 16632 6236 16638 6248
rect 17313 6239 17371 6245
rect 17313 6236 17325 6239
rect 16632 6208 17325 6236
rect 16632 6196 16638 6208
rect 17313 6205 17325 6208
rect 17359 6205 17371 6239
rect 19518 6236 19524 6248
rect 19479 6208 19524 6236
rect 17313 6199 17371 6205
rect 19518 6196 19524 6208
rect 19576 6236 19582 6248
rect 20257 6239 20315 6245
rect 20257 6236 20269 6239
rect 19576 6208 20269 6236
rect 19576 6196 19582 6208
rect 20257 6205 20269 6208
rect 20303 6205 20315 6239
rect 20257 6199 20315 6205
rect 12713 6171 12771 6177
rect 12713 6137 12725 6171
rect 12759 6168 12771 6171
rect 13087 6168 13115 6196
rect 15473 6171 15531 6177
rect 15473 6168 15485 6171
rect 12759 6140 13115 6168
rect 14844 6140 15485 6168
rect 12759 6137 12771 6140
rect 12713 6131 12771 6137
rect 10778 6100 10784 6112
rect 8772 6072 10784 6100
rect 3237 6063 3295 6069
rect 10778 6060 10784 6072
rect 10836 6060 10842 6112
rect 11146 6100 11152 6112
rect 11107 6072 11152 6100
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 12253 6103 12311 6109
rect 12253 6069 12265 6103
rect 12299 6100 12311 6103
rect 12894 6100 12900 6112
rect 12299 6072 12900 6100
rect 12299 6069 12311 6072
rect 12253 6063 12311 6069
rect 12894 6060 12900 6072
rect 12952 6100 12958 6112
rect 14185 6103 14243 6109
rect 14185 6100 14197 6103
rect 12952 6072 14197 6100
rect 12952 6060 12958 6072
rect 14185 6069 14197 6072
rect 14231 6069 14243 6103
rect 14185 6063 14243 6069
rect 14734 6060 14740 6112
rect 14792 6100 14798 6112
rect 14844 6109 14872 6140
rect 15473 6137 15485 6140
rect 15519 6137 15531 6171
rect 16850 6168 16856 6180
rect 16811 6140 16856 6168
rect 15473 6131 15531 6137
rect 16850 6128 16856 6140
rect 16908 6128 16914 6180
rect 19797 6171 19855 6177
rect 19797 6137 19809 6171
rect 19843 6168 19855 6171
rect 20530 6168 20536 6180
rect 19843 6140 20536 6168
rect 19843 6137 19855 6140
rect 19797 6131 19855 6137
rect 20530 6128 20536 6140
rect 20588 6128 20594 6180
rect 14829 6103 14887 6109
rect 14829 6100 14841 6103
rect 14792 6072 14841 6100
rect 14792 6060 14798 6072
rect 14829 6069 14841 6072
rect 14875 6069 14887 6103
rect 16114 6100 16120 6112
rect 16075 6072 16120 6100
rect 14829 6063 14887 6069
rect 16114 6060 16120 6072
rect 16172 6060 16178 6112
rect 18046 6100 18052 6112
rect 18007 6072 18052 6100
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1397 5899 1455 5905
rect 1397 5865 1409 5899
rect 1443 5896 1455 5899
rect 1762 5896 1768 5908
rect 1443 5868 1768 5896
rect 1443 5865 1455 5868
rect 1397 5859 1455 5865
rect 1762 5856 1768 5868
rect 1820 5856 1826 5908
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5896 2467 5899
rect 2682 5896 2688 5908
rect 2455 5868 2688 5896
rect 2455 5865 2467 5868
rect 2409 5859 2467 5865
rect 2682 5856 2688 5868
rect 2740 5856 2746 5908
rect 2777 5899 2835 5905
rect 2777 5865 2789 5899
rect 2823 5896 2835 5899
rect 3694 5896 3700 5908
rect 2823 5868 3700 5896
rect 2823 5865 2835 5868
rect 2777 5859 2835 5865
rect 3694 5856 3700 5868
rect 3752 5856 3758 5908
rect 4614 5896 4620 5908
rect 4575 5868 4620 5896
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5353 5899 5411 5905
rect 5353 5865 5365 5899
rect 5399 5896 5411 5899
rect 5534 5896 5540 5908
rect 5399 5868 5540 5896
rect 5399 5865 5411 5868
rect 5353 5859 5411 5865
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 5721 5899 5779 5905
rect 5721 5865 5733 5899
rect 5767 5896 5779 5899
rect 5994 5896 6000 5908
rect 5767 5868 6000 5896
rect 5767 5865 5779 5868
rect 5721 5859 5779 5865
rect 5994 5856 6000 5868
rect 6052 5856 6058 5908
rect 7374 5896 7380 5908
rect 7335 5868 7380 5896
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 8110 5856 8116 5908
rect 8168 5896 8174 5908
rect 8205 5899 8263 5905
rect 8205 5896 8217 5899
rect 8168 5868 8217 5896
rect 8168 5856 8174 5868
rect 8205 5865 8217 5868
rect 8251 5865 8263 5899
rect 8754 5896 8760 5908
rect 8715 5868 8760 5896
rect 8205 5859 8263 5865
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 9122 5896 9128 5908
rect 9083 5868 9128 5896
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 10042 5856 10048 5908
rect 10100 5896 10106 5908
rect 11054 5896 11060 5908
rect 10100 5868 11060 5896
rect 10100 5856 10106 5868
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 12618 5896 12624 5908
rect 12492 5868 12624 5896
rect 12492 5856 12498 5868
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 13078 5896 13084 5908
rect 13039 5868 13084 5896
rect 13078 5856 13084 5868
rect 13136 5856 13142 5908
rect 13538 5856 13544 5908
rect 13596 5896 13602 5908
rect 13725 5899 13783 5905
rect 13725 5896 13737 5899
rect 13596 5868 13737 5896
rect 13596 5856 13602 5868
rect 13725 5865 13737 5868
rect 13771 5865 13783 5899
rect 13725 5859 13783 5865
rect 16114 5856 16120 5908
rect 16172 5896 16178 5908
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 16172 5868 17693 5896
rect 16172 5856 16178 5868
rect 17681 5865 17693 5868
rect 17727 5865 17739 5899
rect 17681 5859 17739 5865
rect 6012 5828 6040 5856
rect 6242 5831 6300 5837
rect 6242 5828 6254 5831
rect 6012 5800 6254 5828
rect 6242 5797 6254 5800
rect 6288 5797 6300 5831
rect 6242 5791 6300 5797
rect 11882 5788 11888 5840
rect 11940 5837 11946 5840
rect 11940 5831 12004 5837
rect 11940 5797 11958 5831
rect 11992 5828 12004 5831
rect 11992 5800 12388 5828
rect 11992 5797 12004 5800
rect 11940 5791 12004 5797
rect 11940 5788 11946 5791
rect 12360 5772 12388 5800
rect 14550 5788 14556 5840
rect 14608 5828 14614 5840
rect 15013 5831 15071 5837
rect 15013 5828 15025 5831
rect 14608 5800 15025 5828
rect 14608 5788 14614 5800
rect 15013 5797 15025 5800
rect 15059 5797 15071 5831
rect 15013 5791 15071 5797
rect 3234 5720 3240 5772
rect 3292 5760 3298 5772
rect 3513 5763 3571 5769
rect 3513 5760 3525 5763
rect 3292 5732 3525 5760
rect 3292 5720 3298 5732
rect 3513 5729 3525 5732
rect 3559 5760 3571 5763
rect 3881 5763 3939 5769
rect 3881 5760 3893 5763
rect 3559 5732 3893 5760
rect 3559 5729 3571 5732
rect 3513 5723 3571 5729
rect 3881 5729 3893 5732
rect 3927 5760 3939 5763
rect 5442 5760 5448 5772
rect 3927 5732 5448 5760
rect 3927 5729 3939 5732
rect 3881 5723 3939 5729
rect 5442 5720 5448 5732
rect 5500 5760 5506 5772
rect 5997 5763 6055 5769
rect 5997 5760 6009 5763
rect 5500 5732 6009 5760
rect 5500 5720 5506 5732
rect 5997 5729 6009 5732
rect 6043 5760 6055 5763
rect 6546 5760 6552 5772
rect 6043 5732 6552 5760
rect 6043 5729 6055 5732
rect 5997 5723 6055 5729
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 7837 5763 7895 5769
rect 7837 5729 7849 5763
rect 7883 5760 7895 5763
rect 8202 5760 8208 5772
rect 7883 5732 8208 5760
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 9398 5720 9404 5772
rect 9456 5760 9462 5772
rect 10045 5763 10103 5769
rect 10045 5760 10057 5763
rect 9456 5732 10057 5760
rect 9456 5720 9462 5732
rect 10045 5729 10057 5732
rect 10091 5729 10103 5763
rect 10045 5723 10103 5729
rect 11149 5763 11207 5769
rect 11149 5729 11161 5763
rect 11195 5760 11207 5763
rect 11425 5763 11483 5769
rect 11425 5760 11437 5763
rect 11195 5732 11437 5760
rect 11195 5729 11207 5732
rect 11149 5723 11207 5729
rect 11425 5729 11437 5732
rect 11471 5760 11483 5763
rect 12250 5760 12256 5772
rect 11471 5732 12256 5760
rect 11471 5729 11483 5732
rect 11425 5723 11483 5729
rect 12250 5720 12256 5732
rect 12308 5720 12314 5772
rect 12342 5720 12348 5772
rect 12400 5720 12406 5772
rect 13909 5763 13967 5769
rect 13909 5729 13921 5763
rect 13955 5760 13967 5763
rect 14182 5760 14188 5772
rect 13955 5732 14188 5760
rect 13955 5729 13967 5732
rect 13909 5723 13967 5729
rect 14182 5720 14188 5732
rect 14240 5720 14246 5772
rect 16574 5769 16580 5772
rect 16568 5760 16580 5769
rect 16535 5732 16580 5760
rect 16568 5723 16580 5732
rect 16574 5720 16580 5723
rect 16632 5720 16638 5772
rect 18138 5720 18144 5772
rect 18196 5760 18202 5772
rect 18509 5763 18567 5769
rect 18509 5760 18521 5763
rect 18196 5732 18521 5760
rect 18196 5720 18202 5732
rect 18509 5729 18521 5732
rect 18555 5729 18567 5763
rect 18509 5723 18567 5729
rect 19613 5763 19671 5769
rect 19613 5729 19625 5763
rect 19659 5760 19671 5763
rect 20622 5760 20628 5772
rect 19659 5732 20628 5760
rect 19659 5729 19671 5732
rect 19613 5723 19671 5729
rect 20622 5720 20628 5732
rect 20680 5720 20686 5772
rect 2866 5692 2872 5704
rect 2148 5664 2872 5692
rect 2148 5568 2176 5664
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5661 3019 5695
rect 2961 5655 3019 5661
rect 2314 5624 2320 5636
rect 2227 5596 2320 5624
rect 2314 5584 2320 5596
rect 2372 5624 2378 5636
rect 2976 5624 3004 5655
rect 4430 5652 4436 5704
rect 4488 5692 4494 5704
rect 4709 5695 4767 5701
rect 4709 5692 4721 5695
rect 4488 5664 4721 5692
rect 4488 5652 4494 5664
rect 4709 5661 4721 5664
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 4798 5652 4804 5704
rect 4856 5692 4862 5704
rect 10137 5695 10195 5701
rect 4856 5664 4901 5692
rect 4856 5652 4862 5664
rect 10137 5661 10149 5695
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 2372 5596 3004 5624
rect 2372 5584 2378 5596
rect 8294 5584 8300 5636
rect 8352 5624 8358 5636
rect 9401 5627 9459 5633
rect 9401 5624 9413 5627
rect 8352 5596 9413 5624
rect 8352 5584 8358 5596
rect 9401 5593 9413 5596
rect 9447 5624 9459 5627
rect 10152 5624 10180 5655
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 10284 5664 10329 5692
rect 10284 5652 10290 5664
rect 11606 5652 11612 5704
rect 11664 5692 11670 5704
rect 11701 5695 11759 5701
rect 11701 5692 11713 5695
rect 11664 5664 11713 5692
rect 11664 5652 11670 5664
rect 11701 5661 11713 5664
rect 11747 5661 11759 5695
rect 11701 5655 11759 5661
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5692 14151 5695
rect 14734 5692 14740 5704
rect 14139 5664 14740 5692
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 10962 5624 10968 5636
rect 9447 5596 10180 5624
rect 10612 5596 10968 5624
rect 9447 5593 9459 5596
rect 9401 5587 9459 5593
rect 1949 5559 2007 5565
rect 1949 5525 1961 5559
rect 1995 5556 2007 5559
rect 2038 5556 2044 5568
rect 1995 5528 2044 5556
rect 1995 5525 2007 5528
rect 1949 5519 2007 5525
rect 2038 5516 2044 5528
rect 2096 5516 2102 5568
rect 2130 5516 2136 5568
rect 2188 5516 2194 5568
rect 4154 5516 4160 5568
rect 4212 5556 4218 5568
rect 4249 5559 4307 5565
rect 4249 5556 4261 5559
rect 4212 5528 4261 5556
rect 4212 5516 4218 5528
rect 4249 5525 4261 5528
rect 4295 5525 4307 5559
rect 4249 5519 4307 5525
rect 9677 5559 9735 5565
rect 9677 5525 9689 5559
rect 9723 5556 9735 5559
rect 10612 5556 10640 5596
rect 10962 5584 10968 5596
rect 11020 5584 11026 5636
rect 10778 5556 10784 5568
rect 9723 5528 10640 5556
rect 10739 5528 10784 5556
rect 9723 5525 9735 5528
rect 9677 5519 9735 5525
rect 10778 5516 10784 5528
rect 10836 5556 10842 5568
rect 11241 5559 11299 5565
rect 11241 5556 11253 5559
rect 10836 5528 11253 5556
rect 10836 5516 10842 5528
rect 11241 5525 11253 5528
rect 11287 5556 11299 5559
rect 11716 5556 11744 5655
rect 14734 5652 14740 5664
rect 14792 5652 14798 5704
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5692 15347 5695
rect 16206 5692 16212 5704
rect 15335 5664 16212 5692
rect 15335 5661 15347 5664
rect 15289 5655 15347 5661
rect 16206 5652 16212 5664
rect 16264 5652 16270 5704
rect 16301 5695 16359 5701
rect 16301 5661 16313 5695
rect 16347 5661 16359 5695
rect 16301 5655 16359 5661
rect 16316 5624 16344 5655
rect 15764 5596 16344 5624
rect 13357 5559 13415 5565
rect 13357 5556 13369 5559
rect 11287 5528 13369 5556
rect 11287 5525 11299 5528
rect 11241 5519 11299 5525
rect 13357 5525 13369 5528
rect 13403 5525 13415 5559
rect 13357 5519 13415 5525
rect 15470 5516 15476 5568
rect 15528 5556 15534 5568
rect 15764 5565 15792 5596
rect 15749 5559 15807 5565
rect 15749 5556 15761 5559
rect 15528 5528 15761 5556
rect 15528 5516 15534 5528
rect 15749 5525 15761 5528
rect 15795 5525 15807 5559
rect 15749 5519 15807 5525
rect 16209 5559 16267 5565
rect 16209 5525 16221 5559
rect 16255 5556 16267 5559
rect 16482 5556 16488 5568
rect 16255 5528 16488 5556
rect 16255 5525 16267 5528
rect 16209 5519 16267 5525
rect 16482 5516 16488 5528
rect 16540 5516 16546 5568
rect 18693 5559 18751 5565
rect 18693 5525 18705 5559
rect 18739 5556 18751 5559
rect 18782 5556 18788 5568
rect 18739 5528 18788 5556
rect 18739 5525 18751 5528
rect 18693 5519 18751 5525
rect 18782 5516 18788 5528
rect 18840 5516 18846 5568
rect 19797 5559 19855 5565
rect 19797 5525 19809 5559
rect 19843 5556 19855 5559
rect 20990 5556 20996 5568
rect 19843 5528 20996 5556
rect 19843 5525 19855 5528
rect 19797 5519 19855 5525
rect 20990 5516 20996 5528
rect 21048 5516 21054 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 4614 5352 4620 5364
rect 4575 5324 4620 5352
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 5169 5355 5227 5361
rect 5169 5321 5181 5355
rect 5215 5352 5227 5355
rect 5350 5352 5356 5364
rect 5215 5324 5356 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 6546 5312 6552 5364
rect 6604 5352 6610 5364
rect 7929 5355 7987 5361
rect 7929 5352 7941 5355
rect 6604 5324 7941 5352
rect 6604 5312 6610 5324
rect 7929 5321 7941 5324
rect 7975 5352 7987 5355
rect 8297 5355 8355 5361
rect 8297 5352 8309 5355
rect 7975 5324 8309 5352
rect 7975 5321 7987 5324
rect 7929 5315 7987 5321
rect 8297 5321 8309 5324
rect 8343 5352 8355 5355
rect 8754 5352 8760 5364
rect 8343 5324 8760 5352
rect 8343 5321 8355 5324
rect 8297 5315 8355 5321
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 11330 5312 11336 5364
rect 11388 5352 11394 5364
rect 12250 5352 12256 5364
rect 11388 5324 12256 5352
rect 11388 5312 11394 5324
rect 12250 5312 12256 5324
rect 12308 5312 12314 5364
rect 12437 5355 12495 5361
rect 12437 5321 12449 5355
rect 12483 5352 12495 5355
rect 13262 5352 13268 5364
rect 12483 5324 13268 5352
rect 12483 5321 12495 5324
rect 12437 5315 12495 5321
rect 13262 5312 13268 5324
rect 13320 5312 13326 5364
rect 13909 5355 13967 5361
rect 13909 5321 13921 5355
rect 13955 5352 13967 5355
rect 13998 5352 14004 5364
rect 13955 5324 14004 5352
rect 13955 5321 13967 5324
rect 13909 5315 13967 5321
rect 13998 5312 14004 5324
rect 14056 5312 14062 5364
rect 14182 5312 14188 5364
rect 14240 5352 14246 5364
rect 15013 5355 15071 5361
rect 15013 5352 15025 5355
rect 14240 5324 15025 5352
rect 14240 5312 14246 5324
rect 15013 5321 15025 5324
rect 15059 5321 15071 5355
rect 15013 5315 15071 5321
rect 18138 5312 18144 5364
rect 18196 5352 18202 5364
rect 18785 5355 18843 5361
rect 18785 5352 18797 5355
rect 18196 5324 18797 5352
rect 18196 5312 18202 5324
rect 18785 5321 18797 5324
rect 18831 5321 18843 5355
rect 18785 5315 18843 5321
rect 11790 5284 11796 5296
rect 11751 5256 11796 5284
rect 11790 5244 11796 5256
rect 11848 5244 11854 5296
rect 5534 5176 5540 5228
rect 5592 5216 5598 5228
rect 5721 5219 5779 5225
rect 5721 5216 5733 5219
rect 5592 5188 5733 5216
rect 5592 5176 5598 5188
rect 5721 5185 5733 5188
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 7098 5176 7104 5228
rect 7156 5216 7162 5228
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 7156 5188 7389 5216
rect 7156 5176 7162 5188
rect 7377 5185 7389 5188
rect 7423 5185 7435 5219
rect 7377 5179 7435 5185
rect 8478 5176 8484 5228
rect 8536 5216 8542 5228
rect 8573 5219 8631 5225
rect 8573 5216 8585 5219
rect 8536 5188 8585 5216
rect 8536 5176 8542 5188
rect 8573 5185 8585 5188
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 1762 5108 1768 5160
rect 1820 5148 1826 5160
rect 1949 5151 2007 5157
rect 1949 5148 1961 5151
rect 1820 5120 1961 5148
rect 1820 5108 1826 5120
rect 1949 5117 1961 5120
rect 1995 5148 2007 5151
rect 3234 5148 3240 5160
rect 1995 5120 3240 5148
rect 1995 5117 2007 5120
rect 1949 5111 2007 5117
rect 3234 5108 3240 5120
rect 3292 5108 3298 5160
rect 3694 5148 3700 5160
rect 3655 5120 3700 5148
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 4982 5108 4988 5160
rect 5040 5148 5046 5160
rect 5077 5151 5135 5157
rect 5077 5148 5089 5151
rect 5040 5120 5089 5148
rect 5040 5108 5046 5120
rect 5077 5117 5089 5120
rect 5123 5148 5135 5151
rect 5629 5151 5687 5157
rect 5629 5148 5641 5151
rect 5123 5120 5641 5148
rect 5123 5117 5135 5120
rect 5077 5111 5135 5117
rect 5629 5117 5641 5120
rect 5675 5148 5687 5151
rect 6086 5148 6092 5160
rect 5675 5120 6092 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 6086 5108 6092 5120
rect 6144 5108 6150 5160
rect 7193 5151 7251 5157
rect 7193 5148 7205 5151
rect 6196 5120 7205 5148
rect 2038 5040 2044 5092
rect 2096 5080 2102 5092
rect 2216 5083 2274 5089
rect 2216 5080 2228 5083
rect 2096 5052 2228 5080
rect 2096 5040 2102 5052
rect 2216 5049 2228 5052
rect 2262 5080 2274 5083
rect 3142 5080 3148 5092
rect 2262 5052 3148 5080
rect 2262 5049 2274 5052
rect 2216 5043 2274 5049
rect 3142 5040 3148 5052
rect 3200 5040 3206 5092
rect 1857 5015 1915 5021
rect 1857 4981 1869 5015
rect 1903 5012 1915 5015
rect 2130 5012 2136 5024
rect 1903 4984 2136 5012
rect 1903 4981 1915 4984
rect 1857 4975 1915 4981
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 3326 5012 3332 5024
rect 3287 4984 3332 5012
rect 3326 4972 3332 4984
rect 3384 4972 3390 5024
rect 4341 5015 4399 5021
rect 4341 4981 4353 5015
rect 4387 5012 4399 5015
rect 4430 5012 4436 5024
rect 4387 4984 4436 5012
rect 4387 4981 4399 4984
rect 4341 4975 4399 4981
rect 4430 4972 4436 4984
rect 4488 4972 4494 5024
rect 5166 4972 5172 5024
rect 5224 5012 5230 5024
rect 5537 5015 5595 5021
rect 5537 5012 5549 5015
rect 5224 4984 5549 5012
rect 5224 4972 5230 4984
rect 5537 4981 5549 4984
rect 5583 4981 5595 5015
rect 5537 4975 5595 4981
rect 6086 4972 6092 5024
rect 6144 5012 6150 5024
rect 6196 5021 6224 5120
rect 7193 5117 7205 5120
rect 7239 5148 7251 5151
rect 7926 5148 7932 5160
rect 7239 5120 7932 5148
rect 7239 5117 7251 5120
rect 7193 5111 7251 5117
rect 7926 5108 7932 5120
rect 7984 5108 7990 5160
rect 9585 5151 9643 5157
rect 9585 5117 9597 5151
rect 9631 5148 9643 5151
rect 10778 5148 10784 5160
rect 9631 5120 10784 5148
rect 9631 5117 9643 5120
rect 9585 5111 9643 5117
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 11808 5148 11836 5244
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 12989 5219 13047 5225
rect 12989 5216 13001 5219
rect 12492 5188 13001 5216
rect 12492 5176 12498 5188
rect 12989 5185 13001 5188
rect 13035 5216 13047 5219
rect 13449 5219 13507 5225
rect 13449 5216 13461 5219
rect 13035 5188 13461 5216
rect 13035 5185 13047 5188
rect 12989 5179 13047 5185
rect 13449 5185 13461 5188
rect 13495 5185 13507 5219
rect 13449 5179 13507 5185
rect 14090 5176 14096 5228
rect 14148 5216 14154 5228
rect 14553 5219 14611 5225
rect 14553 5216 14565 5219
rect 14148 5188 14565 5216
rect 14148 5176 14154 5188
rect 14553 5185 14565 5188
rect 14599 5185 14611 5219
rect 14553 5179 14611 5185
rect 16025 5219 16083 5225
rect 16025 5185 16037 5219
rect 16071 5216 16083 5219
rect 16574 5216 16580 5228
rect 16071 5188 16580 5216
rect 16071 5185 16083 5188
rect 16025 5179 16083 5185
rect 16574 5176 16580 5188
rect 16632 5216 16638 5228
rect 16761 5219 16819 5225
rect 16761 5216 16773 5219
rect 16632 5188 16773 5216
rect 16632 5176 16638 5188
rect 16761 5185 16773 5188
rect 16807 5216 16819 5219
rect 16807 5188 17264 5216
rect 16807 5185 16819 5188
rect 16761 5179 16819 5185
rect 12805 5151 12863 5157
rect 12805 5148 12817 5151
rect 11808 5120 12817 5148
rect 12805 5117 12817 5120
rect 12851 5117 12863 5151
rect 12805 5111 12863 5117
rect 13998 5108 14004 5160
rect 14056 5148 14062 5160
rect 14369 5151 14427 5157
rect 14369 5148 14381 5151
rect 14056 5120 14381 5148
rect 14056 5108 14062 5120
rect 14369 5117 14381 5120
rect 14415 5117 14427 5151
rect 14369 5111 14427 5117
rect 6546 5040 6552 5092
rect 6604 5080 6610 5092
rect 6641 5083 6699 5089
rect 6641 5080 6653 5083
rect 6604 5052 6653 5080
rect 6604 5040 6610 5052
rect 6641 5049 6653 5052
rect 6687 5080 6699 5083
rect 7285 5083 7343 5089
rect 7285 5080 7297 5083
rect 6687 5052 7297 5080
rect 6687 5049 6699 5052
rect 6641 5043 6699 5049
rect 7285 5049 7297 5052
rect 7331 5080 7343 5083
rect 8110 5080 8116 5092
rect 7331 5052 8116 5080
rect 7331 5049 7343 5052
rect 7285 5043 7343 5049
rect 8110 5040 8116 5052
rect 8168 5040 8174 5092
rect 9125 5083 9183 5089
rect 9125 5049 9137 5083
rect 9171 5080 9183 5083
rect 9171 5052 9536 5080
rect 9171 5049 9183 5052
rect 9125 5043 9183 5049
rect 6181 5015 6239 5021
rect 6181 5012 6193 5015
rect 6144 4984 6193 5012
rect 6144 4972 6150 4984
rect 6181 4981 6193 4984
rect 6227 4981 6239 5015
rect 6822 5012 6828 5024
rect 6783 4984 6828 5012
rect 6181 4975 6239 4981
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 8294 4972 8300 5024
rect 8352 5012 8358 5024
rect 9398 5012 9404 5024
rect 8352 4984 9404 5012
rect 8352 4972 8358 4984
rect 9398 4972 9404 4984
rect 9456 4972 9462 5024
rect 9508 5012 9536 5052
rect 9766 5040 9772 5092
rect 9824 5089 9830 5092
rect 9824 5083 9888 5089
rect 9824 5049 9842 5083
rect 9876 5080 9888 5083
rect 11241 5083 11299 5089
rect 11241 5080 11253 5083
rect 9876 5052 11253 5080
rect 9876 5049 9888 5052
rect 9824 5043 9888 5049
rect 11241 5049 11253 5052
rect 11287 5049 11299 5083
rect 11241 5043 11299 5049
rect 9824 5040 9830 5043
rect 13814 5040 13820 5092
rect 13872 5080 13878 5092
rect 14458 5080 14464 5092
rect 13872 5052 14464 5080
rect 13872 5040 13878 5052
rect 14458 5040 14464 5052
rect 14516 5040 14522 5092
rect 15657 5083 15715 5089
rect 15657 5049 15669 5083
rect 15703 5080 15715 5083
rect 16022 5080 16028 5092
rect 15703 5052 16028 5080
rect 15703 5049 15715 5052
rect 15657 5043 15715 5049
rect 16022 5040 16028 5052
rect 16080 5080 16086 5092
rect 16485 5083 16543 5089
rect 16485 5080 16497 5083
rect 16080 5052 16497 5080
rect 16080 5040 16086 5052
rect 16485 5049 16497 5052
rect 16531 5049 16543 5083
rect 16485 5043 16543 5049
rect 10134 5012 10140 5024
rect 9508 4984 10140 5012
rect 10134 4972 10140 4984
rect 10192 4972 10198 5024
rect 10686 4972 10692 5024
rect 10744 5012 10750 5024
rect 10965 5015 11023 5021
rect 10965 5012 10977 5015
rect 10744 4984 10977 5012
rect 10744 4972 10750 4984
rect 10965 4981 10977 4984
rect 11011 4981 11023 5015
rect 10965 4975 11023 4981
rect 12253 5015 12311 5021
rect 12253 4981 12265 5015
rect 12299 5012 12311 5015
rect 12894 5012 12900 5024
rect 12299 4984 12900 5012
rect 12299 4981 12311 4984
rect 12253 4975 12311 4981
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 14001 5015 14059 5021
rect 14001 4981 14013 5015
rect 14047 5012 14059 5015
rect 14826 5012 14832 5024
rect 14047 4984 14832 5012
rect 14047 4981 14059 4984
rect 14001 4975 14059 4981
rect 14826 4972 14832 4984
rect 14884 4972 14890 5024
rect 16114 5012 16120 5024
rect 16075 4984 16120 5012
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 16574 5012 16580 5024
rect 16535 4984 16580 5012
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 17236 5021 17264 5188
rect 17865 5151 17923 5157
rect 17865 5117 17877 5151
rect 17911 5148 17923 5151
rect 18046 5148 18052 5160
rect 17911 5120 18052 5148
rect 17911 5117 17923 5120
rect 17865 5111 17923 5117
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 19337 5151 19395 5157
rect 19337 5117 19349 5151
rect 19383 5148 19395 5151
rect 19426 5148 19432 5160
rect 19383 5120 19432 5148
rect 19383 5117 19395 5120
rect 19337 5111 19395 5117
rect 19426 5108 19432 5120
rect 19484 5148 19490 5160
rect 19889 5151 19947 5157
rect 19889 5148 19901 5151
rect 19484 5120 19901 5148
rect 19484 5108 19490 5120
rect 19889 5117 19901 5120
rect 19935 5117 19947 5151
rect 20530 5148 20536 5160
rect 20491 5120 20536 5148
rect 19889 5111 19947 5117
rect 20530 5108 20536 5120
rect 20588 5148 20594 5160
rect 21085 5151 21143 5157
rect 21085 5148 21097 5151
rect 20588 5120 21097 5148
rect 20588 5108 20594 5120
rect 21085 5117 21097 5120
rect 21131 5117 21143 5151
rect 21085 5111 21143 5117
rect 18322 5080 18328 5092
rect 18283 5052 18328 5080
rect 18322 5040 18328 5052
rect 18380 5040 18386 5092
rect 17221 5015 17279 5021
rect 17221 4981 17233 5015
rect 17267 5012 17279 5015
rect 17402 5012 17408 5024
rect 17267 4984 17408 5012
rect 17267 4981 17279 4984
rect 17221 4975 17279 4981
rect 17402 4972 17408 4984
rect 17460 4972 17466 5024
rect 19334 4972 19340 5024
rect 19392 5012 19398 5024
rect 19521 5015 19579 5021
rect 19521 5012 19533 5015
rect 19392 4984 19533 5012
rect 19392 4972 19398 4984
rect 19521 4981 19533 4984
rect 19567 4981 19579 5015
rect 19521 4975 19579 4981
rect 20349 5015 20407 5021
rect 20349 4981 20361 5015
rect 20395 5012 20407 5015
rect 20622 5012 20628 5024
rect 20395 4984 20628 5012
rect 20395 4981 20407 4984
rect 20349 4975 20407 4981
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 20717 5015 20775 5021
rect 20717 4981 20729 5015
rect 20763 5012 20775 5015
rect 22554 5012 22560 5024
rect 20763 4984 22560 5012
rect 20763 4981 20775 4984
rect 20717 4975 20775 4981
rect 22554 4972 22560 4984
rect 22612 4972 22618 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 3142 4808 3148 4820
rect 3103 4780 3148 4808
rect 3142 4768 3148 4780
rect 3200 4808 3206 4820
rect 3421 4811 3479 4817
rect 3421 4808 3433 4811
rect 3200 4780 3433 4808
rect 3200 4768 3206 4780
rect 3421 4777 3433 4780
rect 3467 4777 3479 4811
rect 3421 4771 3479 4777
rect 3881 4811 3939 4817
rect 3881 4777 3893 4811
rect 3927 4808 3939 4811
rect 4062 4808 4068 4820
rect 3927 4780 4068 4808
rect 3927 4777 3939 4780
rect 3881 4771 3939 4777
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 6730 4768 6736 4820
rect 6788 4808 6794 4820
rect 6917 4811 6975 4817
rect 6917 4808 6929 4811
rect 6788 4780 6929 4808
rect 6788 4768 6794 4780
rect 6917 4777 6929 4780
rect 6963 4777 6975 4811
rect 6917 4771 6975 4777
rect 8021 4811 8079 4817
rect 8021 4777 8033 4811
rect 8067 4808 8079 4811
rect 8202 4808 8208 4820
rect 8067 4780 8208 4808
rect 8067 4777 8079 4780
rect 8021 4771 8079 4777
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 8754 4768 8760 4820
rect 8812 4808 8818 4820
rect 9033 4811 9091 4817
rect 9033 4808 9045 4811
rect 8812 4780 9045 4808
rect 8812 4768 8818 4780
rect 9033 4777 9045 4780
rect 9079 4777 9091 4811
rect 9033 4771 9091 4777
rect 11054 4768 11060 4820
rect 11112 4808 11118 4820
rect 11609 4811 11667 4817
rect 11609 4808 11621 4811
rect 11112 4780 11621 4808
rect 11112 4768 11118 4780
rect 11609 4777 11621 4780
rect 11655 4777 11667 4811
rect 12802 4808 12808 4820
rect 12763 4780 12808 4808
rect 11609 4771 11667 4777
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 13262 4768 13268 4820
rect 13320 4808 13326 4820
rect 13446 4808 13452 4820
rect 13320 4780 13452 4808
rect 13320 4768 13326 4780
rect 13446 4768 13452 4780
rect 13504 4768 13510 4820
rect 14090 4808 14096 4820
rect 14051 4780 14096 4808
rect 14090 4768 14096 4780
rect 14148 4768 14154 4820
rect 14458 4808 14464 4820
rect 14419 4780 14464 4808
rect 14458 4768 14464 4780
rect 14516 4768 14522 4820
rect 17402 4808 17408 4820
rect 17363 4780 17408 4808
rect 17402 4768 17408 4780
rect 17460 4768 17466 4820
rect 2032 4743 2090 4749
rect 2032 4709 2044 4743
rect 2078 4740 2090 4743
rect 2314 4740 2320 4752
rect 2078 4712 2320 4740
rect 2078 4709 2090 4712
rect 2032 4703 2090 4709
rect 2314 4700 2320 4712
rect 2372 4700 2378 4752
rect 5534 4700 5540 4752
rect 5592 4740 5598 4752
rect 5782 4743 5840 4749
rect 5782 4740 5794 4743
rect 5592 4712 5794 4740
rect 5592 4700 5598 4712
rect 5782 4709 5794 4712
rect 5828 4709 5840 4743
rect 5782 4703 5840 4709
rect 12710 4700 12716 4752
rect 12768 4740 12774 4752
rect 13173 4743 13231 4749
rect 13173 4740 13185 4743
rect 12768 4712 13185 4740
rect 12768 4700 12774 4712
rect 13173 4709 13185 4712
rect 13219 4709 13231 4743
rect 13173 4703 13231 4709
rect 14642 4700 14648 4752
rect 14700 4740 14706 4752
rect 18049 4743 18107 4749
rect 18049 4740 18061 4743
rect 14700 4712 18061 4740
rect 14700 4700 14706 4712
rect 18049 4709 18061 4712
rect 18095 4740 18107 4743
rect 18414 4740 18420 4752
rect 18095 4712 18420 4740
rect 18095 4709 18107 4712
rect 18049 4703 18107 4709
rect 18414 4700 18420 4712
rect 18472 4700 18478 4752
rect 4706 4632 4712 4684
rect 4764 4672 4770 4684
rect 8389 4675 8447 4681
rect 8389 4672 8401 4675
rect 4764 4644 8401 4672
rect 4764 4632 4770 4644
rect 8389 4641 8401 4644
rect 8435 4672 8447 4675
rect 8570 4672 8576 4684
rect 8435 4644 8576 4672
rect 8435 4641 8447 4644
rect 8389 4635 8447 4641
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 9398 4632 9404 4684
rect 9456 4672 9462 4684
rect 10045 4675 10103 4681
rect 10045 4672 10057 4675
rect 9456 4644 10057 4672
rect 9456 4632 9462 4644
rect 10045 4641 10057 4644
rect 10091 4641 10103 4675
rect 11701 4675 11759 4681
rect 11701 4672 11713 4675
rect 10045 4635 10103 4641
rect 11072 4644 11713 4672
rect 1762 4604 1768 4616
rect 1723 4576 1768 4604
rect 1762 4564 1768 4576
rect 1820 4564 1826 4616
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 4614 4604 4620 4616
rect 4387 4576 4620 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 4614 4564 4620 4576
rect 4672 4604 4678 4616
rect 4798 4604 4804 4616
rect 4672 4576 4804 4604
rect 4672 4564 4678 4576
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 5442 4564 5448 4616
rect 5500 4604 5506 4616
rect 5537 4607 5595 4613
rect 5537 4604 5549 4607
rect 5500 4576 5549 4604
rect 5500 4564 5506 4576
rect 5537 4573 5549 4576
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 8481 4607 8539 4613
rect 8481 4604 8493 4607
rect 8352 4576 8493 4604
rect 8352 4564 8358 4576
rect 8481 4573 8493 4576
rect 8527 4573 8539 4607
rect 8662 4604 8668 4616
rect 8623 4576 8668 4604
rect 8481 4567 8539 4573
rect 8662 4564 8668 4576
rect 8720 4564 8726 4616
rect 10134 4604 10140 4616
rect 10095 4576 10140 4604
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 10226 4564 10232 4616
rect 10284 4604 10290 4616
rect 10284 4576 10329 4604
rect 10284 4564 10290 4576
rect 4709 4539 4767 4545
rect 4709 4505 4721 4539
rect 4755 4536 4767 4539
rect 5460 4536 5488 4564
rect 11072 4545 11100 4644
rect 11701 4641 11713 4644
rect 11747 4641 11759 4675
rect 11701 4635 11759 4641
rect 13265 4675 13323 4681
rect 13265 4641 13277 4675
rect 13311 4672 13323 4675
rect 13446 4672 13452 4684
rect 13311 4644 13452 4672
rect 13311 4641 13323 4644
rect 13265 4635 13323 4641
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 16298 4681 16304 4684
rect 16292 4672 16304 4681
rect 16259 4644 16304 4672
rect 16292 4635 16304 4644
rect 16298 4632 16304 4635
rect 16356 4632 16362 4684
rect 18230 4672 18236 4684
rect 18191 4644 18236 4672
rect 18230 4632 18236 4644
rect 18288 4632 18294 4684
rect 19518 4672 19524 4684
rect 19479 4644 19524 4672
rect 19518 4632 19524 4644
rect 19576 4632 19582 4684
rect 20898 4672 20904 4684
rect 20859 4644 20904 4672
rect 20898 4632 20904 4644
rect 20956 4632 20962 4684
rect 22005 4675 22063 4681
rect 22005 4641 22017 4675
rect 22051 4672 22063 4675
rect 22051 4644 22085 4672
rect 22051 4641 22063 4644
rect 22005 4635 22063 4641
rect 11882 4604 11888 4616
rect 11843 4576 11888 4604
rect 11882 4564 11888 4576
rect 11940 4564 11946 4616
rect 12986 4564 12992 4616
rect 13044 4604 13050 4616
rect 13357 4607 13415 4613
rect 13357 4604 13369 4607
rect 13044 4576 13369 4604
rect 13044 4564 13050 4576
rect 13357 4573 13369 4576
rect 13403 4573 13415 4607
rect 16025 4607 16083 4613
rect 16025 4604 16037 4607
rect 13357 4567 13415 4573
rect 15856 4576 16037 4604
rect 4755 4508 5488 4536
rect 9677 4539 9735 4545
rect 4755 4505 4767 4508
rect 4709 4499 4767 4505
rect 9677 4505 9689 4539
rect 9723 4536 9735 4539
rect 11057 4539 11115 4545
rect 11057 4536 11069 4539
rect 9723 4508 11069 4536
rect 9723 4505 9735 4508
rect 9677 4499 9735 4505
rect 11057 4505 11069 4508
rect 11103 4505 11115 4539
rect 11057 4499 11115 4505
rect 1670 4468 1676 4480
rect 1631 4440 1676 4468
rect 1670 4428 1676 4440
rect 1728 4468 1734 4480
rect 5166 4468 5172 4480
rect 1728 4440 5172 4468
rect 1728 4428 1734 4440
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 7098 4428 7104 4480
rect 7156 4468 7162 4480
rect 7193 4471 7251 4477
rect 7193 4468 7205 4471
rect 7156 4440 7205 4468
rect 7156 4428 7162 4440
rect 7193 4437 7205 4440
rect 7239 4437 7251 4471
rect 7193 4431 7251 4437
rect 7282 4428 7288 4480
rect 7340 4468 7346 4480
rect 7561 4471 7619 4477
rect 7561 4468 7573 4471
rect 7340 4440 7573 4468
rect 7340 4428 7346 4440
rect 7561 4437 7573 4440
rect 7607 4437 7619 4471
rect 9398 4468 9404 4480
rect 9359 4440 9404 4468
rect 7561 4431 7619 4437
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 10778 4468 10784 4480
rect 10739 4440 10784 4468
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 11238 4468 11244 4480
rect 11199 4440 11244 4468
rect 11238 4428 11244 4440
rect 11296 4428 11302 4480
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 14829 4471 14887 4477
rect 12492 4440 12537 4468
rect 12492 4428 12498 4440
rect 14829 4437 14841 4471
rect 14875 4468 14887 4471
rect 15470 4468 15476 4480
rect 14875 4440 15476 4468
rect 14875 4437 14887 4440
rect 14829 4431 14887 4437
rect 15470 4428 15476 4440
rect 15528 4468 15534 4480
rect 15856 4477 15884 4576
rect 16025 4573 16037 4576
rect 16071 4573 16083 4607
rect 18506 4604 18512 4616
rect 18467 4576 18512 4604
rect 16025 4567 16083 4573
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 19797 4607 19855 4613
rect 19797 4573 19809 4607
rect 19843 4604 19855 4607
rect 22020 4604 22048 4635
rect 22186 4604 22192 4616
rect 19843 4576 22192 4604
rect 19843 4573 19855 4576
rect 19797 4567 19855 4573
rect 22186 4564 22192 4576
rect 22244 4564 22250 4616
rect 15841 4471 15899 4477
rect 15841 4468 15853 4471
rect 15528 4440 15853 4468
rect 15528 4428 15534 4440
rect 15841 4437 15853 4440
rect 15887 4437 15899 4471
rect 15841 4431 15899 4437
rect 21085 4471 21143 4477
rect 21085 4437 21097 4471
rect 21131 4468 21143 4471
rect 21542 4468 21548 4480
rect 21131 4440 21548 4468
rect 21131 4437 21143 4440
rect 21085 4431 21143 4437
rect 21542 4428 21548 4440
rect 21600 4428 21606 4480
rect 22094 4428 22100 4480
rect 22152 4468 22158 4480
rect 22189 4471 22247 4477
rect 22189 4468 22201 4471
rect 22152 4440 22201 4468
rect 22152 4428 22158 4440
rect 22189 4437 22201 4440
rect 22235 4437 22247 4471
rect 22189 4431 22247 4437
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1578 4264 1584 4276
rect 1539 4236 1584 4264
rect 1578 4224 1584 4236
rect 1636 4224 1642 4276
rect 2314 4224 2320 4276
rect 2372 4264 2378 4276
rect 2593 4267 2651 4273
rect 2593 4264 2605 4267
rect 2372 4236 2605 4264
rect 2372 4224 2378 4236
rect 2593 4233 2605 4236
rect 2639 4233 2651 4267
rect 2593 4227 2651 4233
rect 3053 4267 3111 4273
rect 3053 4233 3065 4267
rect 3099 4264 3111 4267
rect 3326 4264 3332 4276
rect 3099 4236 3332 4264
rect 3099 4233 3111 4236
rect 3053 4227 3111 4233
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 4798 4224 4804 4276
rect 4856 4264 4862 4276
rect 4893 4267 4951 4273
rect 4893 4264 4905 4267
rect 4856 4236 4905 4264
rect 4856 4224 4862 4236
rect 4893 4233 4905 4236
rect 4939 4264 4951 4267
rect 5442 4264 5448 4276
rect 4939 4236 5448 4264
rect 4939 4233 4951 4236
rect 4893 4227 4951 4233
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 7926 4264 7932 4276
rect 7887 4236 7932 4264
rect 7926 4224 7932 4236
rect 7984 4224 7990 4276
rect 8481 4267 8539 4273
rect 8481 4233 8493 4267
rect 8527 4264 8539 4267
rect 9398 4264 9404 4276
rect 8527 4236 9404 4264
rect 8527 4233 8539 4236
rect 8481 4227 8539 4233
rect 9398 4224 9404 4236
rect 9456 4224 9462 4276
rect 10778 4264 10784 4276
rect 10152 4236 10784 4264
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4128 2283 4131
rect 2332 4128 2360 4224
rect 6840 4168 7420 4196
rect 2271 4100 2360 4128
rect 2271 4097 2283 4100
rect 2225 4091 2283 4097
rect 4706 4088 4712 4140
rect 4764 4128 4770 4140
rect 6641 4131 6699 4137
rect 6641 4128 6653 4131
rect 4764 4100 6653 4128
rect 4764 4088 4770 4100
rect 6641 4097 6653 4100
rect 6687 4128 6699 4131
rect 6840 4128 6868 4168
rect 7282 4128 7288 4140
rect 6687 4100 6868 4128
rect 7243 4100 7288 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 7392 4137 7420 4168
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 9125 4131 9183 4137
rect 9125 4097 9137 4131
rect 9171 4128 9183 4131
rect 9398 4128 9404 4140
rect 9171 4100 9404 4128
rect 9171 4097 9183 4100
rect 9125 4091 9183 4097
rect 9398 4088 9404 4100
rect 9456 4088 9462 4140
rect 10152 4137 10180 4236
rect 10778 4224 10784 4236
rect 10836 4224 10842 4276
rect 15654 4224 15660 4276
rect 15712 4264 15718 4276
rect 17681 4267 17739 4273
rect 17681 4264 17693 4267
rect 15712 4236 17693 4264
rect 15712 4224 15718 4236
rect 17681 4233 17693 4236
rect 17727 4264 17739 4267
rect 17773 4267 17831 4273
rect 17773 4264 17785 4267
rect 17727 4236 17785 4264
rect 17727 4233 17739 4236
rect 17681 4227 17739 4233
rect 17773 4233 17785 4236
rect 17819 4233 17831 4267
rect 17773 4227 17831 4233
rect 18230 4224 18236 4276
rect 18288 4264 18294 4276
rect 19061 4267 19119 4273
rect 19061 4264 19073 4267
rect 18288 4236 19073 4264
rect 18288 4224 18294 4236
rect 19061 4233 19073 4236
rect 19107 4233 19119 4267
rect 19518 4264 19524 4276
rect 19479 4236 19524 4264
rect 19061 4227 19119 4233
rect 19518 4224 19524 4236
rect 19576 4224 19582 4276
rect 20809 4267 20867 4273
rect 20809 4233 20821 4267
rect 20855 4264 20867 4267
rect 20898 4264 20904 4276
rect 20855 4236 20904 4264
rect 20855 4233 20867 4236
rect 20809 4227 20867 4233
rect 17972 4168 18644 4196
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 12526 4088 12532 4140
rect 12584 4128 12590 4140
rect 13081 4131 13139 4137
rect 13081 4128 13093 4131
rect 12584 4100 13093 4128
rect 12584 4088 12590 4100
rect 13081 4097 13093 4100
rect 13127 4128 13139 4131
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13127 4100 13829 4128
rect 13127 4097 13139 4100
rect 13081 4091 13139 4097
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 17402 4128 17408 4140
rect 17363 4100 17408 4128
rect 13817 4091 13875 4097
rect 17402 4088 17408 4100
rect 17460 4128 17466 4140
rect 17972 4128 18000 4168
rect 18616 4137 18644 4168
rect 17460 4100 18000 4128
rect 18601 4131 18659 4137
rect 17460 4088 17466 4100
rect 18601 4097 18613 4131
rect 18647 4097 18659 4131
rect 18601 4091 18659 4097
rect 19889 4131 19947 4137
rect 19889 4097 19901 4131
rect 19935 4128 19947 4131
rect 20824 4128 20852 4227
rect 20898 4224 20904 4236
rect 20956 4224 20962 4276
rect 19935 4100 20852 4128
rect 19935 4097 19947 4100
rect 19889 4091 19947 4097
rect 22186 4088 22192 4140
rect 22244 4128 22250 4140
rect 22557 4131 22615 4137
rect 22557 4128 22569 4131
rect 22244 4100 22569 4128
rect 22244 4088 22250 4100
rect 22557 4097 22569 4100
rect 22603 4097 22615 4131
rect 22557 4091 22615 4097
rect 3145 4063 3203 4069
rect 3145 4029 3157 4063
rect 3191 4060 3203 4063
rect 4798 4060 4804 4072
rect 3191 4032 4804 4060
rect 3191 4029 3203 4032
rect 3145 4023 3203 4029
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 5994 4060 6000 4072
rect 5955 4032 6000 4060
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 6822 4020 6828 4072
rect 6880 4060 6886 4072
rect 7193 4063 7251 4069
rect 7193 4060 7205 4063
rect 6880 4032 7205 4060
rect 6880 4020 6886 4032
rect 7193 4029 7205 4032
rect 7239 4029 7251 4063
rect 7193 4023 7251 4029
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 8849 4063 8907 4069
rect 8849 4060 8861 4063
rect 7984 4032 8861 4060
rect 7984 4020 7990 4032
rect 8849 4029 8861 4032
rect 8895 4060 8907 4063
rect 10404 4063 10462 4069
rect 8895 4032 10364 4060
rect 8895 4029 8907 4032
rect 8849 4023 8907 4029
rect 1210 3952 1216 4004
rect 1268 3992 1274 4004
rect 1670 3992 1676 4004
rect 1268 3964 1676 3992
rect 1268 3952 1274 3964
rect 1670 3952 1676 3964
rect 1728 3992 1734 4004
rect 1949 3995 2007 4001
rect 1949 3992 1961 3995
rect 1728 3964 1961 3992
rect 1728 3952 1734 3964
rect 1949 3961 1961 3964
rect 1995 3961 2007 3995
rect 1949 3955 2007 3961
rect 3326 3952 3332 4004
rect 3384 4001 3390 4004
rect 3384 3995 3448 4001
rect 3384 3961 3402 3995
rect 3436 3961 3448 3995
rect 3384 3955 3448 3961
rect 3384 3952 3390 3955
rect 4338 3952 4344 4004
rect 4396 3992 4402 4004
rect 5166 3992 5172 4004
rect 4396 3964 5172 3992
rect 4396 3952 4402 3964
rect 5166 3952 5172 3964
rect 5224 3952 5230 4004
rect 8110 3952 8116 4004
rect 8168 3992 8174 4004
rect 8389 3995 8447 4001
rect 8389 3992 8401 3995
rect 8168 3964 8401 3992
rect 8168 3952 8174 3964
rect 8389 3961 8401 3964
rect 8435 3992 8447 3995
rect 8435 3964 8984 3992
rect 8435 3961 8447 3964
rect 8389 3955 8447 3961
rect 4525 3927 4583 3933
rect 4525 3893 4537 3927
rect 4571 3924 4583 3927
rect 4614 3924 4620 3936
rect 4571 3896 4620 3924
rect 4571 3893 4583 3896
rect 4525 3887 4583 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 5442 3884 5448 3936
rect 5500 3924 5506 3936
rect 5537 3927 5595 3933
rect 5537 3924 5549 3927
rect 5500 3896 5549 3924
rect 5500 3884 5506 3896
rect 5537 3893 5549 3896
rect 5583 3893 5595 3927
rect 5537 3887 5595 3893
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 8956 3933 8984 3964
rect 9030 3952 9036 4004
rect 9088 3992 9094 4004
rect 9953 3995 10011 4001
rect 9953 3992 9965 3995
rect 9088 3964 9965 3992
rect 9088 3952 9094 3964
rect 9953 3961 9965 3964
rect 9999 3992 10011 3995
rect 10226 3992 10232 4004
rect 9999 3964 10232 3992
rect 9999 3961 10011 3964
rect 9953 3955 10011 3961
rect 10226 3952 10232 3964
rect 10284 3952 10290 4004
rect 10336 3992 10364 4032
rect 10404 4029 10416 4063
rect 10450 4060 10462 4063
rect 10686 4060 10692 4072
rect 10450 4032 10692 4060
rect 10450 4029 10462 4032
rect 10404 4023 10462 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 11072 4032 12173 4060
rect 11072 3992 11100 4032
rect 12161 4029 12173 4032
rect 12207 4029 12219 4063
rect 12161 4023 12219 4029
rect 10336 3964 11100 3992
rect 11330 3952 11336 4004
rect 11388 3992 11394 4004
rect 11793 3995 11851 4001
rect 11793 3992 11805 3995
rect 11388 3964 11805 3992
rect 11388 3952 11394 3964
rect 11793 3961 11805 3964
rect 11839 3992 11851 3995
rect 11882 3992 11888 4004
rect 11839 3964 11888 3992
rect 11839 3961 11851 3964
rect 11793 3955 11851 3961
rect 11882 3952 11888 3964
rect 11940 3952 11946 4004
rect 12176 3992 12204 4023
rect 12434 4020 12440 4072
rect 12492 4060 12498 4072
rect 12805 4063 12863 4069
rect 12805 4060 12817 4063
rect 12492 4032 12817 4060
rect 12492 4020 12498 4032
rect 12805 4029 12817 4032
rect 12851 4029 12863 4063
rect 14093 4063 14151 4069
rect 14093 4060 14105 4063
rect 12805 4023 12863 4029
rect 13832 4032 14105 4060
rect 13832 4004 13860 4032
rect 14093 4029 14105 4032
rect 14139 4060 14151 4063
rect 14829 4063 14887 4069
rect 14829 4060 14841 4063
rect 14139 4032 14841 4060
rect 14139 4029 14151 4032
rect 14093 4023 14151 4029
rect 14829 4029 14841 4032
rect 14875 4029 14887 4063
rect 14829 4023 14887 4029
rect 15381 4063 15439 4069
rect 15381 4029 15393 4063
rect 15427 4060 15439 4063
rect 15470 4060 15476 4072
rect 15427 4032 15476 4060
rect 15427 4029 15439 4032
rect 15381 4023 15439 4029
rect 15470 4020 15476 4032
rect 15528 4020 15534 4072
rect 17681 4063 17739 4069
rect 17681 4029 17693 4063
rect 17727 4060 17739 4063
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 17727 4032 18521 4060
rect 17727 4029 17739 4032
rect 17681 4023 17739 4029
rect 18509 4029 18521 4032
rect 18555 4029 18567 4063
rect 18509 4023 18567 4029
rect 19518 4020 19524 4072
rect 19576 4060 19582 4072
rect 19613 4063 19671 4069
rect 19613 4060 19625 4063
rect 19576 4032 19625 4060
rect 19576 4020 19582 4032
rect 19613 4029 19625 4032
rect 19659 4060 19671 4063
rect 20349 4063 20407 4069
rect 20349 4060 20361 4063
rect 19659 4032 20361 4060
rect 19659 4029 19671 4032
rect 19613 4023 19671 4029
rect 20349 4029 20361 4032
rect 20395 4029 20407 4063
rect 20898 4060 20904 4072
rect 20859 4032 20904 4060
rect 20349 4023 20407 4029
rect 20898 4020 20904 4032
rect 20956 4060 20962 4072
rect 21453 4063 21511 4069
rect 21453 4060 21465 4063
rect 20956 4032 21465 4060
rect 20956 4020 20962 4032
rect 21453 4029 21465 4032
rect 21499 4029 21511 4063
rect 22005 4063 22063 4069
rect 22005 4060 22017 4063
rect 21453 4023 21511 4029
rect 21836 4032 22017 4060
rect 12897 3995 12955 4001
rect 12897 3992 12909 3995
rect 12176 3964 12909 3992
rect 12897 3961 12909 3964
rect 12943 3961 12955 3995
rect 12897 3955 12955 3961
rect 13814 3952 13820 4004
rect 13872 3952 13878 4004
rect 14369 3995 14427 4001
rect 14369 3961 14381 3995
rect 14415 3992 14427 3995
rect 15102 3992 15108 4004
rect 14415 3964 15108 3992
rect 14415 3961 14427 3964
rect 14369 3955 14427 3961
rect 15102 3952 15108 3964
rect 15160 3952 15166 4004
rect 15626 3995 15684 4001
rect 15626 3992 15638 3995
rect 15304 3964 15638 3992
rect 15304 3936 15332 3964
rect 15626 3961 15638 3964
rect 15672 3961 15684 3995
rect 17129 3995 17187 4001
rect 17129 3992 17141 3995
rect 15626 3955 15684 3961
rect 16776 3964 17141 3992
rect 6825 3927 6883 3933
rect 6825 3924 6837 3927
rect 6788 3896 6837 3924
rect 6788 3884 6794 3896
rect 6825 3893 6837 3896
rect 6871 3893 6883 3927
rect 6825 3887 6883 3893
rect 8941 3927 8999 3933
rect 8941 3893 8953 3927
rect 8987 3924 8999 3927
rect 9122 3924 9128 3936
rect 8987 3896 9128 3924
rect 8987 3893 8999 3896
rect 8941 3887 8999 3893
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 9493 3927 9551 3933
rect 9493 3924 9505 3927
rect 9456 3896 9505 3924
rect 9456 3884 9462 3896
rect 9493 3893 9505 3896
rect 9539 3893 9551 3927
rect 11514 3924 11520 3936
rect 11475 3896 11520 3924
rect 9493 3887 9551 3893
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 13446 3924 13452 3936
rect 12492 3896 12537 3924
rect 13407 3896 13452 3924
rect 12492 3884 12498 3896
rect 13446 3884 13452 3896
rect 13504 3884 13510 3936
rect 15286 3924 15292 3936
rect 15247 3896 15292 3924
rect 15286 3884 15292 3896
rect 15344 3884 15350 3936
rect 16298 3884 16304 3936
rect 16356 3924 16362 3936
rect 16666 3924 16672 3936
rect 16356 3896 16672 3924
rect 16356 3884 16362 3896
rect 16666 3884 16672 3896
rect 16724 3924 16730 3936
rect 16776 3933 16804 3964
rect 17129 3961 17141 3964
rect 17175 3992 17187 3995
rect 18138 3992 18144 4004
rect 17175 3964 18144 3992
rect 17175 3961 17187 3964
rect 17129 3955 17187 3961
rect 18138 3952 18144 3964
rect 18196 3952 18202 4004
rect 18414 3992 18420 4004
rect 18375 3964 18420 3992
rect 18414 3952 18420 3964
rect 18472 3952 18478 4004
rect 21836 3936 21864 4032
rect 22005 4029 22017 4032
rect 22051 4029 22063 4063
rect 22005 4023 22063 4029
rect 23198 3992 23204 4004
rect 22204 3964 23204 3992
rect 16761 3927 16819 3933
rect 16761 3924 16773 3927
rect 16724 3896 16773 3924
rect 16724 3884 16730 3896
rect 16761 3893 16773 3896
rect 16807 3893 16819 3927
rect 16761 3887 16819 3893
rect 18049 3927 18107 3933
rect 18049 3893 18061 3927
rect 18095 3924 18107 3927
rect 18322 3924 18328 3936
rect 18095 3896 18328 3924
rect 18095 3893 18107 3896
rect 18049 3887 18107 3893
rect 18322 3884 18328 3896
rect 18380 3884 18386 3936
rect 19978 3884 19984 3936
rect 20036 3924 20042 3936
rect 21085 3927 21143 3933
rect 21085 3924 21097 3927
rect 20036 3896 21097 3924
rect 20036 3884 20042 3896
rect 21085 3893 21097 3896
rect 21131 3893 21143 3927
rect 21818 3924 21824 3936
rect 21779 3896 21824 3924
rect 21085 3887 21143 3893
rect 21818 3884 21824 3896
rect 21876 3884 21882 3936
rect 22204 3933 22232 3964
rect 23198 3952 23204 3964
rect 23256 3952 23262 4004
rect 22189 3927 22247 3933
rect 22189 3893 22201 3927
rect 22235 3893 22247 3927
rect 22189 3887 22247 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 198 3680 204 3732
rect 256 3720 262 3732
rect 1673 3723 1731 3729
rect 1673 3720 1685 3723
rect 256 3692 1685 3720
rect 256 3680 262 3692
rect 1673 3689 1685 3692
rect 1719 3720 1731 3723
rect 2038 3720 2044 3732
rect 1719 3692 2044 3720
rect 1719 3689 1731 3692
rect 1673 3683 1731 3689
rect 2038 3680 2044 3692
rect 2096 3680 2102 3732
rect 2314 3680 2320 3732
rect 2372 3720 2378 3732
rect 3145 3723 3203 3729
rect 3145 3720 3157 3723
rect 2372 3692 3157 3720
rect 2372 3680 2378 3692
rect 3145 3689 3157 3692
rect 3191 3720 3203 3723
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 3191 3692 3433 3720
rect 3191 3689 3203 3692
rect 3145 3683 3203 3689
rect 3421 3689 3433 3692
rect 3467 3689 3479 3723
rect 4706 3720 4712 3732
rect 4667 3692 4712 3720
rect 3421 3683 3479 3689
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 5166 3680 5172 3732
rect 5224 3720 5230 3732
rect 5537 3723 5595 3729
rect 5537 3720 5549 3723
rect 5224 3692 5549 3720
rect 5224 3680 5230 3692
rect 5537 3689 5549 3692
rect 5583 3689 5595 3723
rect 5537 3683 5595 3689
rect 6733 3723 6791 3729
rect 6733 3689 6745 3723
rect 6779 3720 6791 3723
rect 7282 3720 7288 3732
rect 6779 3692 7288 3720
rect 6779 3689 6791 3692
rect 6733 3683 6791 3689
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 8110 3720 8116 3732
rect 8071 3692 8116 3720
rect 8110 3680 8116 3692
rect 8168 3720 8174 3732
rect 8294 3720 8300 3732
rect 8168 3692 8300 3720
rect 8168 3680 8174 3692
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 8481 3723 8539 3729
rect 8481 3689 8493 3723
rect 8527 3720 8539 3723
rect 8570 3720 8576 3732
rect 8527 3692 8576 3720
rect 8527 3689 8539 3692
rect 8481 3683 8539 3689
rect 8570 3680 8576 3692
rect 8628 3680 8634 3732
rect 9493 3723 9551 3729
rect 9493 3689 9505 3723
rect 9539 3720 9551 3723
rect 10134 3720 10140 3732
rect 9539 3692 10140 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 10686 3720 10692 3732
rect 10647 3692 10692 3720
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 11054 3720 11060 3732
rect 11015 3692 11060 3720
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 12526 3720 12532 3732
rect 12487 3692 12532 3720
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 12710 3680 12716 3732
rect 12768 3720 12774 3732
rect 12805 3723 12863 3729
rect 12805 3720 12817 3723
rect 12768 3692 12817 3720
rect 12768 3680 12774 3692
rect 12805 3689 12817 3692
rect 12851 3689 12863 3723
rect 12805 3683 12863 3689
rect 12986 3680 12992 3732
rect 13044 3720 13050 3732
rect 13173 3723 13231 3729
rect 13173 3720 13185 3723
rect 13044 3692 13185 3720
rect 13044 3680 13050 3692
rect 13173 3689 13185 3692
rect 13219 3689 13231 3723
rect 13173 3683 13231 3689
rect 13722 3680 13728 3732
rect 13780 3720 13786 3732
rect 13817 3723 13875 3729
rect 13817 3720 13829 3723
rect 13780 3692 13829 3720
rect 13780 3680 13786 3692
rect 13817 3689 13829 3692
rect 13863 3689 13875 3723
rect 13817 3683 13875 3689
rect 15933 3723 15991 3729
rect 15933 3689 15945 3723
rect 15979 3720 15991 3723
rect 16022 3720 16028 3732
rect 15979 3692 16028 3720
rect 15979 3689 15991 3692
rect 15933 3683 15991 3689
rect 16022 3680 16028 3692
rect 16080 3680 16086 3732
rect 16206 3680 16212 3732
rect 16264 3720 16270 3732
rect 16301 3723 16359 3729
rect 16301 3720 16313 3723
rect 16264 3692 16313 3720
rect 16264 3680 16270 3692
rect 16301 3689 16313 3692
rect 16347 3689 16359 3723
rect 16301 3683 16359 3689
rect 16574 3680 16580 3732
rect 16632 3720 16638 3732
rect 17497 3723 17555 3729
rect 17497 3720 17509 3723
rect 16632 3692 17509 3720
rect 16632 3680 16638 3692
rect 17497 3689 17509 3692
rect 17543 3689 17555 3723
rect 17862 3720 17868 3732
rect 17823 3692 17868 3720
rect 17497 3683 17555 3689
rect 17862 3680 17868 3692
rect 17920 3680 17926 3732
rect 18322 3680 18328 3732
rect 18380 3720 18386 3732
rect 18877 3723 18935 3729
rect 18877 3720 18889 3723
rect 18380 3692 18889 3720
rect 18380 3680 18386 3692
rect 18877 3689 18889 3692
rect 18923 3689 18935 3723
rect 18877 3683 18935 3689
rect 5077 3655 5135 3661
rect 5077 3621 5089 3655
rect 5123 3652 5135 3655
rect 6641 3655 6699 3661
rect 5123 3624 5672 3652
rect 5123 3621 5135 3624
rect 5077 3615 5135 3621
rect 1762 3584 1768 3596
rect 1723 3556 1768 3584
rect 1762 3544 1768 3556
rect 1820 3544 1826 3596
rect 2038 3593 2044 3596
rect 2032 3584 2044 3593
rect 1999 3556 2044 3584
rect 2032 3547 2044 3556
rect 2038 3544 2044 3547
rect 2096 3544 2102 3596
rect 5644 3593 5672 3624
rect 6641 3621 6653 3655
rect 6687 3652 6699 3655
rect 6822 3652 6828 3664
rect 6687 3624 6828 3652
rect 6687 3621 6699 3624
rect 6641 3615 6699 3621
rect 6822 3612 6828 3624
rect 6880 3612 6886 3664
rect 7006 3612 7012 3664
rect 7064 3652 7070 3664
rect 7101 3655 7159 3661
rect 7101 3652 7113 3655
rect 7064 3624 7113 3652
rect 7064 3612 7070 3624
rect 7101 3621 7113 3624
rect 7147 3621 7159 3655
rect 7101 3615 7159 3621
rect 11416 3655 11474 3661
rect 11416 3621 11428 3655
rect 11462 3652 11474 3655
rect 11514 3652 11520 3664
rect 11462 3624 11520 3652
rect 11462 3621 11474 3624
rect 11416 3615 11474 3621
rect 11514 3612 11520 3624
rect 11572 3612 11578 3664
rect 14734 3612 14740 3664
rect 14792 3652 14798 3664
rect 16390 3652 16396 3664
rect 14792 3624 16396 3652
rect 14792 3612 14798 3624
rect 16390 3612 16396 3624
rect 16448 3612 16454 3664
rect 19337 3655 19395 3661
rect 19337 3621 19349 3655
rect 19383 3652 19395 3655
rect 19426 3652 19432 3664
rect 19383 3624 19432 3652
rect 19383 3621 19395 3624
rect 19337 3615 19395 3621
rect 19426 3612 19432 3624
rect 19484 3612 19490 3664
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3584 5687 3587
rect 6730 3584 6736 3596
rect 5675 3556 6736 3584
rect 5675 3553 5687 3556
rect 5629 3547 5687 3553
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 7190 3584 7196 3596
rect 7151 3556 7196 3584
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 9766 3544 9772 3596
rect 9824 3584 9830 3596
rect 9861 3587 9919 3593
rect 9861 3584 9873 3587
rect 9824 3556 9873 3584
rect 9824 3544 9830 3556
rect 9861 3553 9873 3556
rect 9907 3553 9919 3587
rect 9861 3547 9919 3553
rect 10778 3544 10784 3596
rect 10836 3584 10842 3596
rect 11149 3587 11207 3593
rect 11149 3584 11161 3587
rect 10836 3556 11161 3584
rect 10836 3544 10842 3556
rect 11149 3553 11161 3556
rect 11195 3584 11207 3587
rect 12342 3584 12348 3596
rect 11195 3556 12348 3584
rect 11195 3553 11207 3556
rect 11149 3547 11207 3553
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 12618 3544 12624 3596
rect 12676 3584 12682 3596
rect 13725 3587 13783 3593
rect 13725 3584 13737 3587
rect 12676 3556 13737 3584
rect 12676 3544 12682 3556
rect 13725 3553 13737 3556
rect 13771 3584 13783 3587
rect 14458 3584 14464 3596
rect 13771 3556 14464 3584
rect 13771 3553 13783 3556
rect 13725 3547 13783 3553
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 19058 3584 19064 3596
rect 19019 3556 19064 3584
rect 19058 3544 19064 3556
rect 19116 3544 19122 3596
rect 20898 3584 20904 3596
rect 20859 3556 20904 3584
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 22002 3584 22008 3596
rect 21963 3556 22008 3584
rect 22002 3544 22008 3556
rect 22060 3544 22066 3596
rect 23934 3584 23940 3596
rect 23895 3556 23940 3584
rect 23934 3544 23940 3556
rect 23992 3544 23998 3596
rect 3326 3476 3332 3528
rect 3384 3516 3390 3528
rect 4157 3519 4215 3525
rect 4157 3516 4169 3519
rect 3384 3488 4169 3516
rect 3384 3476 3390 3488
rect 4157 3485 4169 3488
rect 4203 3485 4215 3519
rect 4157 3479 4215 3485
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 5500 3488 5733 3516
rect 5500 3476 5506 3488
rect 5721 3485 5733 3488
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 7285 3519 7343 3525
rect 7285 3485 7297 3519
rect 7331 3485 7343 3519
rect 7285 3479 7343 3485
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3516 8631 3519
rect 9582 3516 9588 3528
rect 8619 3488 9588 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 7098 3408 7104 3460
rect 7156 3448 7162 3460
rect 7300 3448 7328 3479
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 10134 3516 10140 3528
rect 10095 3488 10140 3516
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 14001 3519 14059 3525
rect 14001 3485 14013 3519
rect 14047 3516 14059 3519
rect 16577 3519 16635 3525
rect 14047 3488 14228 3516
rect 14047 3485 14059 3488
rect 14001 3479 14059 3485
rect 7156 3420 7328 3448
rect 7156 3408 7162 3420
rect 14200 3392 14228 3488
rect 16577 3485 16589 3519
rect 16623 3516 16635 3519
rect 16666 3516 16672 3528
rect 16623 3488 16672 3516
rect 16623 3485 16635 3488
rect 16577 3479 16635 3485
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 17770 3476 17776 3528
rect 17828 3516 17834 3528
rect 17957 3519 18015 3525
rect 17957 3516 17969 3519
rect 17828 3488 17969 3516
rect 17828 3476 17834 3488
rect 17957 3485 17969 3488
rect 18003 3485 18015 3519
rect 18138 3516 18144 3528
rect 18099 3488 18144 3516
rect 17957 3479 18015 3485
rect 18138 3476 18144 3488
rect 18196 3476 18202 3528
rect 16942 3448 16948 3460
rect 16903 3420 16948 3448
rect 16942 3408 16948 3420
rect 17000 3408 17006 3460
rect 3510 3340 3516 3392
rect 3568 3380 3574 3392
rect 3789 3383 3847 3389
rect 3789 3380 3801 3383
rect 3568 3352 3801 3380
rect 3568 3340 3574 3352
rect 3789 3349 3801 3352
rect 3835 3349 3847 3383
rect 3789 3343 3847 3349
rect 4430 3340 4436 3392
rect 4488 3380 4494 3392
rect 4798 3380 4804 3392
rect 4488 3352 4804 3380
rect 4488 3340 4494 3352
rect 4798 3340 4804 3352
rect 4856 3340 4862 3392
rect 5166 3380 5172 3392
rect 5127 3352 5172 3380
rect 5166 3340 5172 3352
rect 5224 3340 5230 3392
rect 6273 3383 6331 3389
rect 6273 3349 6285 3383
rect 6319 3380 6331 3383
rect 7466 3380 7472 3392
rect 6319 3352 7472 3380
rect 6319 3349 6331 3352
rect 6273 3343 6331 3349
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 8662 3340 8668 3392
rect 8720 3380 8726 3392
rect 9033 3383 9091 3389
rect 9033 3380 9045 3383
rect 8720 3352 9045 3380
rect 8720 3340 8726 3352
rect 9033 3349 9045 3352
rect 9079 3380 9091 3383
rect 9398 3380 9404 3392
rect 9079 3352 9404 3380
rect 9079 3349 9091 3352
rect 9033 3343 9091 3349
rect 9398 3340 9404 3352
rect 9456 3380 9462 3392
rect 9950 3380 9956 3392
rect 9456 3352 9956 3380
rect 9456 3340 9462 3352
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 13357 3383 13415 3389
rect 13357 3349 13369 3383
rect 13403 3380 13415 3383
rect 13630 3380 13636 3392
rect 13403 3352 13636 3380
rect 13403 3349 13415 3352
rect 13357 3343 13415 3349
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 14182 3340 14188 3392
rect 14240 3380 14246 3392
rect 14369 3383 14427 3389
rect 14369 3380 14381 3383
rect 14240 3352 14381 3380
rect 14240 3340 14246 3352
rect 14369 3349 14381 3352
rect 14415 3380 14427 3383
rect 14737 3383 14795 3389
rect 14737 3380 14749 3383
rect 14415 3352 14749 3380
rect 14415 3349 14427 3352
rect 14369 3343 14427 3349
rect 14737 3349 14749 3352
rect 14783 3349 14795 3383
rect 15470 3380 15476 3392
rect 15431 3352 15476 3380
rect 14737 3343 14795 3349
rect 15470 3340 15476 3352
rect 15528 3380 15534 3392
rect 17313 3383 17371 3389
rect 17313 3380 17325 3383
rect 15528 3352 17325 3380
rect 15528 3340 15534 3352
rect 17313 3349 17325 3352
rect 17359 3349 17371 3383
rect 18598 3380 18604 3392
rect 18559 3352 18604 3380
rect 17313 3343 17371 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 21082 3380 21088 3392
rect 21043 3352 21088 3380
rect 21082 3340 21088 3352
rect 21140 3340 21146 3392
rect 22186 3380 22192 3392
rect 22147 3352 22192 3380
rect 22186 3340 22192 3352
rect 22244 3340 22250 3392
rect 24118 3380 24124 3392
rect 24079 3352 24124 3380
rect 24118 3340 24124 3352
rect 24176 3340 24182 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1397 3179 1455 3185
rect 1397 3145 1409 3179
rect 1443 3176 1455 3179
rect 1486 3176 1492 3188
rect 1443 3148 1492 3176
rect 1443 3145 1455 3148
rect 1397 3139 1455 3145
rect 1486 3136 1492 3148
rect 1544 3136 1550 3188
rect 2222 3136 2228 3188
rect 2280 3176 2286 3188
rect 2409 3179 2467 3185
rect 2409 3176 2421 3179
rect 2280 3148 2421 3176
rect 2280 3136 2286 3148
rect 2409 3145 2421 3148
rect 2455 3145 2467 3179
rect 2409 3139 2467 3145
rect 2961 3179 3019 3185
rect 2961 3145 2973 3179
rect 3007 3176 3019 3179
rect 4338 3176 4344 3188
rect 3007 3148 4344 3176
rect 3007 3145 3019 3148
rect 2961 3139 3019 3145
rect 4338 3136 4344 3148
rect 4396 3136 4402 3188
rect 4433 3179 4491 3185
rect 4433 3145 4445 3179
rect 4479 3176 4491 3179
rect 5442 3176 5448 3188
rect 4479 3148 5448 3176
rect 4479 3145 4491 3148
rect 4433 3139 4491 3145
rect 5442 3136 5448 3148
rect 5500 3176 5506 3188
rect 5905 3179 5963 3185
rect 5905 3176 5917 3179
rect 5500 3148 5917 3176
rect 5500 3136 5506 3148
rect 5905 3145 5917 3148
rect 5951 3145 5963 3179
rect 5905 3139 5963 3145
rect 6641 3179 6699 3185
rect 6641 3145 6653 3179
rect 6687 3176 6699 3179
rect 7190 3176 7196 3188
rect 6687 3148 7196 3176
rect 6687 3145 6699 3148
rect 6641 3139 6699 3145
rect 7190 3136 7196 3148
rect 7248 3136 7254 3188
rect 10226 3136 10232 3188
rect 10284 3176 10290 3188
rect 10413 3179 10471 3185
rect 10413 3176 10425 3179
rect 10284 3148 10425 3176
rect 10284 3136 10290 3148
rect 10413 3145 10425 3148
rect 10459 3145 10471 3179
rect 12434 3176 12440 3188
rect 10413 3139 10471 3145
rect 11808 3148 12440 3176
rect 8202 3108 8208 3120
rect 7208 3080 8208 3108
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 1946 3040 1952 3052
rect 1903 3012 1952 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3040 2099 3043
rect 3510 3040 3516 3052
rect 2087 3012 3516 3040
rect 2087 3009 2099 3012
rect 2041 3003 2099 3009
rect 3510 3000 3516 3012
rect 3568 3000 3574 3052
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3040 3663 3043
rect 3651 3012 4200 3040
rect 3651 3009 3663 3012
rect 3605 3003 3663 3009
rect 1765 2975 1823 2981
rect 1765 2941 1777 2975
rect 1811 2972 1823 2975
rect 2222 2972 2228 2984
rect 1811 2944 2228 2972
rect 1811 2941 1823 2944
rect 1765 2935 1823 2941
rect 2222 2932 2228 2944
rect 2280 2932 2286 2984
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2972 2927 2975
rect 3326 2972 3332 2984
rect 2915 2944 3332 2972
rect 2915 2941 2927 2944
rect 2869 2935 2927 2941
rect 3326 2932 3332 2944
rect 3384 2932 3390 2984
rect 3421 2975 3479 2981
rect 3421 2941 3433 2975
rect 3467 2972 3479 2975
rect 4062 2972 4068 2984
rect 3467 2944 4068 2972
rect 3467 2941 3479 2944
rect 3421 2935 3479 2941
rect 4062 2932 4068 2944
rect 4120 2932 4126 2984
rect 3973 2907 4031 2913
rect 3973 2873 3985 2907
rect 4019 2904 4031 2907
rect 4172 2904 4200 3012
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 7208 3049 7236 3080
rect 8202 3068 8208 3080
rect 8260 3068 8266 3120
rect 9398 3068 9404 3120
rect 9456 3108 9462 3120
rect 9585 3111 9643 3117
rect 9585 3108 9597 3111
rect 9456 3080 9597 3108
rect 9456 3068 9462 3080
rect 9585 3077 9597 3080
rect 9631 3077 9643 3111
rect 9950 3108 9956 3120
rect 9863 3080 9956 3108
rect 9585 3071 9643 3077
rect 9950 3068 9956 3080
rect 10008 3108 10014 3120
rect 11514 3108 11520 3120
rect 10008 3080 11008 3108
rect 11475 3080 11520 3108
rect 10008 3068 10014 3080
rect 10980 3052 11008 3080
rect 11514 3068 11520 3080
rect 11572 3068 11578 3120
rect 4525 3043 4583 3049
rect 4525 3040 4537 3043
rect 4488 3012 4537 3040
rect 4488 3000 4494 3012
rect 4525 3009 4537 3012
rect 4571 3009 4583 3043
rect 4525 3003 4583 3009
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3040 8171 3043
rect 10870 3040 10876 3052
rect 8159 3012 8340 3040
rect 10831 3012 10876 3040
rect 8159 3009 8171 3012
rect 8113 3003 8171 3009
rect 4614 2932 4620 2984
rect 4672 2972 4678 2984
rect 6181 2975 6239 2981
rect 6181 2972 6193 2975
rect 4672 2944 6193 2972
rect 4672 2932 4678 2944
rect 6181 2941 6193 2944
rect 6227 2972 6239 2975
rect 7098 2972 7104 2984
rect 6227 2944 7104 2972
rect 6227 2941 6239 2944
rect 6181 2935 6239 2941
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 7466 2932 7472 2984
rect 7524 2972 7530 2984
rect 7745 2975 7803 2981
rect 7745 2972 7757 2975
rect 7524 2944 7757 2972
rect 7524 2932 7530 2944
rect 7745 2941 7757 2944
rect 7791 2972 7803 2975
rect 8205 2975 8263 2981
rect 8205 2972 8217 2975
rect 7791 2944 8217 2972
rect 7791 2941 7803 2944
rect 7745 2935 7803 2941
rect 8205 2941 8217 2944
rect 8251 2941 8263 2975
rect 8312 2972 8340 3012
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 10962 3000 10968 3052
rect 11020 3040 11026 3052
rect 11020 3012 11065 3040
rect 11020 3000 11026 3012
rect 8472 2975 8530 2981
rect 8472 2972 8484 2975
rect 8312 2944 8484 2972
rect 8205 2935 8263 2941
rect 8472 2941 8484 2944
rect 8518 2972 8530 2975
rect 9030 2972 9036 2984
rect 8518 2944 9036 2972
rect 8518 2941 8530 2944
rect 8472 2935 8530 2941
rect 4706 2904 4712 2916
rect 4019 2876 4712 2904
rect 4019 2873 4031 2876
rect 3973 2867 4031 2873
rect 4706 2864 4712 2876
rect 4764 2913 4770 2916
rect 4764 2907 4828 2913
rect 4764 2873 4782 2907
rect 4816 2904 4828 2907
rect 5718 2904 5724 2916
rect 4816 2876 5724 2904
rect 4816 2873 4828 2876
rect 4764 2867 4828 2873
rect 4764 2864 4770 2867
rect 5718 2864 5724 2876
rect 5776 2864 5782 2916
rect 8220 2904 8248 2935
rect 9030 2932 9036 2944
rect 9088 2932 9094 2984
rect 11422 2932 11428 2984
rect 11480 2972 11486 2984
rect 11808 2981 11836 3148
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 13722 3136 13728 3188
rect 13780 3176 13786 3188
rect 14093 3179 14151 3185
rect 14093 3176 14105 3179
rect 13780 3148 14105 3176
rect 13780 3136 13786 3148
rect 14093 3145 14105 3148
rect 14139 3145 14151 3179
rect 14458 3176 14464 3188
rect 14419 3148 14464 3176
rect 14093 3139 14151 3145
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 16206 3136 16212 3188
rect 16264 3176 16270 3188
rect 16669 3179 16727 3185
rect 16669 3176 16681 3179
rect 16264 3148 16681 3176
rect 16264 3136 16270 3148
rect 16669 3145 16681 3148
rect 16715 3145 16727 3179
rect 16669 3139 16727 3145
rect 17589 3179 17647 3185
rect 17589 3145 17601 3179
rect 17635 3176 17647 3179
rect 17862 3176 17868 3188
rect 17635 3148 17868 3176
rect 17635 3145 17647 3148
rect 17589 3139 17647 3145
rect 17862 3136 17868 3148
rect 17920 3136 17926 3188
rect 18046 3176 18052 3188
rect 18007 3148 18052 3176
rect 18046 3136 18052 3148
rect 18104 3136 18110 3188
rect 18138 3136 18144 3188
rect 18196 3176 18202 3188
rect 19061 3179 19119 3185
rect 19061 3176 19073 3179
rect 18196 3148 19073 3176
rect 18196 3136 18202 3148
rect 19061 3145 19073 3148
rect 19107 3145 19119 3179
rect 21358 3176 21364 3188
rect 21319 3148 21364 3176
rect 19061 3139 19119 3145
rect 21358 3136 21364 3148
rect 21416 3136 21422 3188
rect 22002 3136 22008 3188
rect 22060 3176 22066 3188
rect 22097 3179 22155 3185
rect 22097 3176 22109 3179
rect 22060 3148 22109 3176
rect 22060 3136 22066 3148
rect 22097 3145 22109 3148
rect 22143 3145 22155 3179
rect 24762 3176 24768 3188
rect 24723 3148 24768 3176
rect 22097 3139 22155 3145
rect 24762 3136 24768 3148
rect 24820 3136 24826 3188
rect 16114 3068 16120 3120
rect 16172 3108 16178 3120
rect 17037 3111 17095 3117
rect 17037 3108 17049 3111
rect 16172 3080 17049 3108
rect 16172 3068 16178 3080
rect 17037 3077 17049 3080
rect 17083 3077 17095 3111
rect 17037 3071 17095 3077
rect 12253 3043 12311 3049
rect 12253 3009 12265 3043
rect 12299 3040 12311 3043
rect 16390 3040 16396 3052
rect 12299 3012 12572 3040
rect 16351 3012 16396 3040
rect 12299 3009 12311 3012
rect 12253 3003 12311 3009
rect 12544 2984 12572 3012
rect 16390 3000 16396 3012
rect 16448 3000 16454 3052
rect 18322 3000 18328 3052
rect 18380 3040 18386 3052
rect 18509 3043 18567 3049
rect 18509 3040 18521 3043
rect 18380 3012 18521 3040
rect 18380 3000 18386 3012
rect 18509 3009 18521 3012
rect 18555 3009 18567 3043
rect 18509 3003 18567 3009
rect 18598 3000 18604 3052
rect 18656 3040 18662 3052
rect 18656 3012 18701 3040
rect 18656 3000 18662 3012
rect 19058 3000 19064 3052
rect 19116 3040 19122 3052
rect 19429 3043 19487 3049
rect 19429 3040 19441 3043
rect 19116 3012 19441 3040
rect 19116 3000 19122 3012
rect 19429 3009 19441 3012
rect 19475 3009 19487 3043
rect 19429 3003 19487 3009
rect 20533 3043 20591 3049
rect 20533 3009 20545 3043
rect 20579 3040 20591 3043
rect 21818 3040 21824 3052
rect 20579 3012 21824 3040
rect 20579 3009 20591 3012
rect 20533 3003 20591 3009
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 11793 2975 11851 2981
rect 11793 2972 11805 2975
rect 11480 2944 11805 2972
rect 11480 2932 11486 2944
rect 11793 2941 11805 2944
rect 11839 2941 11851 2975
rect 11793 2935 11851 2941
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12400 2944 12449 2972
rect 12400 2932 12406 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 8754 2904 8760 2916
rect 8220 2876 8760 2904
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 12452 2904 12480 2935
rect 12526 2932 12532 2984
rect 12584 2972 12590 2984
rect 12693 2975 12751 2981
rect 12693 2972 12705 2975
rect 12584 2944 12705 2972
rect 12584 2932 12590 2944
rect 12693 2941 12705 2944
rect 12739 2941 12751 2975
rect 14645 2975 14703 2981
rect 14645 2972 14657 2975
rect 12693 2935 12751 2941
rect 14108 2944 14657 2972
rect 14108 2904 14136 2944
rect 14645 2941 14657 2944
rect 14691 2972 14703 2975
rect 15470 2972 15476 2984
rect 14691 2944 15476 2972
rect 14691 2941 14703 2944
rect 14645 2935 14703 2941
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 16853 2975 16911 2981
rect 16853 2941 16865 2975
rect 16899 2972 16911 2975
rect 16942 2972 16948 2984
rect 16899 2944 16948 2972
rect 16899 2941 16911 2944
rect 16853 2935 16911 2941
rect 16942 2932 16948 2944
rect 17000 2932 17006 2984
rect 20254 2972 20260 2984
rect 20215 2944 20260 2972
rect 20254 2932 20260 2944
rect 20312 2972 20318 2984
rect 20993 2975 21051 2981
rect 20993 2972 21005 2975
rect 20312 2944 21005 2972
rect 20312 2932 20318 2944
rect 20993 2941 21005 2944
rect 21039 2941 21051 2975
rect 20993 2935 21051 2941
rect 21358 2932 21364 2984
rect 21416 2972 21422 2984
rect 21545 2975 21603 2981
rect 21545 2972 21557 2975
rect 21416 2944 21557 2972
rect 21416 2932 21422 2944
rect 21545 2941 21557 2944
rect 21591 2941 21603 2975
rect 21545 2935 21603 2941
rect 24581 2975 24639 2981
rect 24581 2941 24593 2975
rect 24627 2941 24639 2975
rect 24581 2935 24639 2941
rect 12452 2876 14136 2904
rect 14182 2864 14188 2916
rect 14240 2904 14246 2916
rect 14890 2907 14948 2913
rect 14890 2904 14902 2907
rect 14240 2876 14902 2904
rect 14240 2864 14246 2876
rect 14890 2873 14902 2876
rect 14936 2873 14948 2907
rect 24596 2904 24624 2935
rect 25222 2904 25228 2916
rect 24596 2876 25228 2904
rect 14890 2867 14948 2873
rect 25222 2864 25228 2876
rect 25280 2864 25286 2916
rect 7006 2836 7012 2848
rect 6967 2808 7012 2836
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 10229 2839 10287 2845
rect 10229 2836 10241 2839
rect 10192 2808 10241 2836
rect 10192 2796 10198 2808
rect 10229 2805 10241 2808
rect 10275 2836 10287 2839
rect 10781 2839 10839 2845
rect 10781 2836 10793 2839
rect 10275 2808 10793 2836
rect 10275 2805 10287 2808
rect 10229 2799 10287 2805
rect 10781 2805 10793 2808
rect 10827 2805 10839 2839
rect 13814 2836 13820 2848
rect 13775 2808 13820 2836
rect 10781 2799 10839 2805
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 16022 2836 16028 2848
rect 15983 2808 16028 2836
rect 16022 2796 16028 2808
rect 16080 2796 16086 2848
rect 18138 2796 18144 2848
rect 18196 2836 18202 2848
rect 18417 2839 18475 2845
rect 18417 2836 18429 2839
rect 18196 2808 18429 2836
rect 18196 2796 18202 2808
rect 18417 2805 18429 2808
rect 18463 2805 18475 2839
rect 21726 2836 21732 2848
rect 21687 2808 21732 2836
rect 18417 2799 18475 2805
rect 21726 2796 21732 2808
rect 21784 2796 21790 2848
rect 23934 2836 23940 2848
rect 23895 2808 23940 2836
rect 23934 2796 23940 2808
rect 23992 2796 23998 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1673 2635 1731 2641
rect 1673 2601 1685 2635
rect 1719 2632 1731 2635
rect 1946 2632 1952 2644
rect 1719 2604 1952 2632
rect 1719 2601 1731 2604
rect 1673 2595 1731 2601
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 2498 2592 2504 2644
rect 2556 2632 2562 2644
rect 2593 2635 2651 2641
rect 2593 2632 2605 2635
rect 2556 2604 2605 2632
rect 2556 2592 2562 2604
rect 2593 2601 2605 2604
rect 2639 2601 2651 2635
rect 3234 2632 3240 2644
rect 3195 2604 3240 2632
rect 2593 2595 2651 2601
rect 3234 2592 3240 2604
rect 3292 2592 3298 2644
rect 5718 2632 5724 2644
rect 5679 2604 5724 2632
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 5994 2632 6000 2644
rect 5955 2604 6000 2632
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 8849 2635 8907 2641
rect 8849 2601 8861 2635
rect 8895 2632 8907 2635
rect 9030 2632 9036 2644
rect 8895 2604 9036 2632
rect 8895 2601 8907 2604
rect 8849 2595 8907 2601
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 10505 2635 10563 2641
rect 10505 2601 10517 2635
rect 10551 2632 10563 2635
rect 10870 2632 10876 2644
rect 10551 2604 10876 2632
rect 10551 2601 10563 2604
rect 10505 2595 10563 2601
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 11422 2632 11428 2644
rect 11383 2604 11428 2632
rect 11422 2592 11428 2604
rect 11480 2592 11486 2644
rect 12437 2635 12495 2641
rect 12437 2601 12449 2635
rect 12483 2632 12495 2635
rect 14182 2632 14188 2644
rect 12483 2604 12517 2632
rect 14143 2604 14188 2632
rect 12483 2601 12495 2604
rect 12437 2595 12495 2601
rect 4614 2573 4620 2576
rect 3881 2567 3939 2573
rect 3881 2533 3893 2567
rect 3927 2564 3939 2567
rect 4586 2567 4620 2573
rect 4586 2564 4598 2567
rect 3927 2536 4598 2564
rect 3927 2533 3939 2536
rect 3881 2527 3939 2533
rect 4586 2533 4598 2536
rect 4672 2564 4678 2576
rect 7377 2567 7435 2573
rect 4672 2536 4734 2564
rect 4586 2527 4620 2533
rect 4614 2524 4620 2527
rect 4672 2524 4678 2536
rect 7377 2533 7389 2567
rect 7423 2564 7435 2567
rect 7714 2567 7772 2573
rect 7714 2564 7726 2567
rect 7423 2536 7726 2564
rect 7423 2533 7435 2536
rect 7377 2527 7435 2533
rect 7714 2533 7726 2536
rect 7760 2564 7772 2567
rect 8662 2564 8668 2576
rect 7760 2536 8668 2564
rect 7760 2533 7772 2536
rect 7714 2527 7772 2533
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 9674 2524 9680 2576
rect 9732 2564 9738 2576
rect 10781 2567 10839 2573
rect 10781 2564 10793 2567
rect 9732 2536 10793 2564
rect 9732 2524 9738 2536
rect 10781 2533 10793 2536
rect 10827 2564 10839 2567
rect 11333 2567 11391 2573
rect 11333 2564 11345 2567
rect 10827 2536 11345 2564
rect 10827 2533 10839 2536
rect 10781 2527 10839 2533
rect 11333 2533 11345 2536
rect 11379 2533 11391 2567
rect 11333 2527 11391 2533
rect 12069 2567 12127 2573
rect 12069 2533 12081 2567
rect 12115 2564 12127 2567
rect 12452 2564 12480 2595
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 15289 2635 15347 2641
rect 15289 2601 15301 2635
rect 15335 2632 15347 2635
rect 15838 2632 15844 2644
rect 15335 2604 15844 2632
rect 15335 2601 15347 2604
rect 15289 2595 15347 2601
rect 15838 2592 15844 2604
rect 15896 2592 15902 2644
rect 16577 2635 16635 2641
rect 16577 2601 16589 2635
rect 16623 2632 16635 2635
rect 16666 2632 16672 2644
rect 16623 2604 16672 2632
rect 16623 2601 16635 2604
rect 16577 2595 16635 2601
rect 16666 2592 16672 2604
rect 16724 2592 16730 2644
rect 17681 2635 17739 2641
rect 17681 2601 17693 2635
rect 17727 2632 17739 2635
rect 17770 2632 17776 2644
rect 17727 2604 17776 2632
rect 17727 2601 17739 2604
rect 17681 2595 17739 2601
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 18138 2632 18144 2644
rect 18099 2604 18144 2632
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 20898 2632 20904 2644
rect 20859 2604 20904 2632
rect 20898 2592 20904 2604
rect 20956 2592 20962 2644
rect 24762 2632 24768 2644
rect 24723 2604 24768 2632
rect 24762 2592 24768 2604
rect 24820 2592 24826 2644
rect 13072 2567 13130 2573
rect 13072 2564 13084 2567
rect 12115 2536 13084 2564
rect 12115 2533 12127 2536
rect 12069 2527 12127 2533
rect 13072 2533 13084 2536
rect 13118 2564 13130 2567
rect 13814 2564 13820 2576
rect 13118 2536 13820 2564
rect 13118 2533 13130 2536
rect 13072 2527 13130 2533
rect 1394 2456 1400 2508
rect 1452 2496 1458 2508
rect 2501 2499 2559 2505
rect 2501 2496 2513 2499
rect 1452 2468 2513 2496
rect 1452 2456 1458 2468
rect 2501 2465 2513 2468
rect 2547 2496 2559 2499
rect 2958 2496 2964 2508
rect 2547 2468 2964 2496
rect 2547 2465 2559 2468
rect 2501 2459 2559 2465
rect 2958 2456 2964 2468
rect 3016 2456 3022 2508
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2496 4399 2499
rect 4430 2496 4436 2508
rect 4387 2468 4436 2496
rect 4387 2465 4399 2468
rect 4341 2459 4399 2465
rect 4430 2456 4436 2468
rect 4488 2456 4494 2508
rect 7466 2496 7472 2508
rect 7427 2468 7472 2496
rect 7466 2456 7472 2468
rect 7524 2456 7530 2508
rect 9217 2499 9275 2505
rect 9217 2465 9229 2499
rect 9263 2496 9275 2499
rect 9861 2499 9919 2505
rect 9861 2496 9873 2499
rect 9263 2468 9873 2496
rect 9263 2465 9275 2468
rect 9217 2459 9275 2465
rect 9861 2465 9873 2468
rect 9907 2496 9919 2499
rect 9950 2496 9956 2508
rect 9907 2468 9956 2496
rect 9907 2465 9919 2468
rect 9861 2459 9919 2465
rect 9950 2456 9956 2468
rect 10008 2456 10014 2508
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2428 2835 2431
rect 3234 2428 3240 2440
rect 2823 2400 3240 2428
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 6362 2428 6368 2440
rect 6323 2400 6368 2428
rect 6362 2388 6368 2400
rect 6420 2388 6426 2440
rect 9582 2428 9588 2440
rect 9543 2400 9588 2428
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 11609 2431 11667 2437
rect 11609 2397 11621 2431
rect 11655 2428 11667 2431
rect 12084 2428 12112 2527
rect 13814 2524 13820 2536
rect 13872 2524 13878 2576
rect 15933 2567 15991 2573
rect 15933 2564 15945 2567
rect 14476 2536 15945 2564
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 12805 2499 12863 2505
rect 12805 2496 12817 2499
rect 12492 2468 12817 2496
rect 12492 2456 12498 2468
rect 12805 2465 12817 2468
rect 12851 2465 12863 2499
rect 12805 2459 12863 2465
rect 13630 2456 13636 2508
rect 13688 2496 13694 2508
rect 14476 2505 14504 2536
rect 15933 2533 15945 2536
rect 15979 2533 15991 2567
rect 19889 2567 19947 2573
rect 19889 2564 19901 2567
rect 15933 2527 15991 2533
rect 17052 2536 19901 2564
rect 17052 2505 17080 2536
rect 19889 2533 19901 2536
rect 19935 2533 19947 2567
rect 19889 2527 19947 2533
rect 20714 2524 20720 2576
rect 20772 2564 20778 2576
rect 21453 2567 21511 2573
rect 21453 2564 21465 2567
rect 20772 2536 21465 2564
rect 20772 2524 20778 2536
rect 21453 2533 21465 2536
rect 21499 2533 21511 2567
rect 21453 2527 21511 2533
rect 14461 2499 14519 2505
rect 14461 2496 14473 2499
rect 13688 2468 14473 2496
rect 13688 2456 13694 2468
rect 14461 2465 14473 2468
rect 14507 2465 14519 2499
rect 14461 2459 14519 2465
rect 16945 2499 17003 2505
rect 16945 2465 16957 2499
rect 16991 2496 17003 2499
rect 17037 2499 17095 2505
rect 17037 2496 17049 2499
rect 16991 2468 17049 2496
rect 16991 2465 17003 2468
rect 16945 2459 17003 2465
rect 17037 2465 17049 2468
rect 17083 2465 17095 2499
rect 18322 2496 18328 2508
rect 18283 2468 18328 2496
rect 17037 2459 17095 2465
rect 18322 2456 18328 2468
rect 18380 2496 18386 2508
rect 19061 2499 19119 2505
rect 19061 2496 19073 2499
rect 18380 2468 19073 2496
rect 18380 2456 18386 2468
rect 19061 2465 19073 2468
rect 19107 2465 19119 2499
rect 19610 2496 19616 2508
rect 19571 2468 19616 2496
rect 19061 2459 19119 2465
rect 19610 2456 19616 2468
rect 19668 2496 19674 2508
rect 20349 2499 20407 2505
rect 20349 2496 20361 2499
rect 19668 2468 20361 2496
rect 19668 2456 19674 2468
rect 20349 2465 20361 2468
rect 20395 2465 20407 2499
rect 21174 2496 21180 2508
rect 21135 2468 21180 2496
rect 20349 2459 20407 2465
rect 21174 2456 21180 2468
rect 21232 2496 21238 2508
rect 21913 2499 21971 2505
rect 21913 2496 21925 2499
rect 21232 2468 21925 2496
rect 21232 2456 21238 2468
rect 21913 2465 21925 2468
rect 21959 2465 21971 2499
rect 22462 2496 22468 2508
rect 22423 2468 22468 2496
rect 21913 2459 21971 2465
rect 22462 2456 22468 2468
rect 22520 2496 22526 2508
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22520 2468 23029 2496
rect 22520 2456 22526 2468
rect 23017 2465 23029 2468
rect 23063 2465 23075 2499
rect 23017 2459 23075 2465
rect 11655 2400 12112 2428
rect 14921 2431 14979 2437
rect 11655 2397 11667 2400
rect 11609 2391 11667 2397
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 15286 2428 15292 2440
rect 14967 2400 15292 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 15286 2388 15292 2400
rect 15344 2428 15350 2440
rect 16022 2428 16028 2440
rect 15344 2400 16028 2428
rect 15344 2388 15350 2400
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 18506 2428 18512 2440
rect 18467 2400 18512 2428
rect 18506 2388 18512 2400
rect 18564 2388 18570 2440
rect 2130 2360 2136 2372
rect 2091 2332 2136 2360
rect 2130 2320 2136 2332
rect 2188 2320 2194 2372
rect 10045 2363 10103 2369
rect 10045 2329 10057 2363
rect 10091 2360 10103 2363
rect 10686 2360 10692 2372
rect 10091 2332 10692 2360
rect 10091 2329 10103 2332
rect 10045 2323 10103 2329
rect 10686 2320 10692 2332
rect 10744 2320 10750 2372
rect 15470 2360 15476 2372
rect 15431 2332 15476 2360
rect 15470 2320 15476 2332
rect 15528 2320 15534 2372
rect 15562 2320 15568 2372
rect 15620 2360 15626 2372
rect 17221 2363 17279 2369
rect 17221 2360 17233 2363
rect 15620 2332 17233 2360
rect 15620 2320 15626 2332
rect 17221 2329 17233 2332
rect 17267 2329 17279 2363
rect 17221 2323 17279 2329
rect 2038 2292 2044 2304
rect 1951 2264 2044 2292
rect 2038 2252 2044 2264
rect 2096 2292 2102 2304
rect 9398 2292 9404 2304
rect 2096 2264 9404 2292
rect 2096 2252 2102 2264
rect 9398 2252 9404 2264
rect 9456 2252 9462 2304
rect 10962 2292 10968 2304
rect 10923 2264 10968 2292
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 22646 2292 22652 2304
rect 22607 2264 22652 2292
rect 22646 2252 22652 2264
rect 22704 2252 22710 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 5626 1980 5632 2032
rect 5684 2020 5690 2032
rect 6270 2020 6276 2032
rect 5684 1992 6276 2020
rect 5684 1980 5690 1992
rect 6270 1980 6276 1992
rect 6328 1980 6334 2032
rect 14274 1980 14280 2032
rect 14332 2020 14338 2032
rect 14918 2020 14924 2032
rect 14332 1992 14924 2020
rect 14332 1980 14338 1992
rect 14918 1980 14924 1992
rect 14976 1980 14982 2032
rect 23474 1980 23480 2032
rect 23532 2020 23538 2032
rect 24302 2020 24308 2032
rect 23532 1992 24308 2020
rect 23532 1980 23538 1992
rect 24302 1980 24308 1992
rect 24360 1980 24366 2032
rect 9858 1368 9864 1420
rect 9916 1408 9922 1420
rect 10594 1408 10600 1420
rect 9916 1380 10600 1408
rect 9916 1368 9922 1380
rect 10594 1368 10600 1380
rect 10652 1368 10658 1420
rect 11606 552 11612 604
rect 11664 592 11670 604
rect 11698 592 11704 604
rect 11664 564 11704 592
rect 11664 552 11670 564
rect 11698 552 11704 564
rect 11756 552 11762 604
rect 23566 552 23572 604
rect 23624 592 23630 604
rect 23750 592 23756 604
rect 23624 564 23756 592
rect 23624 552 23630 564
rect 23750 552 23756 564
rect 23808 552 23814 604
rect 24946 552 24952 604
rect 25004 592 25010 604
rect 25406 592 25412 604
rect 25004 564 25412 592
rect 25004 552 25010 564
rect 25406 552 25412 564
rect 25464 552 25470 604
<< via1 >>
rect 4068 26528 4120 26580
rect 5540 26528 5592 26580
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1584 24395 1636 24404
rect 1584 24361 1593 24395
rect 1593 24361 1627 24395
rect 1627 24361 1636 24395
rect 1584 24352 1636 24361
rect 1400 24259 1452 24268
rect 1400 24225 1409 24259
rect 1409 24225 1443 24259
rect 1443 24225 1452 24259
rect 1400 24216 1452 24225
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1400 23808 1452 23860
rect 1860 23808 1912 23860
rect 2688 23851 2740 23860
rect 2688 23817 2697 23851
rect 2697 23817 2731 23851
rect 2731 23817 2740 23851
rect 2688 23808 2740 23817
rect 3792 23851 3844 23860
rect 3792 23817 3801 23851
rect 3801 23817 3835 23851
rect 3835 23817 3844 23851
rect 3792 23808 3844 23817
rect 20996 23808 21048 23860
rect 1952 23604 2004 23656
rect 1584 23511 1636 23520
rect 1584 23477 1593 23511
rect 1593 23477 1627 23511
rect 1627 23477 1636 23511
rect 1584 23468 1636 23477
rect 2596 23468 2648 23520
rect 4436 23468 4488 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 8300 23307 8352 23316
rect 8300 23273 8309 23307
rect 8309 23273 8343 23307
rect 8343 23273 8352 23307
rect 8300 23264 8352 23273
rect 1952 23239 2004 23248
rect 1952 23205 1961 23239
rect 1961 23205 1995 23239
rect 1995 23205 2004 23239
rect 1952 23196 2004 23205
rect 2872 23128 2924 23180
rect 8116 23171 8168 23180
rect 8116 23137 8125 23171
rect 8125 23137 8159 23171
rect 8159 23137 8168 23171
rect 8116 23128 8168 23137
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 4160 22720 4212 22772
rect 7472 22763 7524 22772
rect 7472 22729 7481 22763
rect 7481 22729 7515 22763
rect 7515 22729 7524 22763
rect 7472 22720 7524 22729
rect 8116 22720 8168 22772
rect 1860 22627 1912 22636
rect 1860 22593 1869 22627
rect 1869 22593 1903 22627
rect 1903 22593 1912 22627
rect 1860 22584 1912 22593
rect 2780 22516 2832 22568
rect 2504 22423 2556 22432
rect 2504 22389 2513 22423
rect 2513 22389 2547 22423
rect 2547 22389 2556 22423
rect 2504 22380 2556 22389
rect 2872 22423 2924 22432
rect 2872 22389 2881 22423
rect 2881 22389 2915 22423
rect 2915 22389 2924 22423
rect 2872 22380 2924 22389
rect 3148 22423 3200 22432
rect 3148 22389 3157 22423
rect 3157 22389 3191 22423
rect 3191 22389 3200 22423
rect 3148 22380 3200 22389
rect 4712 22423 4764 22432
rect 4712 22389 4721 22423
rect 4721 22389 4755 22423
rect 4755 22389 4764 22423
rect 4712 22380 4764 22389
rect 8116 22380 8168 22432
rect 9588 22423 9640 22432
rect 9588 22389 9597 22423
rect 9597 22389 9631 22423
rect 9631 22389 9640 22423
rect 9588 22380 9640 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 2044 22040 2096 22092
rect 2504 22083 2556 22092
rect 2504 22049 2513 22083
rect 2513 22049 2547 22083
rect 2547 22049 2556 22083
rect 2504 22040 2556 22049
rect 4068 22083 4120 22092
rect 4068 22049 4077 22083
rect 4077 22049 4111 22083
rect 4111 22049 4120 22083
rect 4068 22040 4120 22049
rect 6000 22040 6052 22092
rect 7840 22040 7892 22092
rect 2136 21972 2188 22024
rect 8300 22015 8352 22024
rect 8300 21981 8309 22015
rect 8309 21981 8343 22015
rect 8343 21981 8352 22015
rect 8300 21972 8352 21981
rect 2228 21904 2280 21956
rect 4252 21947 4304 21956
rect 4252 21913 4261 21947
rect 4261 21913 4295 21947
rect 4295 21913 4304 21947
rect 4252 21904 4304 21913
rect 5540 21904 5592 21956
rect 2044 21836 2096 21888
rect 2872 21836 2924 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 4068 21632 4120 21684
rect 4528 21632 4580 21684
rect 5264 21675 5316 21684
rect 5264 21641 5273 21675
rect 5273 21641 5307 21675
rect 5307 21641 5316 21675
rect 5264 21632 5316 21641
rect 6000 21675 6052 21684
rect 6000 21641 6009 21675
rect 6009 21641 6043 21675
rect 6043 21641 6052 21675
rect 6000 21632 6052 21641
rect 2688 21496 2740 21548
rect 8116 21539 8168 21548
rect 8116 21505 8125 21539
rect 8125 21505 8159 21539
rect 8159 21505 8168 21539
rect 8116 21496 8168 21505
rect 2136 21428 2188 21480
rect 2780 21428 2832 21480
rect 3976 21471 4028 21480
rect 3976 21437 3985 21471
rect 3985 21437 4019 21471
rect 4019 21437 4028 21471
rect 3976 21428 4028 21437
rect 5080 21471 5132 21480
rect 5080 21437 5089 21471
rect 5089 21437 5123 21471
rect 5123 21437 5132 21471
rect 5080 21428 5132 21437
rect 7932 21471 7984 21480
rect 7932 21437 7941 21471
rect 7941 21437 7975 21471
rect 7975 21437 7984 21471
rect 7932 21428 7984 21437
rect 2504 21335 2556 21344
rect 2504 21301 2513 21335
rect 2513 21301 2547 21335
rect 2547 21301 2556 21335
rect 2504 21292 2556 21301
rect 3056 21335 3108 21344
rect 3056 21301 3065 21335
rect 3065 21301 3099 21335
rect 3099 21301 3108 21335
rect 3056 21292 3108 21301
rect 4160 21335 4212 21344
rect 4160 21301 4169 21335
rect 4169 21301 4203 21335
rect 4203 21301 4212 21335
rect 4160 21292 4212 21301
rect 7840 21335 7892 21344
rect 7840 21301 7849 21335
rect 7849 21301 7883 21335
rect 7883 21301 7892 21335
rect 7840 21292 7892 21301
rect 10048 21292 10100 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 9680 21131 9732 21140
rect 9680 21097 9689 21131
rect 9689 21097 9723 21131
rect 9723 21097 9732 21131
rect 9680 21088 9732 21097
rect 10048 21131 10100 21140
rect 10048 21097 10057 21131
rect 10057 21097 10091 21131
rect 10091 21097 10100 21131
rect 10048 21088 10100 21097
rect 1952 21063 2004 21072
rect 1952 21029 1961 21063
rect 1961 21029 1995 21063
rect 1995 21029 2004 21063
rect 1952 21020 2004 21029
rect 4436 21063 4488 21072
rect 4436 21029 4445 21063
rect 4445 21029 4479 21063
rect 4479 21029 4488 21063
rect 4436 21020 4488 21029
rect 6000 21020 6052 21072
rect 1676 20995 1728 21004
rect 1676 20961 1685 20995
rect 1685 20961 1719 20995
rect 1719 20961 1728 20995
rect 1676 20952 1728 20961
rect 4252 20952 4304 21004
rect 6092 20995 6144 21004
rect 6092 20961 6101 20995
rect 6101 20961 6135 20995
rect 6135 20961 6144 20995
rect 6092 20952 6144 20961
rect 7196 20884 7248 20936
rect 10140 20927 10192 20936
rect 10140 20893 10149 20927
rect 10149 20893 10183 20927
rect 10183 20893 10192 20927
rect 10140 20884 10192 20893
rect 10692 20884 10744 20936
rect 6920 20791 6972 20800
rect 6920 20757 6929 20791
rect 6929 20757 6963 20791
rect 6963 20757 6972 20791
rect 6920 20748 6972 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 10048 20587 10100 20596
rect 10048 20553 10057 20587
rect 10057 20553 10091 20587
rect 10091 20553 10100 20587
rect 10048 20544 10100 20553
rect 10140 20544 10192 20596
rect 10692 20476 10744 20528
rect 1952 20451 2004 20460
rect 1952 20417 1961 20451
rect 1961 20417 1995 20451
rect 1995 20417 2004 20451
rect 1952 20408 2004 20417
rect 2596 20408 2648 20460
rect 4528 20451 4580 20460
rect 4528 20417 4537 20451
rect 4537 20417 4571 20451
rect 4571 20417 4580 20451
rect 4528 20408 4580 20417
rect 1768 20340 1820 20392
rect 2320 20272 2372 20324
rect 5540 20383 5592 20392
rect 5540 20349 5549 20383
rect 5549 20349 5583 20383
rect 5583 20349 5592 20383
rect 5540 20340 5592 20349
rect 6920 20340 6972 20392
rect 7380 20340 7432 20392
rect 5448 20272 5500 20324
rect 2412 20204 2464 20256
rect 2596 20204 2648 20256
rect 3608 20204 3660 20256
rect 4160 20247 4212 20256
rect 4160 20213 4169 20247
rect 4169 20213 4203 20247
rect 4203 20213 4212 20247
rect 4160 20204 4212 20213
rect 5080 20247 5132 20256
rect 5080 20213 5089 20247
rect 5089 20213 5123 20247
rect 5123 20213 5132 20247
rect 5080 20204 5132 20213
rect 5356 20247 5408 20256
rect 5356 20213 5365 20247
rect 5365 20213 5399 20247
rect 5399 20213 5408 20247
rect 5356 20204 5408 20213
rect 5724 20247 5776 20256
rect 5724 20213 5733 20247
rect 5733 20213 5767 20247
rect 5767 20213 5776 20247
rect 5724 20204 5776 20213
rect 8208 20247 8260 20256
rect 8208 20213 8217 20247
rect 8217 20213 8251 20247
rect 8251 20213 8260 20247
rect 8208 20204 8260 20213
rect 9312 20204 9364 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 2688 20000 2740 20052
rect 4160 20000 4212 20052
rect 6092 20000 6144 20052
rect 10692 20000 10744 20052
rect 3976 19932 4028 19984
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 2688 19907 2740 19916
rect 2688 19873 2697 19907
rect 2697 19873 2731 19907
rect 2731 19873 2740 19907
rect 2688 19864 2740 19873
rect 5080 19932 5132 19984
rect 5356 19932 5408 19984
rect 9864 19932 9916 19984
rect 4712 19864 4764 19916
rect 8208 19864 8260 19916
rect 5356 19839 5408 19848
rect 5356 19805 5365 19839
rect 5365 19805 5399 19839
rect 5399 19805 5408 19839
rect 5356 19796 5408 19805
rect 5448 19839 5500 19848
rect 5448 19805 5457 19839
rect 5457 19805 5491 19839
rect 5491 19805 5500 19839
rect 7380 19839 7432 19848
rect 5448 19796 5500 19805
rect 7380 19805 7389 19839
rect 7389 19805 7423 19839
rect 7423 19805 7432 19839
rect 7380 19796 7432 19805
rect 1676 19660 1728 19712
rect 2136 19703 2188 19712
rect 2136 19669 2145 19703
rect 2145 19669 2179 19703
rect 2179 19669 2188 19703
rect 2136 19660 2188 19669
rect 2412 19660 2464 19712
rect 3516 19703 3568 19712
rect 3516 19669 3525 19703
rect 3525 19669 3559 19703
rect 3559 19669 3568 19703
rect 3516 19660 3568 19669
rect 4160 19660 4212 19712
rect 6000 19703 6052 19712
rect 6000 19669 6009 19703
rect 6009 19669 6043 19703
rect 6043 19669 6052 19703
rect 6000 19660 6052 19669
rect 6920 19703 6972 19712
rect 6920 19669 6929 19703
rect 6929 19669 6963 19703
rect 6963 19669 6972 19703
rect 6920 19660 6972 19669
rect 7288 19703 7340 19712
rect 7288 19669 7297 19703
rect 7297 19669 7331 19703
rect 7331 19669 7340 19703
rect 7288 19660 7340 19669
rect 8668 19660 8720 19712
rect 9036 19703 9088 19712
rect 9036 19669 9045 19703
rect 9045 19669 9079 19703
rect 9079 19669 9088 19703
rect 9036 19660 9088 19669
rect 9312 19660 9364 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1400 19456 1452 19508
rect 4712 19499 4764 19508
rect 4712 19465 4721 19499
rect 4721 19465 4755 19499
rect 4755 19465 4764 19499
rect 4712 19456 4764 19465
rect 5172 19499 5224 19508
rect 5172 19465 5181 19499
rect 5181 19465 5215 19499
rect 5215 19465 5224 19499
rect 5172 19456 5224 19465
rect 6092 19456 6144 19508
rect 10140 19456 10192 19508
rect 1492 19320 1544 19372
rect 2688 19363 2740 19372
rect 2688 19329 2697 19363
rect 2697 19329 2731 19363
rect 2731 19329 2740 19363
rect 2688 19320 2740 19329
rect 6000 19388 6052 19440
rect 6736 19388 6788 19440
rect 6920 19388 6972 19440
rect 6828 19320 6880 19372
rect 7288 19363 7340 19372
rect 7288 19329 7297 19363
rect 7297 19329 7331 19363
rect 7331 19329 7340 19363
rect 7288 19320 7340 19329
rect 1584 19295 1636 19304
rect 1584 19261 1593 19295
rect 1593 19261 1627 19295
rect 1627 19261 1636 19295
rect 1584 19252 1636 19261
rect 2044 19252 2096 19304
rect 2872 19295 2924 19304
rect 2872 19261 2881 19295
rect 2881 19261 2915 19295
rect 2915 19261 2924 19295
rect 2872 19252 2924 19261
rect 7196 19295 7248 19304
rect 7196 19261 7205 19295
rect 7205 19261 7239 19295
rect 7239 19261 7248 19295
rect 7196 19252 7248 19261
rect 9864 19320 9916 19372
rect 8668 19295 8720 19304
rect 8668 19261 8691 19295
rect 8691 19261 8720 19295
rect 2504 19184 2556 19236
rect 5356 19184 5408 19236
rect 8668 19252 8720 19261
rect 10968 19252 11020 19304
rect 9312 19184 9364 19236
rect 2136 19116 2188 19168
rect 2596 19116 2648 19168
rect 5632 19116 5684 19168
rect 8208 19116 8260 19168
rect 9496 19116 9548 19168
rect 9864 19116 9916 19168
rect 10048 19116 10100 19168
rect 12808 19116 12860 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 5448 18912 5500 18964
rect 7288 18912 7340 18964
rect 9496 18955 9548 18964
rect 9496 18921 9505 18955
rect 9505 18921 9539 18955
rect 9539 18921 9548 18955
rect 9496 18912 9548 18921
rect 9772 18912 9824 18964
rect 2044 18776 2096 18828
rect 2320 18819 2372 18828
rect 2320 18785 2329 18819
rect 2329 18785 2363 18819
rect 2363 18785 2372 18819
rect 2320 18776 2372 18785
rect 4068 18819 4120 18828
rect 4068 18785 4077 18819
rect 4077 18785 4111 18819
rect 4111 18785 4120 18819
rect 4068 18776 4120 18785
rect 5540 18819 5592 18828
rect 5540 18785 5574 18819
rect 5574 18785 5592 18819
rect 5540 18776 5592 18785
rect 7380 18776 7432 18828
rect 8392 18776 8444 18828
rect 9220 18776 9272 18828
rect 2412 18751 2464 18760
rect 2412 18717 2421 18751
rect 2421 18717 2455 18751
rect 2455 18717 2464 18751
rect 2412 18708 2464 18717
rect 2504 18751 2556 18760
rect 2504 18717 2513 18751
rect 2513 18717 2547 18751
rect 2547 18717 2556 18751
rect 2504 18708 2556 18717
rect 5172 18708 5224 18760
rect 8208 18708 8260 18760
rect 10140 18751 10192 18760
rect 10140 18717 10149 18751
rect 10149 18717 10183 18751
rect 10183 18717 10192 18751
rect 10140 18708 10192 18717
rect 10324 18751 10376 18760
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 10968 18708 11020 18760
rect 1952 18615 2004 18624
rect 1952 18581 1961 18615
rect 1961 18581 1995 18615
rect 1995 18581 2004 18615
rect 1952 18572 2004 18581
rect 2964 18615 3016 18624
rect 2964 18581 2973 18615
rect 2973 18581 3007 18615
rect 3007 18581 3016 18615
rect 2964 18572 3016 18581
rect 3700 18615 3752 18624
rect 3700 18581 3709 18615
rect 3709 18581 3743 18615
rect 3743 18581 3752 18615
rect 3700 18572 3752 18581
rect 4252 18615 4304 18624
rect 4252 18581 4261 18615
rect 4261 18581 4295 18615
rect 4295 18581 4304 18615
rect 4252 18572 4304 18581
rect 7380 18572 7432 18624
rect 8484 18615 8536 18624
rect 8484 18581 8493 18615
rect 8493 18581 8527 18615
rect 8527 18581 8536 18615
rect 8484 18572 8536 18581
rect 9036 18572 9088 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 3608 18411 3660 18420
rect 3608 18377 3617 18411
rect 3617 18377 3651 18411
rect 3651 18377 3660 18411
rect 3608 18368 3660 18377
rect 5356 18368 5408 18420
rect 6736 18368 6788 18420
rect 9220 18411 9272 18420
rect 9220 18377 9229 18411
rect 9229 18377 9263 18411
rect 9263 18377 9272 18411
rect 9220 18368 9272 18377
rect 10232 18368 10284 18420
rect 10692 18343 10744 18352
rect 10692 18309 10701 18343
rect 10701 18309 10735 18343
rect 10735 18309 10744 18343
rect 10692 18300 10744 18309
rect 2504 18232 2556 18284
rect 2136 18028 2188 18080
rect 2320 18071 2372 18080
rect 2320 18037 2329 18071
rect 2329 18037 2363 18071
rect 2363 18037 2372 18071
rect 2320 18028 2372 18037
rect 2504 18028 2556 18080
rect 3700 18232 3752 18284
rect 5540 18232 5592 18284
rect 5816 18275 5868 18284
rect 5816 18241 5825 18275
rect 5825 18241 5859 18275
rect 5859 18241 5868 18275
rect 6276 18275 6328 18284
rect 5816 18232 5868 18241
rect 6276 18241 6285 18275
rect 6285 18241 6319 18275
rect 6319 18241 6328 18275
rect 6276 18232 6328 18241
rect 7748 18275 7800 18284
rect 7748 18241 7757 18275
rect 7757 18241 7791 18275
rect 7791 18241 7800 18275
rect 7748 18232 7800 18241
rect 8392 18164 8444 18216
rect 9312 18207 9364 18216
rect 9312 18173 9321 18207
rect 9321 18173 9355 18207
rect 9355 18173 9364 18207
rect 9312 18164 9364 18173
rect 9404 18164 9456 18216
rect 10324 18164 10376 18216
rect 2780 18096 2832 18148
rect 3332 18028 3384 18080
rect 4068 18071 4120 18080
rect 4068 18037 4077 18071
rect 4077 18037 4111 18071
rect 4111 18037 4120 18071
rect 4068 18028 4120 18037
rect 4620 18071 4672 18080
rect 4620 18037 4629 18071
rect 4629 18037 4663 18071
rect 4663 18037 4672 18071
rect 7380 18096 7432 18148
rect 4620 18028 4672 18037
rect 6000 18028 6052 18080
rect 7656 18071 7708 18080
rect 7656 18037 7665 18071
rect 7665 18037 7699 18071
rect 7699 18037 7708 18071
rect 7656 18028 7708 18037
rect 12072 18028 12124 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2688 17824 2740 17876
rect 5816 17867 5868 17876
rect 5816 17833 5825 17867
rect 5825 17833 5859 17867
rect 5859 17833 5868 17867
rect 5816 17824 5868 17833
rect 6092 17824 6144 17876
rect 8300 17867 8352 17876
rect 8300 17833 8309 17867
rect 8309 17833 8343 17867
rect 8343 17833 8352 17867
rect 8300 17824 8352 17833
rect 9220 17824 9272 17876
rect 9404 17867 9456 17876
rect 9404 17833 9413 17867
rect 9413 17833 9447 17867
rect 9447 17833 9456 17867
rect 9404 17824 9456 17833
rect 11060 17824 11112 17876
rect 4068 17756 4120 17808
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 2780 17688 2832 17697
rect 6368 17688 6420 17740
rect 9864 17688 9916 17740
rect 2872 17663 2924 17672
rect 2872 17629 2881 17663
rect 2881 17629 2915 17663
rect 2915 17629 2924 17663
rect 2872 17620 2924 17629
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 3792 17663 3844 17672
rect 2964 17620 3016 17629
rect 3792 17629 3801 17663
rect 3801 17629 3835 17663
rect 3835 17629 3844 17663
rect 3792 17620 3844 17629
rect 3976 17620 4028 17672
rect 1492 17552 1544 17604
rect 9772 17663 9824 17672
rect 9772 17629 9781 17663
rect 9781 17629 9815 17663
rect 9815 17629 9824 17663
rect 9772 17620 9824 17629
rect 7748 17552 7800 17604
rect 1400 17484 1452 17536
rect 2320 17484 2372 17536
rect 5448 17527 5500 17536
rect 5448 17493 5457 17527
rect 5457 17493 5491 17527
rect 5491 17493 5500 17527
rect 5448 17484 5500 17493
rect 6184 17527 6236 17536
rect 6184 17493 6193 17527
rect 6193 17493 6227 17527
rect 6227 17493 6236 17527
rect 6184 17484 6236 17493
rect 7196 17484 7248 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 4068 17280 4120 17332
rect 9956 17280 10008 17332
rect 3792 17212 3844 17264
rect 8116 17212 8168 17264
rect 9312 17255 9364 17264
rect 9312 17221 9321 17255
rect 9321 17221 9355 17255
rect 9355 17221 9364 17255
rect 9312 17212 9364 17221
rect 9772 17212 9824 17264
rect 5448 17144 5500 17196
rect 6368 17187 6420 17196
rect 6368 17153 6377 17187
rect 6377 17153 6411 17187
rect 6411 17153 6420 17187
rect 6368 17144 6420 17153
rect 10692 17144 10744 17196
rect 11244 17187 11296 17196
rect 11244 17153 11253 17187
rect 11253 17153 11287 17187
rect 11287 17153 11296 17187
rect 11244 17144 11296 17153
rect 1584 17076 1636 17128
rect 2504 17076 2556 17128
rect 3976 17076 4028 17128
rect 5816 17076 5868 17128
rect 6184 17076 6236 17128
rect 8208 17076 8260 17128
rect 9312 17076 9364 17128
rect 9864 17076 9916 17128
rect 11336 17076 11388 17128
rect 3056 17051 3108 17060
rect 3056 17017 3090 17051
rect 3090 17017 3108 17051
rect 3056 17008 3108 17017
rect 7196 17008 7248 17060
rect 10784 17008 10836 17060
rect 2780 16940 2832 16992
rect 4068 16940 4120 16992
rect 4620 16940 4672 16992
rect 6000 16940 6052 16992
rect 6920 16940 6972 16992
rect 10140 16983 10192 16992
rect 10140 16949 10149 16983
rect 10149 16949 10183 16983
rect 10183 16949 10192 16983
rect 10140 16940 10192 16949
rect 10692 16983 10744 16992
rect 10692 16949 10701 16983
rect 10701 16949 10735 16983
rect 10735 16949 10744 16983
rect 10692 16940 10744 16949
rect 12072 16940 12124 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1952 16736 2004 16788
rect 2688 16736 2740 16788
rect 2872 16736 2924 16788
rect 7196 16779 7248 16788
rect 7196 16745 7205 16779
rect 7205 16745 7239 16779
rect 7239 16745 7248 16779
rect 7196 16736 7248 16745
rect 8024 16779 8076 16788
rect 8024 16745 8033 16779
rect 8033 16745 8067 16779
rect 8067 16745 8076 16779
rect 8024 16736 8076 16745
rect 10140 16736 10192 16788
rect 11336 16779 11388 16788
rect 11336 16745 11345 16779
rect 11345 16745 11379 16779
rect 11379 16745 11388 16779
rect 11336 16736 11388 16745
rect 2964 16668 3016 16720
rect 3056 16711 3108 16720
rect 3056 16677 3065 16711
rect 3065 16677 3099 16711
rect 3099 16677 3108 16711
rect 3056 16668 3108 16677
rect 4160 16668 4212 16720
rect 6092 16711 6144 16720
rect 2136 16600 2188 16652
rect 3148 16600 3200 16652
rect 4436 16643 4488 16652
rect 4436 16609 4445 16643
rect 4445 16609 4479 16643
rect 4479 16609 4488 16643
rect 4436 16600 4488 16609
rect 6092 16677 6126 16711
rect 6126 16677 6144 16711
rect 6092 16668 6144 16677
rect 6920 16668 6972 16720
rect 7472 16711 7524 16720
rect 7472 16677 7481 16711
rect 7481 16677 7515 16711
rect 7515 16677 7524 16711
rect 7472 16668 7524 16677
rect 8208 16668 8260 16720
rect 5816 16643 5868 16652
rect 5816 16609 5825 16643
rect 5825 16609 5859 16643
rect 5859 16609 5868 16643
rect 5816 16600 5868 16609
rect 8024 16600 8076 16652
rect 2228 16575 2280 16584
rect 2228 16541 2237 16575
rect 2237 16541 2271 16575
rect 2271 16541 2280 16575
rect 2228 16532 2280 16541
rect 4528 16575 4580 16584
rect 4528 16541 4537 16575
rect 4537 16541 4571 16575
rect 4571 16541 4580 16575
rect 4528 16532 4580 16541
rect 3976 16464 4028 16516
rect 4160 16464 4212 16516
rect 5540 16532 5592 16584
rect 8668 16575 8720 16584
rect 5356 16464 5408 16516
rect 8392 16464 8444 16516
rect 8668 16541 8677 16575
rect 8677 16541 8711 16575
rect 8711 16541 8720 16575
rect 9864 16600 9916 16652
rect 10048 16600 10100 16652
rect 10692 16600 10744 16652
rect 8668 16532 8720 16541
rect 9772 16532 9824 16584
rect 9956 16575 10008 16584
rect 9956 16541 9965 16575
rect 9965 16541 9999 16575
rect 9999 16541 10008 16575
rect 9956 16532 10008 16541
rect 1492 16396 1544 16448
rect 5448 16439 5500 16448
rect 5448 16405 5457 16439
rect 5457 16405 5491 16439
rect 5491 16405 5500 16439
rect 5448 16396 5500 16405
rect 9220 16396 9272 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2228 16235 2280 16244
rect 2228 16201 2237 16235
rect 2237 16201 2271 16235
rect 2271 16201 2280 16235
rect 2228 16192 2280 16201
rect 2688 16192 2740 16244
rect 4160 16235 4212 16244
rect 4160 16201 4169 16235
rect 4169 16201 4203 16235
rect 4203 16201 4212 16235
rect 4160 16192 4212 16201
rect 5080 16235 5132 16244
rect 5080 16201 5089 16235
rect 5089 16201 5123 16235
rect 5123 16201 5132 16235
rect 5080 16192 5132 16201
rect 6092 16235 6144 16244
rect 6092 16201 6101 16235
rect 6101 16201 6135 16235
rect 6135 16201 6144 16235
rect 6092 16192 6144 16201
rect 10140 16192 10192 16244
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 5448 16056 5500 16108
rect 6092 16056 6144 16108
rect 10692 16056 10744 16108
rect 12440 16099 12492 16108
rect 12440 16065 12449 16099
rect 12449 16065 12483 16099
rect 12483 16065 12492 16099
rect 12440 16056 12492 16065
rect 1492 15988 1544 16040
rect 3976 15988 4028 16040
rect 4436 15988 4488 16040
rect 2964 15920 3016 15972
rect 4528 15895 4580 15904
rect 4528 15861 4537 15895
rect 4537 15861 4571 15895
rect 4571 15861 4580 15895
rect 4528 15852 4580 15861
rect 4988 15852 5040 15904
rect 5356 15852 5408 15904
rect 6828 15852 6880 15904
rect 7472 15988 7524 16040
rect 8208 15920 8260 15972
rect 11336 15920 11388 15972
rect 8024 15852 8076 15904
rect 8760 15895 8812 15904
rect 8760 15861 8769 15895
rect 8769 15861 8803 15895
rect 8803 15861 8812 15895
rect 8760 15852 8812 15861
rect 9772 15895 9824 15904
rect 9772 15861 9781 15895
rect 9781 15861 9815 15895
rect 9815 15861 9824 15895
rect 9772 15852 9824 15861
rect 11244 15895 11296 15904
rect 11244 15861 11253 15895
rect 11253 15861 11287 15895
rect 11287 15861 11296 15895
rect 11244 15852 11296 15861
rect 11796 15852 11848 15904
rect 12072 15895 12124 15904
rect 12072 15861 12081 15895
rect 12081 15861 12115 15895
rect 12115 15861 12124 15895
rect 12072 15852 12124 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1768 15648 1820 15700
rect 2780 15648 2832 15700
rect 4068 15691 4120 15700
rect 4068 15657 4077 15691
rect 4077 15657 4111 15691
rect 4111 15657 4120 15691
rect 4068 15648 4120 15657
rect 4160 15648 4212 15700
rect 5632 15648 5684 15700
rect 6736 15691 6788 15700
rect 6736 15657 6745 15691
rect 6745 15657 6779 15691
rect 6779 15657 6788 15691
rect 6736 15648 6788 15657
rect 7288 15691 7340 15700
rect 7288 15657 7297 15691
rect 7297 15657 7331 15691
rect 7331 15657 7340 15691
rect 7288 15648 7340 15657
rect 8668 15691 8720 15700
rect 8668 15657 8677 15691
rect 8677 15657 8711 15691
rect 8711 15657 8720 15691
rect 8668 15648 8720 15657
rect 10048 15691 10100 15700
rect 10048 15657 10057 15691
rect 10057 15657 10091 15691
rect 10091 15657 10100 15691
rect 10048 15648 10100 15657
rect 2964 15580 3016 15632
rect 5540 15580 5592 15632
rect 10692 15580 10744 15632
rect 11060 15580 11112 15632
rect 3056 15512 3108 15564
rect 5172 15512 5224 15564
rect 7656 15555 7708 15564
rect 7656 15521 7665 15555
rect 7665 15521 7699 15555
rect 7699 15521 7708 15555
rect 7656 15512 7708 15521
rect 9312 15555 9364 15564
rect 9312 15521 9321 15555
rect 9321 15521 9355 15555
rect 9355 15521 9364 15555
rect 9312 15512 9364 15521
rect 9956 15512 10008 15564
rect 12072 15512 12124 15564
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 1952 15351 2004 15360
rect 1952 15317 1961 15351
rect 1961 15317 1995 15351
rect 1995 15317 2004 15351
rect 1952 15308 2004 15317
rect 4068 15308 4120 15360
rect 7288 15444 7340 15496
rect 7012 15308 7064 15360
rect 8392 15351 8444 15360
rect 8392 15317 8401 15351
rect 8401 15317 8435 15351
rect 8435 15317 8444 15351
rect 8392 15308 8444 15317
rect 9220 15308 9272 15360
rect 12072 15351 12124 15360
rect 12072 15317 12081 15351
rect 12081 15317 12115 15351
rect 12115 15317 12124 15351
rect 12072 15308 12124 15317
rect 12808 15308 12860 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2044 15147 2096 15156
rect 2044 15113 2053 15147
rect 2053 15113 2087 15147
rect 2087 15113 2096 15147
rect 2044 15104 2096 15113
rect 3056 15147 3108 15156
rect 3056 15113 3065 15147
rect 3065 15113 3099 15147
rect 3099 15113 3108 15147
rect 3056 15104 3108 15113
rect 3516 15104 3568 15156
rect 4160 15104 4212 15156
rect 1952 14968 2004 15020
rect 3516 14968 3568 15020
rect 5540 14968 5592 15020
rect 6368 14968 6420 15020
rect 8116 15104 8168 15156
rect 9680 15104 9732 15156
rect 11060 15147 11112 15156
rect 11060 15113 11069 15147
rect 11069 15113 11103 15147
rect 11103 15113 11112 15147
rect 11060 15104 11112 15113
rect 10692 14968 10744 15020
rect 11888 15011 11940 15020
rect 11888 14977 11897 15011
rect 11897 14977 11931 15011
rect 11931 14977 11940 15011
rect 11888 14968 11940 14977
rect 2688 14900 2740 14952
rect 12808 14943 12860 14952
rect 4712 14832 4764 14884
rect 3516 14807 3568 14816
rect 3516 14773 3525 14807
rect 3525 14773 3559 14807
rect 3559 14773 3568 14807
rect 3516 14764 3568 14773
rect 3608 14764 3660 14816
rect 12808 14909 12817 14943
rect 12817 14909 12851 14943
rect 12851 14909 12860 14943
rect 12808 14900 12860 14909
rect 7656 14832 7708 14884
rect 8668 14832 8720 14884
rect 10048 14832 10100 14884
rect 10876 14832 10928 14884
rect 4896 14764 4948 14816
rect 5540 14807 5592 14816
rect 5540 14773 5549 14807
rect 5549 14773 5583 14807
rect 5583 14773 5592 14807
rect 5540 14764 5592 14773
rect 5632 14807 5684 14816
rect 5632 14773 5641 14807
rect 5641 14773 5675 14807
rect 5675 14773 5684 14807
rect 7288 14807 7340 14816
rect 5632 14764 5684 14773
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 9128 14807 9180 14816
rect 9128 14773 9137 14807
rect 9137 14773 9171 14807
rect 9171 14773 9180 14807
rect 9128 14764 9180 14773
rect 10784 14764 10836 14816
rect 11888 14764 11940 14816
rect 12256 14764 12308 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1400 14603 1452 14612
rect 1400 14569 1409 14603
rect 1409 14569 1443 14603
rect 1443 14569 1452 14603
rect 1400 14560 1452 14569
rect 2596 14560 2648 14612
rect 3148 14560 3200 14612
rect 4252 14603 4304 14612
rect 4252 14569 4261 14603
rect 4261 14569 4295 14603
rect 4295 14569 4304 14603
rect 4252 14560 4304 14569
rect 6368 14603 6420 14612
rect 6368 14569 6377 14603
rect 6377 14569 6411 14603
rect 6411 14569 6420 14603
rect 6368 14560 6420 14569
rect 6920 14560 6972 14612
rect 8668 14603 8720 14612
rect 8668 14569 8677 14603
rect 8677 14569 8711 14603
rect 8711 14569 8720 14603
rect 8668 14560 8720 14569
rect 8760 14603 8812 14612
rect 8760 14569 8769 14603
rect 8769 14569 8803 14603
rect 8803 14569 8812 14603
rect 9312 14603 9364 14612
rect 8760 14560 8812 14569
rect 9312 14569 9321 14603
rect 9321 14569 9355 14603
rect 9355 14569 9364 14603
rect 9312 14560 9364 14569
rect 11060 14560 11112 14612
rect 11888 14603 11940 14612
rect 11888 14569 11897 14603
rect 11897 14569 11931 14603
rect 11931 14569 11940 14603
rect 11888 14560 11940 14569
rect 12072 14560 12124 14612
rect 12624 14560 12676 14612
rect 2688 14492 2740 14544
rect 3976 14492 4028 14544
rect 7748 14492 7800 14544
rect 8116 14492 8168 14544
rect 9128 14492 9180 14544
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 3332 14424 3384 14476
rect 5080 14424 5132 14476
rect 5264 14467 5316 14476
rect 5264 14433 5298 14467
rect 5298 14433 5316 14467
rect 5264 14424 5316 14433
rect 10692 14492 10744 14544
rect 11152 14492 11204 14544
rect 10140 14424 10192 14476
rect 12900 14492 12952 14544
rect 23480 14467 23532 14476
rect 23480 14433 23489 14467
rect 23489 14433 23523 14467
rect 23523 14433 23532 14467
rect 23480 14424 23532 14433
rect 3056 14399 3108 14408
rect 3056 14365 3065 14399
rect 3065 14365 3099 14399
rect 3099 14365 3108 14399
rect 3056 14356 3108 14365
rect 4712 14399 4764 14408
rect 4712 14365 4721 14399
rect 4721 14365 4755 14399
rect 4755 14365 4764 14399
rect 4712 14356 4764 14365
rect 6920 14356 6972 14408
rect 7840 14399 7892 14408
rect 7840 14365 7849 14399
rect 7849 14365 7883 14399
rect 7883 14365 7892 14399
rect 7840 14356 7892 14365
rect 12256 14356 12308 14408
rect 12992 14399 13044 14408
rect 12992 14365 13001 14399
rect 13001 14365 13035 14399
rect 13035 14365 13044 14399
rect 12992 14356 13044 14365
rect 6000 14288 6052 14340
rect 8944 14288 8996 14340
rect 6368 14220 6420 14272
rect 24952 14220 25004 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2872 14016 2924 14068
rect 3332 14059 3384 14068
rect 3332 14025 3341 14059
rect 3341 14025 3375 14059
rect 3375 14025 3384 14059
rect 3332 14016 3384 14025
rect 4068 14059 4120 14068
rect 4068 14025 4077 14059
rect 4077 14025 4111 14059
rect 4111 14025 4120 14059
rect 4068 14016 4120 14025
rect 6644 14059 6696 14068
rect 6644 14025 6653 14059
rect 6653 14025 6687 14059
rect 6687 14025 6696 14059
rect 6644 14016 6696 14025
rect 7840 14016 7892 14068
rect 10048 14059 10100 14068
rect 10048 14025 10057 14059
rect 10057 14025 10091 14059
rect 10091 14025 10100 14059
rect 10048 14016 10100 14025
rect 11796 14059 11848 14068
rect 11796 14025 11805 14059
rect 11805 14025 11839 14059
rect 11839 14025 11848 14059
rect 11796 14016 11848 14025
rect 12256 14059 12308 14068
rect 12256 14025 12265 14059
rect 12265 14025 12299 14059
rect 12299 14025 12308 14059
rect 12256 14016 12308 14025
rect 12992 14016 13044 14068
rect 23480 14059 23532 14068
rect 23480 14025 23489 14059
rect 23489 14025 23523 14059
rect 23523 14025 23532 14059
rect 23480 14016 23532 14025
rect 3976 13948 4028 14000
rect 24860 13948 24912 14000
rect 3056 13880 3108 13932
rect 2780 13812 2832 13864
rect 6552 13880 6604 13932
rect 10692 13880 10744 13932
rect 1768 13676 1820 13728
rect 3056 13744 3108 13796
rect 3240 13744 3292 13796
rect 5264 13812 5316 13864
rect 5448 13744 5500 13796
rect 6920 13812 6972 13864
rect 7748 13855 7800 13864
rect 7748 13821 7757 13855
rect 7757 13821 7791 13855
rect 7791 13821 7800 13855
rect 7748 13812 7800 13821
rect 7840 13855 7892 13864
rect 7840 13821 7849 13855
rect 7849 13821 7883 13855
rect 7883 13821 7892 13855
rect 8116 13855 8168 13864
rect 7840 13812 7892 13821
rect 8116 13821 8150 13855
rect 8150 13821 8168 13855
rect 8116 13812 8168 13821
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 23664 13855 23716 13864
rect 23664 13821 23673 13855
rect 23673 13821 23707 13855
rect 23707 13821 23716 13855
rect 23664 13812 23716 13821
rect 6736 13744 6788 13796
rect 11704 13744 11756 13796
rect 2596 13676 2648 13728
rect 6276 13719 6328 13728
rect 6276 13685 6285 13719
rect 6285 13685 6319 13719
rect 6319 13685 6328 13719
rect 6276 13676 6328 13685
rect 6828 13719 6880 13728
rect 6828 13685 6837 13719
rect 6837 13685 6871 13719
rect 6871 13685 6880 13719
rect 6828 13676 6880 13685
rect 8116 13676 8168 13728
rect 9956 13676 10008 13728
rect 11152 13719 11204 13728
rect 11152 13685 11161 13719
rect 11161 13685 11195 13719
rect 11195 13685 11204 13719
rect 11152 13676 11204 13685
rect 11888 13676 11940 13728
rect 12440 13719 12492 13728
rect 12440 13685 12449 13719
rect 12449 13685 12483 13719
rect 12483 13685 12492 13719
rect 12440 13676 12492 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 3056 13472 3108 13524
rect 3884 13472 3936 13524
rect 5448 13472 5500 13524
rect 9312 13472 9364 13524
rect 9956 13472 10008 13524
rect 11152 13472 11204 13524
rect 11888 13515 11940 13524
rect 11888 13481 11897 13515
rect 11897 13481 11931 13515
rect 11931 13481 11940 13515
rect 11888 13472 11940 13481
rect 1952 13404 2004 13456
rect 3240 13404 3292 13456
rect 1768 13379 1820 13388
rect 1768 13345 1777 13379
rect 1777 13345 1811 13379
rect 1811 13345 1820 13379
rect 1768 13336 1820 13345
rect 2504 13336 2556 13388
rect 4068 13379 4120 13388
rect 4068 13345 4077 13379
rect 4077 13345 4111 13379
rect 4111 13345 4120 13379
rect 4068 13336 4120 13345
rect 3608 13268 3660 13320
rect 3884 13311 3936 13320
rect 3884 13277 3893 13311
rect 3893 13277 3927 13311
rect 3927 13277 3936 13311
rect 3884 13268 3936 13277
rect 5264 13268 5316 13320
rect 6368 13404 6420 13456
rect 10692 13404 10744 13456
rect 6000 13336 6052 13388
rect 8576 13336 8628 13388
rect 9312 13379 9364 13388
rect 9312 13345 9321 13379
rect 9321 13345 9355 13379
rect 9355 13345 9364 13379
rect 9312 13336 9364 13345
rect 10140 13336 10192 13388
rect 22284 13379 22336 13388
rect 22284 13345 22293 13379
rect 22293 13345 22327 13379
rect 22327 13345 22336 13379
rect 22284 13336 22336 13345
rect 7656 13268 7708 13320
rect 8208 13311 8260 13320
rect 8208 13277 8217 13311
rect 8217 13277 8251 13311
rect 8251 13277 8260 13311
rect 8208 13268 8260 13277
rect 6736 13243 6788 13252
rect 6736 13209 6745 13243
rect 6745 13209 6779 13243
rect 6779 13209 6788 13243
rect 6736 13200 6788 13209
rect 1768 13132 1820 13184
rect 4804 13132 4856 13184
rect 7380 13132 7432 13184
rect 11980 13132 12032 13184
rect 23480 13132 23532 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2320 12928 2372 12980
rect 3700 12928 3752 12980
rect 4068 12928 4120 12980
rect 8576 12903 8628 12912
rect 8576 12869 8585 12903
rect 8585 12869 8619 12903
rect 8619 12869 8628 12903
rect 8576 12860 8628 12869
rect 10140 12928 10192 12980
rect 10692 12928 10744 12980
rect 11980 12971 12032 12980
rect 11980 12937 11989 12971
rect 11989 12937 12023 12971
rect 12023 12937 12032 12971
rect 11980 12928 12032 12937
rect 11888 12903 11940 12912
rect 11888 12869 11897 12903
rect 11897 12869 11931 12903
rect 11931 12869 11940 12903
rect 11888 12860 11940 12869
rect 2872 12835 2924 12844
rect 2872 12801 2881 12835
rect 2881 12801 2915 12835
rect 2915 12801 2924 12835
rect 2872 12792 2924 12801
rect 7472 12792 7524 12844
rect 9772 12835 9824 12844
rect 9772 12801 9781 12835
rect 9781 12801 9815 12835
rect 9815 12801 9824 12835
rect 9772 12792 9824 12801
rect 1860 12724 1912 12776
rect 2596 12724 2648 12776
rect 3332 12767 3384 12776
rect 3332 12733 3366 12767
rect 3366 12733 3384 12767
rect 3332 12724 3384 12733
rect 4344 12656 4396 12708
rect 12164 12767 12216 12776
rect 12164 12733 12173 12767
rect 12173 12733 12207 12767
rect 12207 12733 12216 12767
rect 12164 12724 12216 12733
rect 12992 12767 13044 12776
rect 12992 12733 13001 12767
rect 13001 12733 13035 12767
rect 13035 12733 13044 12767
rect 12992 12724 13044 12733
rect 22284 12767 22336 12776
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 5540 12656 5592 12708
rect 8392 12656 8444 12708
rect 8668 12656 8720 12708
rect 9312 12656 9364 12708
rect 9680 12699 9732 12708
rect 9680 12665 9689 12699
rect 9689 12665 9723 12699
rect 9723 12665 9732 12699
rect 10048 12699 10100 12708
rect 9680 12656 9732 12665
rect 10048 12665 10082 12699
rect 10082 12665 10100 12699
rect 10048 12656 10100 12665
rect 11888 12656 11940 12708
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 2320 12588 2372 12640
rect 3424 12588 3476 12640
rect 4712 12588 4764 12640
rect 5080 12631 5132 12640
rect 5080 12597 5089 12631
rect 5089 12597 5123 12631
rect 5123 12597 5132 12631
rect 5080 12588 5132 12597
rect 6000 12588 6052 12640
rect 6736 12588 6788 12640
rect 7104 12631 7156 12640
rect 7104 12597 7113 12631
rect 7113 12597 7147 12631
rect 7147 12597 7156 12631
rect 7104 12588 7156 12597
rect 7380 12588 7432 12640
rect 8208 12631 8260 12640
rect 8208 12597 8217 12631
rect 8217 12597 8251 12631
rect 8251 12597 8260 12631
rect 8208 12588 8260 12597
rect 8760 12631 8812 12640
rect 8760 12597 8769 12631
rect 8769 12597 8803 12631
rect 8803 12597 8812 12631
rect 8760 12588 8812 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 3332 12384 3384 12436
rect 4160 12384 4212 12436
rect 4344 12384 4396 12436
rect 5264 12384 5316 12436
rect 2320 12248 2372 12300
rect 4344 12248 4396 12300
rect 5264 12248 5316 12300
rect 6828 12384 6880 12436
rect 7012 12384 7064 12436
rect 7472 12384 7524 12436
rect 7932 12384 7984 12436
rect 8760 12384 8812 12436
rect 10048 12384 10100 12436
rect 10600 12316 10652 12368
rect 6092 12248 6144 12300
rect 9772 12248 9824 12300
rect 11612 12248 11664 12300
rect 12716 12248 12768 12300
rect 21732 12291 21784 12300
rect 21732 12257 21741 12291
rect 21741 12257 21775 12291
rect 21775 12257 21784 12291
rect 21732 12248 21784 12257
rect 3056 12223 3108 12232
rect 3056 12189 3065 12223
rect 3065 12189 3099 12223
rect 3099 12189 3108 12223
rect 3056 12180 3108 12189
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 8484 12223 8536 12232
rect 8484 12189 8493 12223
rect 8493 12189 8527 12223
rect 8527 12189 8536 12223
rect 8484 12180 8536 12189
rect 9128 12223 9180 12232
rect 7748 12112 7800 12164
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 10692 12180 10744 12232
rect 11980 12223 12032 12232
rect 11980 12189 11989 12223
rect 11989 12189 12023 12223
rect 12023 12189 12032 12223
rect 11980 12180 12032 12189
rect 1952 12044 2004 12096
rect 2964 12044 3016 12096
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 4344 12044 4396 12096
rect 4804 12044 4856 12096
rect 5172 12044 5224 12096
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 9680 12044 9732 12096
rect 11152 12044 11204 12096
rect 13268 12044 13320 12096
rect 21916 12087 21968 12096
rect 21916 12053 21925 12087
rect 21925 12053 21959 12087
rect 21959 12053 21968 12087
rect 21916 12044 21968 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2412 11840 2464 11892
rect 3516 11840 3568 11892
rect 1676 11747 1728 11756
rect 1676 11713 1685 11747
rect 1685 11713 1719 11747
rect 1719 11713 1728 11747
rect 1676 11704 1728 11713
rect 3240 11747 3292 11756
rect 3240 11713 3249 11747
rect 3249 11713 3283 11747
rect 3283 11713 3292 11747
rect 3240 11704 3292 11713
rect 6000 11840 6052 11892
rect 6644 11840 6696 11892
rect 7748 11883 7800 11892
rect 7748 11849 7757 11883
rect 7757 11849 7791 11883
rect 7791 11849 7800 11883
rect 7748 11840 7800 11849
rect 8760 11840 8812 11892
rect 11980 11840 12032 11892
rect 21732 11815 21784 11824
rect 21732 11781 21741 11815
rect 21741 11781 21775 11815
rect 21775 11781 21784 11815
rect 21732 11772 21784 11781
rect 3332 11636 3384 11688
rect 9772 11704 9824 11756
rect 10692 11747 10744 11756
rect 10692 11713 10701 11747
rect 10701 11713 10735 11747
rect 10735 11713 10744 11747
rect 10692 11704 10744 11713
rect 2596 11611 2648 11620
rect 2596 11577 2605 11611
rect 2605 11577 2639 11611
rect 2639 11577 2648 11611
rect 2596 11568 2648 11577
rect 5540 11636 5592 11688
rect 12716 11679 12768 11688
rect 12716 11645 12725 11679
rect 12725 11645 12759 11679
rect 12759 11645 12768 11679
rect 12716 11636 12768 11645
rect 5632 11568 5684 11620
rect 2320 11500 2372 11552
rect 2964 11500 3016 11552
rect 5172 11500 5224 11552
rect 8484 11568 8536 11620
rect 8852 11611 8904 11620
rect 8852 11577 8861 11611
rect 8861 11577 8895 11611
rect 8895 11577 8904 11611
rect 8852 11568 8904 11577
rect 9220 11568 9272 11620
rect 11152 11568 11204 11620
rect 6092 11500 6144 11552
rect 6276 11543 6328 11552
rect 6276 11509 6285 11543
rect 6285 11509 6319 11543
rect 6319 11509 6328 11543
rect 6276 11500 6328 11509
rect 6920 11500 6972 11552
rect 10140 11543 10192 11552
rect 10140 11509 10149 11543
rect 10149 11509 10183 11543
rect 10183 11509 10192 11543
rect 10140 11500 10192 11509
rect 10692 11500 10744 11552
rect 12992 11500 13044 11552
rect 13728 11500 13780 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 3148 11296 3200 11348
rect 3332 11339 3384 11348
rect 3332 11305 3341 11339
rect 3341 11305 3375 11339
rect 3375 11305 3384 11339
rect 3332 11296 3384 11305
rect 5264 11339 5316 11348
rect 5264 11305 5273 11339
rect 5273 11305 5307 11339
rect 5307 11305 5316 11339
rect 5264 11296 5316 11305
rect 6276 11296 6328 11348
rect 7104 11296 7156 11348
rect 8300 11296 8352 11348
rect 8484 11296 8536 11348
rect 11244 11339 11296 11348
rect 11244 11305 11253 11339
rect 11253 11305 11287 11339
rect 11287 11305 11296 11339
rect 11244 11296 11296 11305
rect 11612 11296 11664 11348
rect 12808 11339 12860 11348
rect 12808 11305 12817 11339
rect 12817 11305 12851 11339
rect 12851 11305 12860 11339
rect 12808 11296 12860 11305
rect 2504 11228 2556 11280
rect 6000 11228 6052 11280
rect 8116 11271 8168 11280
rect 8116 11237 8150 11271
rect 8150 11237 8168 11271
rect 8116 11228 8168 11237
rect 1768 11160 1820 11212
rect 2964 11160 3016 11212
rect 3148 11160 3200 11212
rect 4160 11160 4212 11212
rect 5632 11203 5684 11212
rect 5632 11169 5641 11203
rect 5641 11169 5675 11203
rect 5675 11169 5684 11203
rect 5632 11160 5684 11169
rect 4068 11092 4120 11144
rect 4620 11135 4672 11144
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 9128 11160 9180 11212
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 11060 11203 11112 11212
rect 11060 11169 11069 11203
rect 11069 11169 11103 11203
rect 11103 11169 11112 11203
rect 11060 11160 11112 11169
rect 11612 11203 11664 11212
rect 11612 11169 11621 11203
rect 11621 11169 11655 11203
rect 11655 11169 11664 11203
rect 11612 11160 11664 11169
rect 13176 11203 13228 11212
rect 13176 11169 13185 11203
rect 13185 11169 13219 11203
rect 13219 11169 13228 11203
rect 13176 11160 13228 11169
rect 13452 11160 13504 11212
rect 4620 11092 4672 11101
rect 9956 11092 10008 11144
rect 10692 11092 10744 11144
rect 13084 11092 13136 11144
rect 9220 11067 9272 11076
rect 1308 10956 1360 11008
rect 3332 10956 3384 11008
rect 7380 10999 7432 11008
rect 7380 10965 7389 10999
rect 7389 10965 7423 10999
rect 7423 10965 7432 10999
rect 7380 10956 7432 10965
rect 8208 10956 8260 11008
rect 9220 11033 9229 11067
rect 9229 11033 9263 11067
rect 9263 11033 9272 11067
rect 9220 11024 9272 11033
rect 9772 11024 9824 11076
rect 10968 11024 11020 11076
rect 12808 10956 12860 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 3056 10795 3108 10804
rect 3056 10761 3065 10795
rect 3065 10761 3099 10795
rect 3099 10761 3108 10795
rect 3056 10752 3108 10761
rect 4252 10752 4304 10804
rect 4620 10752 4672 10804
rect 5540 10752 5592 10804
rect 6000 10795 6052 10804
rect 6000 10761 6009 10795
rect 6009 10761 6043 10795
rect 6043 10761 6052 10795
rect 6000 10752 6052 10761
rect 6920 10752 6972 10804
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 2596 10548 2648 10600
rect 3056 10548 3108 10600
rect 6000 10548 6052 10600
rect 6184 10548 6236 10600
rect 7380 10752 7432 10804
rect 7932 10752 7984 10804
rect 8392 10752 8444 10804
rect 9680 10752 9732 10804
rect 12532 10752 12584 10804
rect 13820 10752 13872 10804
rect 7748 10727 7800 10736
rect 7748 10693 7757 10727
rect 7757 10693 7791 10727
rect 7791 10693 7800 10727
rect 7748 10684 7800 10693
rect 12256 10684 12308 10736
rect 8116 10616 8168 10668
rect 9496 10616 9548 10668
rect 11060 10616 11112 10668
rect 12348 10616 12400 10668
rect 13084 10659 13136 10668
rect 13084 10625 13093 10659
rect 13093 10625 13127 10659
rect 13127 10625 13136 10659
rect 13084 10616 13136 10625
rect 12256 10548 12308 10600
rect 12808 10591 12860 10600
rect 12808 10557 12817 10591
rect 12817 10557 12851 10591
rect 12851 10557 12860 10591
rect 12808 10548 12860 10557
rect 1768 10412 1820 10464
rect 5172 10480 5224 10532
rect 4712 10412 4764 10464
rect 6920 10480 6972 10532
rect 8392 10480 8444 10532
rect 6184 10412 6236 10464
rect 9128 10455 9180 10464
rect 9128 10421 9137 10455
rect 9137 10421 9171 10455
rect 9171 10421 9180 10455
rect 9128 10412 9180 10421
rect 9404 10412 9456 10464
rect 9864 10412 9916 10464
rect 9956 10412 10008 10464
rect 11060 10455 11112 10464
rect 11060 10421 11069 10455
rect 11069 10421 11103 10455
rect 11103 10421 11112 10455
rect 11060 10412 11112 10421
rect 11152 10455 11204 10464
rect 11152 10421 11161 10455
rect 11161 10421 11195 10455
rect 11195 10421 11204 10455
rect 11152 10412 11204 10421
rect 11612 10412 11664 10464
rect 13452 10455 13504 10464
rect 13452 10421 13461 10455
rect 13461 10421 13495 10455
rect 13495 10421 13504 10455
rect 13452 10412 13504 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1768 10251 1820 10260
rect 1768 10217 1777 10251
rect 1777 10217 1811 10251
rect 1811 10217 1820 10251
rect 1768 10208 1820 10217
rect 4068 10251 4120 10260
rect 4068 10217 4077 10251
rect 4077 10217 4111 10251
rect 4111 10217 4120 10251
rect 4068 10208 4120 10217
rect 6092 10208 6144 10260
rect 7196 10208 7248 10260
rect 7932 10251 7984 10260
rect 7932 10217 7941 10251
rect 7941 10217 7975 10251
rect 7975 10217 7984 10251
rect 7932 10208 7984 10217
rect 8116 10208 8168 10260
rect 10048 10208 10100 10260
rect 10692 10208 10744 10260
rect 12348 10251 12400 10260
rect 12348 10217 12357 10251
rect 12357 10217 12391 10251
rect 12391 10217 12400 10251
rect 12348 10208 12400 10217
rect 1492 10140 1544 10192
rect 4160 10140 4212 10192
rect 6368 10140 6420 10192
rect 7748 10140 7800 10192
rect 9404 10140 9456 10192
rect 11060 10140 11112 10192
rect 13176 10208 13228 10260
rect 2412 10115 2464 10124
rect 2412 10081 2421 10115
rect 2421 10081 2455 10115
rect 2455 10081 2464 10115
rect 2412 10072 2464 10081
rect 4068 10072 4120 10124
rect 7380 10072 7432 10124
rect 7840 10072 7892 10124
rect 9128 10072 9180 10124
rect 11244 10115 11296 10124
rect 11244 10081 11278 10115
rect 11278 10081 11296 10115
rect 11244 10072 11296 10081
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 2964 9936 3016 9988
rect 4804 10004 4856 10056
rect 6092 10047 6144 10056
rect 6092 10013 6101 10047
rect 6101 10013 6135 10047
rect 6135 10013 6144 10047
rect 6092 10004 6144 10013
rect 6184 10047 6236 10056
rect 6184 10013 6193 10047
rect 6193 10013 6227 10047
rect 6227 10013 6236 10047
rect 7196 10047 7248 10056
rect 6184 10004 6236 10013
rect 6736 9979 6788 9988
rect 2044 9911 2096 9920
rect 2044 9877 2053 9911
rect 2053 9877 2087 9911
rect 2087 9877 2096 9911
rect 2044 9868 2096 9877
rect 2504 9868 2556 9920
rect 3424 9868 3476 9920
rect 5172 9911 5224 9920
rect 5172 9877 5181 9911
rect 5181 9877 5215 9911
rect 5215 9877 5224 9911
rect 5172 9868 5224 9877
rect 6736 9945 6745 9979
rect 6745 9945 6779 9979
rect 6779 9945 6788 9979
rect 6736 9936 6788 9945
rect 7196 10013 7205 10047
rect 7205 10013 7239 10047
rect 7239 10013 7248 10047
rect 7196 10004 7248 10013
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 10968 10047 11020 10056
rect 10968 10013 10977 10047
rect 10977 10013 11011 10047
rect 11011 10013 11020 10047
rect 10968 10004 11020 10013
rect 13176 10047 13228 10056
rect 13176 10013 13185 10047
rect 13185 10013 13219 10047
rect 13219 10013 13228 10047
rect 13176 10004 13228 10013
rect 9404 9868 9456 9920
rect 13728 9868 13780 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1768 9664 1820 9716
rect 2596 9664 2648 9716
rect 2964 9664 3016 9716
rect 3056 9664 3108 9716
rect 9496 9664 9548 9716
rect 11244 9664 11296 9716
rect 4068 9639 4120 9648
rect 4068 9605 4077 9639
rect 4077 9605 4111 9639
rect 4111 9605 4120 9639
rect 4068 9596 4120 9605
rect 1400 9528 1452 9580
rect 1860 9571 1912 9580
rect 1860 9537 1869 9571
rect 1869 9537 1903 9571
rect 1903 9537 1912 9571
rect 1860 9528 1912 9537
rect 2872 9528 2924 9580
rect 6184 9596 6236 9648
rect 4528 9528 4580 9580
rect 5264 9528 5316 9580
rect 5540 9528 5592 9580
rect 3424 9324 3476 9376
rect 7196 9460 7248 9512
rect 10692 9460 10744 9512
rect 10968 9460 11020 9512
rect 3792 9324 3844 9376
rect 4896 9392 4948 9444
rect 6368 9392 6420 9444
rect 7472 9392 7524 9444
rect 9772 9392 9824 9444
rect 4160 9324 4212 9376
rect 6092 9367 6144 9376
rect 6092 9333 6101 9367
rect 6101 9333 6135 9367
rect 6135 9333 6144 9367
rect 6092 9324 6144 9333
rect 6184 9324 6236 9376
rect 12440 9639 12492 9648
rect 12440 9605 12449 9639
rect 12449 9605 12483 9639
rect 12483 9605 12492 9639
rect 12440 9596 12492 9605
rect 13728 9639 13780 9648
rect 13728 9605 13737 9639
rect 13737 9605 13771 9639
rect 13771 9605 13780 9639
rect 13728 9596 13780 9605
rect 12348 9528 12400 9580
rect 12808 9528 12860 9580
rect 12164 9503 12216 9512
rect 12164 9469 12173 9503
rect 12173 9469 12207 9503
rect 12207 9469 12216 9503
rect 12164 9460 12216 9469
rect 12992 9392 13044 9444
rect 7104 9367 7156 9376
rect 7104 9333 7113 9367
rect 7113 9333 7147 9367
rect 7147 9333 7156 9367
rect 7104 9324 7156 9333
rect 7380 9367 7432 9376
rect 7380 9333 7389 9367
rect 7389 9333 7423 9367
rect 7423 9333 7432 9367
rect 7380 9324 7432 9333
rect 8852 9324 8904 9376
rect 10048 9367 10100 9376
rect 10048 9333 10057 9367
rect 10057 9333 10091 9367
rect 10091 9333 10100 9367
rect 10048 9324 10100 9333
rect 12440 9324 12492 9376
rect 13176 9324 13228 9376
rect 13268 9324 13320 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1584 9120 1636 9172
rect 2044 9120 2096 9172
rect 2872 9120 2924 9172
rect 3056 9120 3108 9172
rect 4068 9120 4120 9172
rect 6552 9120 6604 9172
rect 8116 9120 8168 9172
rect 9128 9120 9180 9172
rect 10140 9120 10192 9172
rect 12808 9163 12860 9172
rect 12808 9129 12817 9163
rect 12817 9129 12851 9163
rect 12851 9129 12860 9163
rect 12808 9120 12860 9129
rect 13728 9120 13780 9172
rect 2688 9052 2740 9104
rect 4344 9095 4396 9104
rect 4344 9061 4353 9095
rect 4353 9061 4387 9095
rect 4387 9061 4396 9095
rect 4344 9052 4396 9061
rect 4896 9052 4948 9104
rect 7380 9052 7432 9104
rect 8484 9052 8536 9104
rect 12440 9095 12492 9104
rect 12440 9061 12449 9095
rect 12449 9061 12483 9095
rect 12483 9061 12492 9095
rect 12440 9052 12492 9061
rect 13452 9052 13504 9104
rect 1952 8984 2004 9036
rect 2504 8984 2556 9036
rect 1768 8916 1820 8968
rect 3976 8984 4028 9036
rect 4712 8984 4764 9036
rect 6368 8984 6420 9036
rect 6736 8984 6788 9036
rect 8024 8984 8076 9036
rect 4344 8916 4396 8968
rect 9680 8984 9732 9036
rect 10692 8984 10744 9036
rect 11520 8984 11572 9036
rect 9772 8959 9824 8968
rect 3056 8780 3108 8832
rect 5172 8848 5224 8900
rect 9772 8925 9781 8959
rect 9781 8925 9815 8959
rect 9815 8925 9824 8959
rect 9772 8916 9824 8925
rect 13268 8916 13320 8968
rect 13636 8959 13688 8968
rect 13636 8925 13645 8959
rect 13645 8925 13679 8959
rect 13679 8925 13688 8959
rect 13636 8916 13688 8925
rect 9312 8848 9364 8900
rect 4804 8823 4856 8832
rect 4804 8789 4813 8823
rect 4813 8789 4847 8823
rect 4847 8789 4856 8823
rect 4804 8780 4856 8789
rect 5356 8780 5408 8832
rect 7748 8823 7800 8832
rect 7748 8789 7757 8823
rect 7757 8789 7791 8823
rect 7791 8789 7800 8823
rect 7748 8780 7800 8789
rect 8024 8823 8076 8832
rect 8024 8789 8033 8823
rect 8033 8789 8067 8823
rect 8067 8789 8076 8823
rect 8024 8780 8076 8789
rect 9496 8780 9548 8832
rect 12164 8823 12216 8832
rect 12164 8789 12173 8823
rect 12173 8789 12207 8823
rect 12207 8789 12216 8823
rect 12164 8780 12216 8789
rect 13728 8780 13780 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2872 8576 2924 8628
rect 3700 8619 3752 8628
rect 3700 8585 3709 8619
rect 3709 8585 3743 8619
rect 3743 8585 3752 8619
rect 3700 8576 3752 8585
rect 3976 8619 4028 8628
rect 3976 8585 3985 8619
rect 3985 8585 4019 8619
rect 4019 8585 4028 8619
rect 3976 8576 4028 8585
rect 4712 8619 4764 8628
rect 4712 8585 4721 8619
rect 4721 8585 4755 8619
rect 4755 8585 4764 8619
rect 4712 8576 4764 8585
rect 6460 8576 6512 8628
rect 7104 8576 7156 8628
rect 8300 8619 8352 8628
rect 8300 8585 8309 8619
rect 8309 8585 8343 8619
rect 8343 8585 8352 8619
rect 8300 8576 8352 8585
rect 8852 8619 8904 8628
rect 8852 8585 8861 8619
rect 8861 8585 8895 8619
rect 8895 8585 8904 8619
rect 8852 8576 8904 8585
rect 9772 8576 9824 8628
rect 5172 8551 5224 8560
rect 5172 8517 5181 8551
rect 5181 8517 5215 8551
rect 5215 8517 5224 8551
rect 5172 8508 5224 8517
rect 1860 8440 1912 8492
rect 4436 8440 4488 8492
rect 6000 8440 6052 8492
rect 3056 8372 3108 8424
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 6920 8440 6972 8492
rect 8300 8440 8352 8492
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 10048 8440 10100 8492
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 12624 8508 12676 8560
rect 5540 8372 5592 8381
rect 7748 8372 7800 8424
rect 9680 8372 9732 8424
rect 10140 8372 10192 8424
rect 11520 8415 11572 8424
rect 11520 8381 11529 8415
rect 11529 8381 11563 8415
rect 11563 8381 11572 8415
rect 11520 8372 11572 8381
rect 12256 8415 12308 8424
rect 12256 8381 12265 8415
rect 12265 8381 12299 8415
rect 12299 8381 12308 8415
rect 12256 8372 12308 8381
rect 5356 8304 5408 8356
rect 2412 8236 2464 8288
rect 2964 8236 3016 8288
rect 7840 8304 7892 8356
rect 8484 8304 8536 8356
rect 7012 8236 7064 8288
rect 9036 8236 9088 8288
rect 13636 8576 13688 8628
rect 13912 8576 13964 8628
rect 14372 8576 14424 8628
rect 17132 8551 17184 8560
rect 17132 8517 17141 8551
rect 17141 8517 17175 8551
rect 17175 8517 17184 8551
rect 17132 8508 17184 8517
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 14004 8415 14056 8424
rect 14004 8381 14013 8415
rect 14013 8381 14047 8415
rect 14047 8381 14056 8415
rect 14004 8372 14056 8381
rect 15752 8415 15804 8424
rect 15752 8381 15761 8415
rect 15761 8381 15795 8415
rect 15795 8381 15804 8415
rect 15752 8372 15804 8381
rect 13544 8304 13596 8356
rect 10692 8236 10744 8288
rect 13176 8236 13228 8288
rect 13452 8279 13504 8288
rect 13452 8245 13461 8279
rect 13461 8245 13495 8279
rect 13495 8245 13504 8279
rect 13452 8236 13504 8245
rect 15660 8279 15712 8288
rect 15660 8245 15669 8279
rect 15669 8245 15703 8279
rect 15703 8245 15712 8279
rect 15660 8236 15712 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2780 8032 2832 8084
rect 4344 8075 4396 8084
rect 4344 8041 4353 8075
rect 4353 8041 4387 8075
rect 4387 8041 4396 8075
rect 4344 8032 4396 8041
rect 5448 8032 5500 8084
rect 1860 7964 1912 8016
rect 2504 7964 2556 8016
rect 5080 8007 5132 8016
rect 5080 7973 5114 8007
rect 5114 7973 5132 8007
rect 5080 7964 5132 7973
rect 5264 7964 5316 8016
rect 6736 8032 6788 8084
rect 7656 8032 7708 8084
rect 9496 8032 9548 8084
rect 9680 8032 9732 8084
rect 12992 8032 13044 8084
rect 12164 7964 12216 8016
rect 13544 7964 13596 8016
rect 15752 8007 15804 8016
rect 15752 7973 15761 8007
rect 15761 7973 15795 8007
rect 15795 7973 15804 8007
rect 15752 7964 15804 7973
rect 2228 7896 2280 7948
rect 2780 7896 2832 7948
rect 7472 7939 7524 7948
rect 7472 7905 7506 7939
rect 7506 7905 7524 7939
rect 7472 7896 7524 7905
rect 10692 7896 10744 7948
rect 12992 7896 13044 7948
rect 7196 7871 7248 7880
rect 2412 7760 2464 7812
rect 4252 7760 4304 7812
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 13176 7828 13228 7880
rect 12532 7803 12584 7812
rect 12532 7769 12541 7803
rect 12541 7769 12575 7803
rect 12575 7769 12584 7803
rect 12532 7760 12584 7769
rect 15844 7828 15896 7880
rect 5448 7692 5500 7744
rect 7012 7692 7064 7744
rect 8576 7735 8628 7744
rect 8576 7701 8585 7735
rect 8585 7701 8619 7735
rect 8619 7701 8628 7735
rect 8576 7692 8628 7701
rect 9036 7692 9088 7744
rect 9312 7735 9364 7744
rect 9312 7701 9321 7735
rect 9321 7701 9355 7735
rect 9355 7701 9364 7735
rect 9312 7692 9364 7701
rect 12900 7692 12952 7744
rect 13820 7692 13872 7744
rect 14096 7692 14148 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2596 7488 2648 7540
rect 2780 7488 2832 7540
rect 3148 7488 3200 7540
rect 4160 7488 4212 7540
rect 2872 7352 2924 7404
rect 2780 7327 2832 7336
rect 2780 7293 2789 7327
rect 2789 7293 2823 7327
rect 2823 7293 2832 7327
rect 2780 7284 2832 7293
rect 7472 7488 7524 7540
rect 6828 7395 6880 7404
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 8760 7488 8812 7540
rect 9680 7531 9732 7540
rect 9680 7497 9689 7531
rect 9689 7497 9723 7531
rect 9723 7497 9732 7531
rect 9680 7488 9732 7497
rect 12164 7488 12216 7540
rect 12992 7531 13044 7540
rect 12992 7497 13001 7531
rect 13001 7497 13035 7531
rect 13035 7497 13044 7531
rect 12992 7488 13044 7497
rect 14464 7488 14516 7540
rect 15844 7531 15896 7540
rect 15844 7497 15853 7531
rect 15853 7497 15887 7531
rect 15887 7497 15896 7531
rect 15844 7488 15896 7497
rect 13452 7352 13504 7404
rect 13544 7352 13596 7404
rect 3056 7216 3108 7268
rect 3884 7216 3936 7268
rect 5264 7216 5316 7268
rect 8576 7284 8628 7336
rect 9680 7284 9732 7336
rect 10784 7284 10836 7336
rect 11244 7327 11296 7336
rect 11244 7293 11253 7327
rect 11253 7293 11287 7327
rect 11287 7293 11296 7327
rect 11244 7284 11296 7293
rect 16488 7395 16540 7404
rect 16488 7361 16497 7395
rect 16497 7361 16531 7395
rect 16531 7361 16540 7395
rect 16488 7352 16540 7361
rect 14096 7216 14148 7268
rect 15660 7216 15712 7268
rect 16488 7216 16540 7268
rect 2504 7191 2556 7200
rect 2504 7157 2513 7191
rect 2513 7157 2547 7191
rect 2547 7157 2556 7191
rect 2504 7148 2556 7157
rect 3516 7148 3568 7200
rect 4804 7148 4856 7200
rect 5172 7191 5224 7200
rect 5172 7157 5181 7191
rect 5181 7157 5215 7191
rect 5215 7157 5224 7191
rect 5172 7148 5224 7157
rect 5448 7148 5500 7200
rect 7196 7148 7248 7200
rect 8208 7148 8260 7200
rect 9404 7191 9456 7200
rect 9404 7157 9413 7191
rect 9413 7157 9447 7191
rect 9447 7157 9456 7191
rect 9404 7148 9456 7157
rect 10140 7148 10192 7200
rect 10784 7191 10836 7200
rect 10784 7157 10793 7191
rect 10793 7157 10827 7191
rect 10827 7157 10836 7191
rect 10784 7148 10836 7157
rect 13176 7148 13228 7200
rect 15936 7191 15988 7200
rect 15936 7157 15945 7191
rect 15945 7157 15979 7191
rect 15979 7157 15988 7191
rect 15936 7148 15988 7157
rect 16396 7191 16448 7200
rect 16396 7157 16405 7191
rect 16405 7157 16439 7191
rect 16439 7157 16448 7191
rect 16396 7148 16448 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 2872 6987 2924 6996
rect 2872 6953 2881 6987
rect 2881 6953 2915 6987
rect 2915 6953 2924 6987
rect 2872 6944 2924 6953
rect 2320 6876 2372 6928
rect 5080 6944 5132 6996
rect 9036 6944 9088 6996
rect 9680 6944 9732 6996
rect 3884 6919 3936 6928
rect 3884 6885 3893 6919
rect 3893 6885 3927 6919
rect 3927 6885 3936 6919
rect 3884 6876 3936 6885
rect 10140 6876 10192 6928
rect 13544 6944 13596 6996
rect 15660 6944 15712 6996
rect 1768 6851 1820 6860
rect 1768 6817 1777 6851
rect 1777 6817 1811 6851
rect 1811 6817 1820 6851
rect 1768 6808 1820 6817
rect 2228 6808 2280 6860
rect 1584 6740 1636 6792
rect 4344 6808 4396 6860
rect 5448 6851 5500 6860
rect 5448 6817 5457 6851
rect 5457 6817 5491 6851
rect 5491 6817 5500 6851
rect 5448 6808 5500 6817
rect 6736 6808 6788 6860
rect 7104 6851 7156 6860
rect 7104 6817 7113 6851
rect 7113 6817 7147 6851
rect 7147 6817 7156 6851
rect 7104 6808 7156 6817
rect 8116 6851 8168 6860
rect 8116 6817 8125 6851
rect 8125 6817 8159 6851
rect 8159 6817 8168 6851
rect 8116 6808 8168 6817
rect 8208 6851 8260 6860
rect 8208 6817 8217 6851
rect 8217 6817 8251 6851
rect 8251 6817 8260 6851
rect 8208 6808 8260 6817
rect 10324 6851 10376 6860
rect 10324 6817 10358 6851
rect 10358 6817 10376 6851
rect 10324 6808 10376 6817
rect 12256 6808 12308 6860
rect 12900 6808 12952 6860
rect 14832 6808 14884 6860
rect 16396 6876 16448 6928
rect 8576 6740 8628 6792
rect 7748 6715 7800 6724
rect 7748 6681 7757 6715
rect 7757 6681 7791 6715
rect 7791 6681 7800 6715
rect 7748 6672 7800 6681
rect 8300 6672 8352 6724
rect 1400 6647 1452 6656
rect 1400 6613 1409 6647
rect 1409 6613 1443 6647
rect 1443 6613 1452 6647
rect 1400 6604 1452 6613
rect 2412 6647 2464 6656
rect 2412 6613 2421 6647
rect 2421 6613 2455 6647
rect 2455 6613 2464 6647
rect 2412 6604 2464 6613
rect 3516 6647 3568 6656
rect 3516 6613 3525 6647
rect 3525 6613 3559 6647
rect 3559 6613 3568 6647
rect 3516 6604 3568 6613
rect 5448 6604 5500 6656
rect 6092 6604 6144 6656
rect 7472 6647 7524 6656
rect 7472 6613 7481 6647
rect 7481 6613 7515 6647
rect 7515 6613 7524 6647
rect 7472 6604 7524 6613
rect 8760 6647 8812 6656
rect 8760 6613 8769 6647
rect 8769 6613 8803 6647
rect 8803 6613 8812 6647
rect 8760 6604 8812 6613
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 9128 6604 9180 6613
rect 12808 6740 12860 6792
rect 15752 6808 15804 6860
rect 17868 6851 17920 6860
rect 17868 6817 17877 6851
rect 17877 6817 17911 6851
rect 17911 6817 17920 6851
rect 17868 6808 17920 6817
rect 15660 6783 15712 6792
rect 15660 6749 15676 6783
rect 15676 6749 15710 6783
rect 15710 6749 15712 6783
rect 18144 6783 18196 6792
rect 15660 6740 15712 6749
rect 18144 6749 18153 6783
rect 18153 6749 18187 6783
rect 18187 6749 18196 6783
rect 18144 6740 18196 6749
rect 10784 6604 10836 6656
rect 11428 6647 11480 6656
rect 11428 6613 11437 6647
rect 11437 6613 11471 6647
rect 11471 6613 11480 6647
rect 11428 6604 11480 6613
rect 11612 6604 11664 6656
rect 14096 6604 14148 6656
rect 16580 6604 16632 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 1768 6400 1820 6452
rect 4160 6400 4212 6452
rect 6828 6443 6880 6452
rect 4344 6332 4396 6384
rect 2044 6264 2096 6316
rect 2412 6264 2464 6316
rect 2688 6196 2740 6248
rect 6828 6409 6837 6443
rect 6837 6409 6871 6443
rect 6871 6409 6880 6443
rect 6828 6400 6880 6409
rect 8116 6400 8168 6452
rect 8576 6400 8628 6452
rect 9772 6400 9824 6452
rect 10324 6400 10376 6452
rect 11428 6400 11480 6452
rect 11888 6400 11940 6452
rect 13084 6400 13136 6452
rect 13452 6400 13504 6452
rect 14832 6400 14884 6452
rect 15660 6400 15712 6452
rect 17868 6400 17920 6452
rect 5540 6332 5592 6384
rect 6736 6332 6788 6384
rect 6000 6264 6052 6316
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 12808 6307 12860 6316
rect 7472 6196 7524 6248
rect 12808 6273 12817 6307
rect 12817 6273 12851 6307
rect 12851 6273 12860 6307
rect 12808 6264 12860 6273
rect 15752 6264 15804 6316
rect 16120 6264 16172 6316
rect 1676 6128 1728 6180
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 2412 6060 2464 6112
rect 7104 6128 7156 6180
rect 9404 6196 9456 6248
rect 13084 6239 13136 6248
rect 13084 6205 13118 6239
rect 13118 6205 13136 6239
rect 13084 6196 13136 6205
rect 13636 6196 13688 6248
rect 14556 6196 14608 6248
rect 16580 6239 16632 6248
rect 16580 6205 16589 6239
rect 16589 6205 16623 6239
rect 16623 6205 16632 6239
rect 16580 6196 16632 6205
rect 19524 6239 19576 6248
rect 19524 6205 19533 6239
rect 19533 6205 19567 6239
rect 19567 6205 19576 6239
rect 19524 6196 19576 6205
rect 10784 6103 10836 6112
rect 10784 6069 10793 6103
rect 10793 6069 10827 6103
rect 10827 6069 10836 6103
rect 10784 6060 10836 6069
rect 11152 6103 11204 6112
rect 11152 6069 11161 6103
rect 11161 6069 11195 6103
rect 11195 6069 11204 6103
rect 11152 6060 11204 6069
rect 12900 6060 12952 6112
rect 14740 6060 14792 6112
rect 16856 6171 16908 6180
rect 16856 6137 16865 6171
rect 16865 6137 16899 6171
rect 16899 6137 16908 6171
rect 16856 6128 16908 6137
rect 20536 6128 20588 6180
rect 16120 6103 16172 6112
rect 16120 6069 16129 6103
rect 16129 6069 16163 6103
rect 16163 6069 16172 6103
rect 16120 6060 16172 6069
rect 18052 6103 18104 6112
rect 18052 6069 18061 6103
rect 18061 6069 18095 6103
rect 18095 6069 18104 6103
rect 18052 6060 18104 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1768 5856 1820 5908
rect 2688 5856 2740 5908
rect 3700 5856 3752 5908
rect 4620 5899 4672 5908
rect 4620 5865 4629 5899
rect 4629 5865 4663 5899
rect 4663 5865 4672 5899
rect 4620 5856 4672 5865
rect 5540 5856 5592 5908
rect 6000 5856 6052 5908
rect 7380 5899 7432 5908
rect 7380 5865 7389 5899
rect 7389 5865 7423 5899
rect 7423 5865 7432 5899
rect 7380 5856 7432 5865
rect 8116 5856 8168 5908
rect 8760 5899 8812 5908
rect 8760 5865 8769 5899
rect 8769 5865 8803 5899
rect 8803 5865 8812 5899
rect 8760 5856 8812 5865
rect 9128 5899 9180 5908
rect 9128 5865 9137 5899
rect 9137 5865 9171 5899
rect 9171 5865 9180 5899
rect 9128 5856 9180 5865
rect 10048 5856 10100 5908
rect 11060 5856 11112 5908
rect 12440 5856 12492 5908
rect 12624 5856 12676 5908
rect 13084 5899 13136 5908
rect 13084 5865 13093 5899
rect 13093 5865 13127 5899
rect 13127 5865 13136 5899
rect 13084 5856 13136 5865
rect 13544 5856 13596 5908
rect 16120 5856 16172 5908
rect 11888 5788 11940 5840
rect 14556 5788 14608 5840
rect 3240 5720 3292 5772
rect 5448 5720 5500 5772
rect 6552 5720 6604 5772
rect 8208 5720 8260 5772
rect 9404 5720 9456 5772
rect 12256 5720 12308 5772
rect 12348 5720 12400 5772
rect 14188 5720 14240 5772
rect 16580 5763 16632 5772
rect 16580 5729 16614 5763
rect 16614 5729 16632 5763
rect 16580 5720 16632 5729
rect 18144 5720 18196 5772
rect 20628 5720 20680 5772
rect 2872 5695 2924 5704
rect 2872 5661 2881 5695
rect 2881 5661 2915 5695
rect 2915 5661 2924 5695
rect 2872 5652 2924 5661
rect 2320 5627 2372 5636
rect 2320 5593 2329 5627
rect 2329 5593 2363 5627
rect 2363 5593 2372 5627
rect 4436 5652 4488 5704
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 2320 5584 2372 5593
rect 8300 5584 8352 5636
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 11612 5652 11664 5704
rect 2044 5516 2096 5568
rect 2136 5516 2188 5568
rect 4160 5516 4212 5568
rect 10968 5584 11020 5636
rect 10784 5559 10836 5568
rect 10784 5525 10793 5559
rect 10793 5525 10827 5559
rect 10827 5525 10836 5559
rect 10784 5516 10836 5525
rect 14740 5652 14792 5704
rect 16212 5652 16264 5704
rect 15476 5516 15528 5568
rect 16488 5516 16540 5568
rect 18788 5516 18840 5568
rect 20996 5516 21048 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 4620 5355 4672 5364
rect 4620 5321 4629 5355
rect 4629 5321 4663 5355
rect 4663 5321 4672 5355
rect 4620 5312 4672 5321
rect 5356 5312 5408 5364
rect 6552 5312 6604 5364
rect 8760 5312 8812 5364
rect 11336 5312 11388 5364
rect 12256 5312 12308 5364
rect 13268 5312 13320 5364
rect 14004 5312 14056 5364
rect 14188 5312 14240 5364
rect 18144 5312 18196 5364
rect 11796 5287 11848 5296
rect 11796 5253 11805 5287
rect 11805 5253 11839 5287
rect 11839 5253 11848 5287
rect 11796 5244 11848 5253
rect 5540 5176 5592 5228
rect 7104 5176 7156 5228
rect 8484 5176 8536 5228
rect 1768 5108 1820 5160
rect 3240 5108 3292 5160
rect 3700 5151 3752 5160
rect 3700 5117 3709 5151
rect 3709 5117 3743 5151
rect 3743 5117 3752 5151
rect 3700 5108 3752 5117
rect 4988 5108 5040 5160
rect 6092 5108 6144 5160
rect 2044 5040 2096 5092
rect 3148 5040 3200 5092
rect 2136 4972 2188 5024
rect 3332 5015 3384 5024
rect 3332 4981 3341 5015
rect 3341 4981 3375 5015
rect 3375 4981 3384 5015
rect 3332 4972 3384 4981
rect 4436 4972 4488 5024
rect 5172 4972 5224 5024
rect 6092 4972 6144 5024
rect 7932 5108 7984 5160
rect 10784 5108 10836 5160
rect 12440 5176 12492 5228
rect 14096 5176 14148 5228
rect 16580 5176 16632 5228
rect 14004 5108 14056 5160
rect 6552 5040 6604 5092
rect 8116 5040 8168 5092
rect 6828 5015 6880 5024
rect 6828 4981 6837 5015
rect 6837 4981 6871 5015
rect 6871 4981 6880 5015
rect 6828 4972 6880 4981
rect 8300 4972 8352 5024
rect 9404 5015 9456 5024
rect 9404 4981 9413 5015
rect 9413 4981 9447 5015
rect 9447 4981 9456 5015
rect 9404 4972 9456 4981
rect 9772 5040 9824 5092
rect 13820 5040 13872 5092
rect 14464 5083 14516 5092
rect 14464 5049 14473 5083
rect 14473 5049 14507 5083
rect 14507 5049 14516 5083
rect 14464 5040 14516 5049
rect 16028 5040 16080 5092
rect 10140 4972 10192 5024
rect 10692 4972 10744 5024
rect 12900 5015 12952 5024
rect 12900 4981 12909 5015
rect 12909 4981 12943 5015
rect 12943 4981 12952 5015
rect 12900 4972 12952 4981
rect 14832 4972 14884 5024
rect 16120 5015 16172 5024
rect 16120 4981 16129 5015
rect 16129 4981 16163 5015
rect 16163 4981 16172 5015
rect 16120 4972 16172 4981
rect 16580 5015 16632 5024
rect 16580 4981 16589 5015
rect 16589 4981 16623 5015
rect 16623 4981 16632 5015
rect 16580 4972 16632 4981
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 19432 5108 19484 5160
rect 20536 5151 20588 5160
rect 20536 5117 20545 5151
rect 20545 5117 20579 5151
rect 20579 5117 20588 5151
rect 20536 5108 20588 5117
rect 18328 5083 18380 5092
rect 18328 5049 18337 5083
rect 18337 5049 18371 5083
rect 18371 5049 18380 5083
rect 18328 5040 18380 5049
rect 17408 4972 17460 5024
rect 19340 4972 19392 5024
rect 20628 4972 20680 5024
rect 22560 4972 22612 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 3148 4811 3200 4820
rect 3148 4777 3157 4811
rect 3157 4777 3191 4811
rect 3191 4777 3200 4811
rect 3148 4768 3200 4777
rect 4068 4768 4120 4820
rect 6736 4768 6788 4820
rect 8208 4768 8260 4820
rect 8760 4768 8812 4820
rect 11060 4768 11112 4820
rect 12808 4811 12860 4820
rect 12808 4777 12817 4811
rect 12817 4777 12851 4811
rect 12851 4777 12860 4811
rect 12808 4768 12860 4777
rect 13268 4768 13320 4820
rect 13452 4768 13504 4820
rect 14096 4811 14148 4820
rect 14096 4777 14105 4811
rect 14105 4777 14139 4811
rect 14139 4777 14148 4811
rect 14096 4768 14148 4777
rect 14464 4811 14516 4820
rect 14464 4777 14473 4811
rect 14473 4777 14507 4811
rect 14507 4777 14516 4811
rect 14464 4768 14516 4777
rect 17408 4811 17460 4820
rect 17408 4777 17417 4811
rect 17417 4777 17451 4811
rect 17451 4777 17460 4811
rect 17408 4768 17460 4777
rect 2320 4700 2372 4752
rect 5540 4700 5592 4752
rect 12716 4700 12768 4752
rect 14648 4700 14700 4752
rect 18420 4700 18472 4752
rect 4712 4632 4764 4684
rect 8576 4632 8628 4684
rect 9404 4632 9456 4684
rect 1768 4607 1820 4616
rect 1768 4573 1777 4607
rect 1777 4573 1811 4607
rect 1811 4573 1820 4607
rect 1768 4564 1820 4573
rect 4620 4564 4672 4616
rect 4804 4564 4856 4616
rect 5448 4564 5500 4616
rect 8300 4564 8352 4616
rect 8668 4607 8720 4616
rect 8668 4573 8677 4607
rect 8677 4573 8711 4607
rect 8711 4573 8720 4607
rect 8668 4564 8720 4573
rect 10140 4607 10192 4616
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 13452 4632 13504 4684
rect 16304 4675 16356 4684
rect 16304 4641 16338 4675
rect 16338 4641 16356 4675
rect 16304 4632 16356 4641
rect 18236 4675 18288 4684
rect 18236 4641 18245 4675
rect 18245 4641 18279 4675
rect 18279 4641 18288 4675
rect 18236 4632 18288 4641
rect 19524 4675 19576 4684
rect 19524 4641 19533 4675
rect 19533 4641 19567 4675
rect 19567 4641 19576 4675
rect 19524 4632 19576 4641
rect 20904 4675 20956 4684
rect 20904 4641 20913 4675
rect 20913 4641 20947 4675
rect 20947 4641 20956 4675
rect 20904 4632 20956 4641
rect 11888 4607 11940 4616
rect 11888 4573 11897 4607
rect 11897 4573 11931 4607
rect 11931 4573 11940 4607
rect 11888 4564 11940 4573
rect 12992 4564 13044 4616
rect 1676 4471 1728 4480
rect 1676 4437 1685 4471
rect 1685 4437 1719 4471
rect 1719 4437 1728 4471
rect 5172 4471 5224 4480
rect 1676 4428 1728 4437
rect 5172 4437 5181 4471
rect 5181 4437 5215 4471
rect 5215 4437 5224 4471
rect 5172 4428 5224 4437
rect 7104 4428 7156 4480
rect 7288 4428 7340 4480
rect 9404 4471 9456 4480
rect 9404 4437 9413 4471
rect 9413 4437 9447 4471
rect 9447 4437 9456 4471
rect 9404 4428 9456 4437
rect 10784 4471 10836 4480
rect 10784 4437 10793 4471
rect 10793 4437 10827 4471
rect 10827 4437 10836 4471
rect 10784 4428 10836 4437
rect 11244 4471 11296 4480
rect 11244 4437 11253 4471
rect 11253 4437 11287 4471
rect 11287 4437 11296 4471
rect 11244 4428 11296 4437
rect 12440 4471 12492 4480
rect 12440 4437 12449 4471
rect 12449 4437 12483 4471
rect 12483 4437 12492 4471
rect 12440 4428 12492 4437
rect 15476 4471 15528 4480
rect 15476 4437 15485 4471
rect 15485 4437 15519 4471
rect 15519 4437 15528 4471
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 22192 4564 22244 4616
rect 15476 4428 15528 4437
rect 21548 4428 21600 4480
rect 22100 4428 22152 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1584 4267 1636 4276
rect 1584 4233 1593 4267
rect 1593 4233 1627 4267
rect 1627 4233 1636 4267
rect 1584 4224 1636 4233
rect 2320 4224 2372 4276
rect 3332 4224 3384 4276
rect 4804 4224 4856 4276
rect 5448 4224 5500 4276
rect 7932 4267 7984 4276
rect 7932 4233 7941 4267
rect 7941 4233 7975 4267
rect 7975 4233 7984 4267
rect 7932 4224 7984 4233
rect 9404 4224 9456 4276
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 4712 4088 4764 4140
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 9404 4088 9456 4140
rect 10784 4224 10836 4276
rect 15660 4224 15712 4276
rect 18236 4224 18288 4276
rect 19524 4267 19576 4276
rect 19524 4233 19533 4267
rect 19533 4233 19567 4267
rect 19567 4233 19576 4267
rect 19524 4224 19576 4233
rect 12532 4088 12584 4140
rect 17408 4131 17460 4140
rect 17408 4097 17417 4131
rect 17417 4097 17451 4131
rect 17451 4097 17460 4131
rect 17408 4088 17460 4097
rect 20904 4224 20956 4276
rect 22192 4088 22244 4140
rect 4804 4020 4856 4072
rect 6000 4063 6052 4072
rect 6000 4029 6009 4063
rect 6009 4029 6043 4063
rect 6043 4029 6052 4063
rect 6000 4020 6052 4029
rect 6828 4020 6880 4072
rect 7932 4020 7984 4072
rect 1216 3952 1268 4004
rect 1676 3952 1728 4004
rect 3332 3952 3384 4004
rect 4344 3952 4396 4004
rect 5172 3995 5224 4004
rect 5172 3961 5181 3995
rect 5181 3961 5215 3995
rect 5215 3961 5224 3995
rect 5172 3952 5224 3961
rect 8116 3952 8168 4004
rect 4620 3884 4672 3936
rect 5448 3884 5500 3936
rect 6736 3884 6788 3936
rect 9036 3952 9088 4004
rect 10232 3952 10284 4004
rect 10692 4020 10744 4072
rect 11336 3952 11388 4004
rect 11888 3952 11940 4004
rect 12440 4020 12492 4072
rect 15476 4020 15528 4072
rect 19524 4020 19576 4072
rect 20904 4063 20956 4072
rect 20904 4029 20913 4063
rect 20913 4029 20947 4063
rect 20947 4029 20956 4063
rect 20904 4020 20956 4029
rect 13820 3952 13872 4004
rect 15108 3952 15160 4004
rect 9128 3884 9180 3936
rect 9404 3884 9456 3936
rect 11520 3927 11572 3936
rect 11520 3893 11529 3927
rect 11529 3893 11563 3927
rect 11563 3893 11572 3927
rect 11520 3884 11572 3893
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 13452 3927 13504 3936
rect 12440 3884 12492 3893
rect 13452 3893 13461 3927
rect 13461 3893 13495 3927
rect 13495 3893 13504 3927
rect 13452 3884 13504 3893
rect 15292 3927 15344 3936
rect 15292 3893 15301 3927
rect 15301 3893 15335 3927
rect 15335 3893 15344 3927
rect 15292 3884 15344 3893
rect 16304 3884 16356 3936
rect 16672 3884 16724 3936
rect 18144 3952 18196 4004
rect 18420 3995 18472 4004
rect 18420 3961 18429 3995
rect 18429 3961 18463 3995
rect 18463 3961 18472 3995
rect 18420 3952 18472 3961
rect 18328 3884 18380 3936
rect 19984 3884 20036 3936
rect 21824 3927 21876 3936
rect 21824 3893 21833 3927
rect 21833 3893 21867 3927
rect 21867 3893 21876 3927
rect 21824 3884 21876 3893
rect 23204 3952 23256 4004
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 204 3680 256 3732
rect 2044 3680 2096 3732
rect 2320 3680 2372 3732
rect 4712 3723 4764 3732
rect 4712 3689 4721 3723
rect 4721 3689 4755 3723
rect 4755 3689 4764 3723
rect 4712 3680 4764 3689
rect 5172 3680 5224 3732
rect 7288 3680 7340 3732
rect 8116 3723 8168 3732
rect 8116 3689 8125 3723
rect 8125 3689 8159 3723
rect 8159 3689 8168 3723
rect 8116 3680 8168 3689
rect 8300 3680 8352 3732
rect 8576 3680 8628 3732
rect 10140 3680 10192 3732
rect 10692 3723 10744 3732
rect 10692 3689 10701 3723
rect 10701 3689 10735 3723
rect 10735 3689 10744 3723
rect 10692 3680 10744 3689
rect 11060 3723 11112 3732
rect 11060 3689 11069 3723
rect 11069 3689 11103 3723
rect 11103 3689 11112 3723
rect 11060 3680 11112 3689
rect 12532 3723 12584 3732
rect 12532 3689 12541 3723
rect 12541 3689 12575 3723
rect 12575 3689 12584 3723
rect 12532 3680 12584 3689
rect 12716 3680 12768 3732
rect 12992 3680 13044 3732
rect 13728 3680 13780 3732
rect 16028 3680 16080 3732
rect 16212 3680 16264 3732
rect 16580 3680 16632 3732
rect 17868 3723 17920 3732
rect 17868 3689 17877 3723
rect 17877 3689 17911 3723
rect 17911 3689 17920 3723
rect 17868 3680 17920 3689
rect 18328 3680 18380 3732
rect 1768 3587 1820 3596
rect 1768 3553 1777 3587
rect 1777 3553 1811 3587
rect 1811 3553 1820 3587
rect 1768 3544 1820 3553
rect 2044 3587 2096 3596
rect 2044 3553 2078 3587
rect 2078 3553 2096 3587
rect 2044 3544 2096 3553
rect 6828 3612 6880 3664
rect 7012 3612 7064 3664
rect 11520 3612 11572 3664
rect 14740 3612 14792 3664
rect 16396 3655 16448 3664
rect 16396 3621 16405 3655
rect 16405 3621 16439 3655
rect 16439 3621 16448 3655
rect 16396 3612 16448 3621
rect 19432 3612 19484 3664
rect 6736 3544 6788 3596
rect 7196 3587 7248 3596
rect 7196 3553 7205 3587
rect 7205 3553 7239 3587
rect 7239 3553 7248 3587
rect 7196 3544 7248 3553
rect 9772 3544 9824 3596
rect 10784 3544 10836 3596
rect 12348 3544 12400 3596
rect 12624 3544 12676 3596
rect 14464 3544 14516 3596
rect 19064 3587 19116 3596
rect 19064 3553 19073 3587
rect 19073 3553 19107 3587
rect 19107 3553 19116 3587
rect 19064 3544 19116 3553
rect 20904 3587 20956 3596
rect 20904 3553 20913 3587
rect 20913 3553 20947 3587
rect 20947 3553 20956 3587
rect 20904 3544 20956 3553
rect 22008 3587 22060 3596
rect 22008 3553 22017 3587
rect 22017 3553 22051 3587
rect 22051 3553 22060 3587
rect 22008 3544 22060 3553
rect 23940 3587 23992 3596
rect 23940 3553 23949 3587
rect 23949 3553 23983 3587
rect 23983 3553 23992 3587
rect 23940 3544 23992 3553
rect 3332 3476 3384 3528
rect 5448 3476 5500 3528
rect 7104 3408 7156 3460
rect 9588 3476 9640 3528
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 16672 3476 16724 3528
rect 17776 3476 17828 3528
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 16948 3451 17000 3460
rect 16948 3417 16957 3451
rect 16957 3417 16991 3451
rect 16991 3417 17000 3451
rect 16948 3408 17000 3417
rect 3516 3340 3568 3392
rect 4436 3340 4488 3392
rect 4804 3340 4856 3392
rect 5172 3383 5224 3392
rect 5172 3349 5181 3383
rect 5181 3349 5215 3383
rect 5215 3349 5224 3383
rect 5172 3340 5224 3349
rect 7472 3340 7524 3392
rect 8668 3340 8720 3392
rect 9404 3340 9456 3392
rect 9956 3340 10008 3392
rect 13636 3340 13688 3392
rect 14188 3340 14240 3392
rect 15476 3383 15528 3392
rect 15476 3349 15485 3383
rect 15485 3349 15519 3383
rect 15519 3349 15528 3383
rect 15476 3340 15528 3349
rect 18604 3383 18656 3392
rect 18604 3349 18613 3383
rect 18613 3349 18647 3383
rect 18647 3349 18656 3383
rect 18604 3340 18656 3349
rect 21088 3383 21140 3392
rect 21088 3349 21097 3383
rect 21097 3349 21131 3383
rect 21131 3349 21140 3383
rect 21088 3340 21140 3349
rect 22192 3383 22244 3392
rect 22192 3349 22201 3383
rect 22201 3349 22235 3383
rect 22235 3349 22244 3383
rect 22192 3340 22244 3349
rect 24124 3383 24176 3392
rect 24124 3349 24133 3383
rect 24133 3349 24167 3383
rect 24167 3349 24176 3383
rect 24124 3340 24176 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1492 3136 1544 3188
rect 2228 3136 2280 3188
rect 4344 3136 4396 3188
rect 5448 3136 5500 3188
rect 7196 3136 7248 3188
rect 10232 3136 10284 3188
rect 1952 3000 2004 3052
rect 3516 3000 3568 3052
rect 2228 2932 2280 2984
rect 3332 2975 3384 2984
rect 3332 2941 3341 2975
rect 3341 2941 3375 2975
rect 3375 2941 3384 2975
rect 3332 2932 3384 2941
rect 4068 2932 4120 2984
rect 4436 3000 4488 3052
rect 8208 3068 8260 3120
rect 9404 3068 9456 3120
rect 9956 3111 10008 3120
rect 9956 3077 9965 3111
rect 9965 3077 9999 3111
rect 9999 3077 10008 3111
rect 11520 3111 11572 3120
rect 9956 3068 10008 3077
rect 11520 3077 11529 3111
rect 11529 3077 11563 3111
rect 11563 3077 11572 3111
rect 11520 3068 11572 3077
rect 10876 3043 10928 3052
rect 4620 2932 4672 2984
rect 7104 2932 7156 2984
rect 7472 2932 7524 2984
rect 10876 3009 10885 3043
rect 10885 3009 10919 3043
rect 10919 3009 10928 3043
rect 10876 3000 10928 3009
rect 10968 3043 11020 3052
rect 10968 3009 10977 3043
rect 10977 3009 11011 3043
rect 11011 3009 11020 3043
rect 10968 3000 11020 3009
rect 4712 2864 4764 2916
rect 5724 2864 5776 2916
rect 9036 2932 9088 2984
rect 11428 2932 11480 2984
rect 12440 3136 12492 3188
rect 13728 3136 13780 3188
rect 14464 3179 14516 3188
rect 14464 3145 14473 3179
rect 14473 3145 14507 3179
rect 14507 3145 14516 3179
rect 14464 3136 14516 3145
rect 16212 3136 16264 3188
rect 17868 3136 17920 3188
rect 18052 3179 18104 3188
rect 18052 3145 18061 3179
rect 18061 3145 18095 3179
rect 18095 3145 18104 3179
rect 18052 3136 18104 3145
rect 18144 3136 18196 3188
rect 21364 3179 21416 3188
rect 21364 3145 21373 3179
rect 21373 3145 21407 3179
rect 21407 3145 21416 3179
rect 21364 3136 21416 3145
rect 22008 3136 22060 3188
rect 24768 3179 24820 3188
rect 24768 3145 24777 3179
rect 24777 3145 24811 3179
rect 24811 3145 24820 3179
rect 24768 3136 24820 3145
rect 16120 3068 16172 3120
rect 16396 3043 16448 3052
rect 16396 3009 16405 3043
rect 16405 3009 16439 3043
rect 16439 3009 16448 3043
rect 16396 3000 16448 3009
rect 18328 3000 18380 3052
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 19064 3000 19116 3052
rect 21824 3000 21876 3052
rect 12348 2932 12400 2984
rect 8760 2864 8812 2916
rect 12532 2932 12584 2984
rect 15476 2932 15528 2984
rect 16948 2932 17000 2984
rect 20260 2975 20312 2984
rect 20260 2941 20269 2975
rect 20269 2941 20303 2975
rect 20303 2941 20312 2975
rect 20260 2932 20312 2941
rect 21364 2932 21416 2984
rect 14188 2864 14240 2916
rect 25228 2907 25280 2916
rect 25228 2873 25237 2907
rect 25237 2873 25271 2907
rect 25271 2873 25280 2907
rect 25228 2864 25280 2873
rect 7012 2839 7064 2848
rect 7012 2805 7021 2839
rect 7021 2805 7055 2839
rect 7055 2805 7064 2839
rect 7012 2796 7064 2805
rect 10140 2796 10192 2848
rect 13820 2839 13872 2848
rect 13820 2805 13829 2839
rect 13829 2805 13863 2839
rect 13863 2805 13872 2839
rect 13820 2796 13872 2805
rect 16028 2839 16080 2848
rect 16028 2805 16037 2839
rect 16037 2805 16071 2839
rect 16071 2805 16080 2839
rect 16028 2796 16080 2805
rect 18144 2796 18196 2848
rect 21732 2839 21784 2848
rect 21732 2805 21741 2839
rect 21741 2805 21775 2839
rect 21775 2805 21784 2839
rect 21732 2796 21784 2805
rect 23940 2839 23992 2848
rect 23940 2805 23949 2839
rect 23949 2805 23983 2839
rect 23983 2805 23992 2839
rect 23940 2796 23992 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1952 2592 2004 2644
rect 2504 2592 2556 2644
rect 3240 2635 3292 2644
rect 3240 2601 3249 2635
rect 3249 2601 3283 2635
rect 3283 2601 3292 2635
rect 3240 2592 3292 2601
rect 5724 2635 5776 2644
rect 5724 2601 5733 2635
rect 5733 2601 5767 2635
rect 5767 2601 5776 2635
rect 5724 2592 5776 2601
rect 6000 2635 6052 2644
rect 6000 2601 6009 2635
rect 6009 2601 6043 2635
rect 6043 2601 6052 2635
rect 6000 2592 6052 2601
rect 9036 2592 9088 2644
rect 10876 2592 10928 2644
rect 11428 2635 11480 2644
rect 11428 2601 11437 2635
rect 11437 2601 11471 2635
rect 11471 2601 11480 2635
rect 11428 2592 11480 2601
rect 14188 2635 14240 2644
rect 4620 2567 4672 2576
rect 4620 2533 4632 2567
rect 4632 2533 4672 2567
rect 4620 2524 4672 2533
rect 8668 2524 8720 2576
rect 9680 2524 9732 2576
rect 14188 2601 14197 2635
rect 14197 2601 14231 2635
rect 14231 2601 14240 2635
rect 14188 2592 14240 2601
rect 15844 2635 15896 2644
rect 15844 2601 15853 2635
rect 15853 2601 15887 2635
rect 15887 2601 15896 2635
rect 15844 2592 15896 2601
rect 16672 2592 16724 2644
rect 17776 2592 17828 2644
rect 18144 2635 18196 2644
rect 18144 2601 18153 2635
rect 18153 2601 18187 2635
rect 18187 2601 18196 2635
rect 18144 2592 18196 2601
rect 20904 2635 20956 2644
rect 20904 2601 20913 2635
rect 20913 2601 20947 2635
rect 20947 2601 20956 2635
rect 20904 2592 20956 2601
rect 24768 2635 24820 2644
rect 24768 2601 24777 2635
rect 24777 2601 24811 2635
rect 24811 2601 24820 2635
rect 24768 2592 24820 2601
rect 1400 2456 1452 2508
rect 2964 2456 3016 2508
rect 4436 2456 4488 2508
rect 7472 2499 7524 2508
rect 7472 2465 7481 2499
rect 7481 2465 7515 2499
rect 7515 2465 7524 2499
rect 7472 2456 7524 2465
rect 9956 2456 10008 2508
rect 3240 2388 3292 2440
rect 6368 2431 6420 2440
rect 6368 2397 6377 2431
rect 6377 2397 6411 2431
rect 6411 2397 6420 2431
rect 6368 2388 6420 2397
rect 9588 2431 9640 2440
rect 9588 2397 9597 2431
rect 9597 2397 9631 2431
rect 9631 2397 9640 2431
rect 9588 2388 9640 2397
rect 13820 2524 13872 2576
rect 12440 2456 12492 2508
rect 13636 2456 13688 2508
rect 20720 2524 20772 2576
rect 18328 2499 18380 2508
rect 18328 2465 18337 2499
rect 18337 2465 18371 2499
rect 18371 2465 18380 2499
rect 18328 2456 18380 2465
rect 19616 2499 19668 2508
rect 19616 2465 19625 2499
rect 19625 2465 19659 2499
rect 19659 2465 19668 2499
rect 19616 2456 19668 2465
rect 21180 2499 21232 2508
rect 21180 2465 21189 2499
rect 21189 2465 21223 2499
rect 21223 2465 21232 2499
rect 21180 2456 21232 2465
rect 22468 2499 22520 2508
rect 22468 2465 22477 2499
rect 22477 2465 22511 2499
rect 22511 2465 22520 2499
rect 22468 2456 22520 2465
rect 15292 2388 15344 2440
rect 16028 2431 16080 2440
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 2136 2363 2188 2372
rect 2136 2329 2145 2363
rect 2145 2329 2179 2363
rect 2179 2329 2188 2363
rect 2136 2320 2188 2329
rect 10692 2320 10744 2372
rect 15476 2363 15528 2372
rect 15476 2329 15485 2363
rect 15485 2329 15519 2363
rect 15519 2329 15528 2363
rect 15476 2320 15528 2329
rect 15568 2320 15620 2372
rect 2044 2295 2096 2304
rect 2044 2261 2053 2295
rect 2053 2261 2087 2295
rect 2087 2261 2096 2295
rect 2044 2252 2096 2261
rect 9404 2252 9456 2304
rect 10968 2295 11020 2304
rect 10968 2261 10977 2295
rect 10977 2261 11011 2295
rect 11011 2261 11020 2295
rect 10968 2252 11020 2261
rect 22652 2295 22704 2304
rect 22652 2261 22661 2295
rect 22661 2261 22695 2295
rect 22695 2261 22704 2295
rect 22652 2252 22704 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 5632 1980 5684 2032
rect 6276 1980 6328 2032
rect 14280 1980 14332 2032
rect 14924 1980 14976 2032
rect 23480 1980 23532 2032
rect 24308 1980 24360 2032
rect 9864 1368 9916 1420
rect 10600 1368 10652 1420
rect 11612 552 11664 604
rect 11704 552 11756 604
rect 23572 552 23624 604
rect 23756 552 23808 604
rect 24952 552 25004 604
rect 25412 552 25464 604
<< metal2 >>
rect 2410 27704 2466 27713
rect 2410 27639 2466 27648
rect 1582 24848 1638 24857
rect 1582 24783 1638 24792
rect 1596 24410 1624 24783
rect 1584 24404 1636 24410
rect 1584 24346 1636 24352
rect 1400 24268 1452 24274
rect 1400 24210 1452 24216
rect 1412 23866 1440 24210
rect 1400 23860 1452 23866
rect 1400 23802 1452 23808
rect 1860 23860 1912 23866
rect 1860 23802 1912 23808
rect 1584 23520 1636 23526
rect 1584 23462 1636 23468
rect 1596 21457 1624 23462
rect 1872 22642 1900 23802
rect 1952 23656 2004 23662
rect 1952 23598 2004 23604
rect 1964 23254 1992 23598
rect 1952 23248 2004 23254
rect 1952 23190 2004 23196
rect 1860 22636 1912 22642
rect 1860 22578 1912 22584
rect 2044 22092 2096 22098
rect 2044 22034 2096 22040
rect 2056 21894 2084 22034
rect 2136 22024 2188 22030
rect 2136 21966 2188 21972
rect 2044 21888 2096 21894
rect 2044 21830 2096 21836
rect 1582 21448 1638 21457
rect 1582 21383 1638 21392
rect 1950 21448 2006 21457
rect 1950 21383 2006 21392
rect 1964 21078 1992 21383
rect 1952 21072 2004 21078
rect 1952 21014 2004 21020
rect 1676 21004 1728 21010
rect 1676 20946 1728 20952
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1412 19514 1440 19858
rect 1688 19718 1716 20946
rect 1950 20496 2006 20505
rect 1950 20431 1952 20440
rect 2004 20431 2006 20440
rect 1952 20402 2004 20408
rect 1768 20392 1820 20398
rect 1768 20334 1820 20340
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1400 19508 1452 19514
rect 1400 19450 1452 19456
rect 1412 18465 1440 19450
rect 1504 19378 1532 19417
rect 1492 19372 1544 19378
rect 1492 19314 1544 19320
rect 1398 18456 1454 18465
rect 1398 18391 1454 18400
rect 1504 17610 1532 19314
rect 1584 19304 1636 19310
rect 1582 19272 1584 19281
rect 1636 19272 1638 19281
rect 1582 19207 1638 19216
rect 1582 18320 1638 18329
rect 1582 18255 1638 18264
rect 1492 17604 1544 17610
rect 1492 17546 1544 17552
rect 1400 17536 1452 17542
rect 1400 17478 1452 17484
rect 1412 14618 1440 17478
rect 1596 17134 1624 18255
rect 1674 18184 1730 18193
rect 1674 18119 1730 18128
rect 1584 17128 1636 17134
rect 1584 17070 1636 17076
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 1504 16046 1532 16390
rect 1492 16040 1544 16046
rect 1490 16008 1492 16017
rect 1544 16008 1546 16017
rect 1490 15943 1546 15952
rect 1400 14612 1452 14618
rect 1400 14554 1452 14560
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1306 12336 1362 12345
rect 1306 12271 1362 12280
rect 1320 11014 1348 12271
rect 1308 11008 1360 11014
rect 1308 10950 1360 10956
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1412 9586 1440 10542
rect 1504 10198 1532 12582
rect 1492 10192 1544 10198
rect 1492 10134 1544 10140
rect 1490 9752 1546 9761
rect 1490 9687 1546 9696
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1400 6656 1452 6662
rect 1400 6598 1452 6604
rect 1216 4004 1268 4010
rect 1216 3946 1268 3952
rect 204 3732 256 3738
rect 204 3674 256 3680
rect 216 480 244 3674
rect 662 2816 718 2825
rect 662 2751 718 2760
rect 676 480 704 2751
rect 1228 480 1256 3946
rect 1412 2514 1440 6598
rect 1504 3194 1532 9687
rect 1596 9178 1624 17070
rect 1688 16114 1716 18119
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1780 15706 1808 20334
rect 2056 19310 2084 21830
rect 2148 21486 2176 21966
rect 2228 21956 2280 21962
rect 2228 21898 2280 21904
rect 2136 21480 2188 21486
rect 2136 21422 2188 21428
rect 2148 20097 2176 21422
rect 2134 20088 2190 20097
rect 2134 20023 2190 20032
rect 2136 19712 2188 19718
rect 2136 19654 2188 19660
rect 2148 19417 2176 19654
rect 2134 19408 2190 19417
rect 2134 19343 2190 19352
rect 2044 19304 2096 19310
rect 2044 19246 2096 19252
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 2044 18828 2096 18834
rect 2044 18770 2096 18776
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 1964 16794 1992 18566
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 1964 15026 1992 15302
rect 2056 15162 2084 18770
rect 2148 18170 2176 19110
rect 2240 18601 2268 21898
rect 2320 20324 2372 20330
rect 2320 20266 2372 20272
rect 2332 18834 2360 20266
rect 2424 20262 2452 27639
rect 7010 27520 7066 28000
rect 20994 27520 21050 28000
rect 4066 27160 4122 27169
rect 4122 27118 4200 27146
rect 4066 27095 4122 27104
rect 4066 26616 4122 26625
rect 4066 26551 4068 26560
rect 4120 26551 4122 26560
rect 4068 26522 4120 26528
rect 3790 26072 3846 26081
rect 3790 26007 3846 26016
rect 2686 25392 2742 25401
rect 2686 25327 2742 25336
rect 2700 23866 2728 25327
rect 3804 23866 3832 26007
rect 4066 24304 4122 24313
rect 4066 24239 4122 24248
rect 2688 23860 2740 23866
rect 2688 23802 2740 23808
rect 3792 23860 3844 23866
rect 3792 23802 3844 23808
rect 2596 23520 2648 23526
rect 2596 23462 2648 23468
rect 2504 22432 2556 22438
rect 2502 22400 2504 22409
rect 2556 22400 2558 22409
rect 2502 22335 2558 22344
rect 2504 22092 2556 22098
rect 2504 22034 2556 22040
rect 2516 21350 2544 22034
rect 2504 21344 2556 21350
rect 2504 21286 2556 21292
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 2412 19712 2464 19718
rect 2412 19654 2464 19660
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2424 18766 2452 19654
rect 2516 19242 2544 21286
rect 2608 20466 2636 23462
rect 4080 23361 4108 24239
rect 4066 23352 4122 23361
rect 4066 23287 4122 23296
rect 2872 23180 2924 23186
rect 2872 23122 2924 23128
rect 2780 22568 2832 22574
rect 2700 22516 2780 22522
rect 2700 22510 2832 22516
rect 2700 22494 2820 22510
rect 2700 21554 2728 22494
rect 2884 22438 2912 23122
rect 4172 22778 4200 27118
rect 5540 26580 5592 26586
rect 5540 26522 5592 26528
rect 4436 23520 4488 23526
rect 4436 23462 4488 23468
rect 4160 22772 4212 22778
rect 4160 22714 4212 22720
rect 4250 22536 4306 22545
rect 4250 22471 4306 22480
rect 2872 22432 2924 22438
rect 2872 22374 2924 22380
rect 3148 22432 3200 22438
rect 3148 22374 3200 22380
rect 2884 22137 2912 22374
rect 2870 22128 2926 22137
rect 2870 22063 2926 22072
rect 3160 22001 3188 22374
rect 4068 22092 4120 22098
rect 4068 22034 4120 22040
rect 3146 21992 3202 22001
rect 3146 21927 3202 21936
rect 2872 21888 2924 21894
rect 2872 21830 2924 21836
rect 2688 21548 2740 21554
rect 2688 21490 2740 21496
rect 2780 21480 2832 21486
rect 2700 21428 2780 21434
rect 2700 21422 2832 21428
rect 2700 21406 2820 21422
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 2596 20256 2648 20262
rect 2596 20198 2648 20204
rect 2504 19236 2556 19242
rect 2504 19178 2556 19184
rect 2608 19174 2636 20198
rect 2700 20058 2728 21406
rect 2688 20052 2740 20058
rect 2688 19994 2740 20000
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 2700 19378 2728 19858
rect 2884 19689 2912 21830
rect 4080 21690 4108 22034
rect 4264 21962 4292 22471
rect 4252 21956 4304 21962
rect 4252 21898 4304 21904
rect 4068 21684 4120 21690
rect 4068 21626 4120 21632
rect 3976 21480 4028 21486
rect 3976 21422 4028 21428
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 2870 19680 2926 19689
rect 2870 19615 2926 19624
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 2884 19009 2912 19246
rect 3068 19145 3096 21286
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 3516 19712 3568 19718
rect 3516 19654 3568 19660
rect 3528 19281 3556 19654
rect 3514 19272 3570 19281
rect 3514 19207 3570 19216
rect 3054 19136 3110 19145
rect 3054 19071 3110 19080
rect 2594 19000 2650 19009
rect 2594 18935 2650 18944
rect 2870 19000 2926 19009
rect 2870 18935 2926 18944
rect 2412 18760 2464 18766
rect 2412 18702 2464 18708
rect 2504 18760 2556 18766
rect 2504 18702 2556 18708
rect 2226 18592 2282 18601
rect 2226 18527 2282 18536
rect 2148 18142 2268 18170
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 2148 16658 2176 18022
rect 2240 16674 2268 18142
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 2332 17542 2360 18022
rect 2320 17536 2372 17542
rect 2320 17478 2372 17484
rect 2136 16652 2188 16658
rect 2240 16646 2360 16674
rect 2136 16594 2188 16600
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2240 16250 2268 16526
rect 2228 16244 2280 16250
rect 2228 16186 2280 16192
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1780 13394 1808 13670
rect 1964 13462 1992 14962
rect 1952 13456 2004 13462
rect 1952 13398 2004 13404
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1768 13184 1820 13190
rect 1820 13144 1900 13172
rect 1768 13126 1820 13132
rect 1872 12782 1900 13144
rect 2332 12986 2360 16646
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1674 12472 1730 12481
rect 1674 12407 1730 12416
rect 1688 11762 1716 12407
rect 1872 12186 1900 12718
rect 2332 12646 2360 12922
rect 2320 12640 2372 12646
rect 2320 12582 2372 12588
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 1872 12158 2176 12186
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1780 10470 1808 11154
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1780 10266 1808 10406
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1780 9722 1808 10202
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1780 8974 1808 9658
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1872 8498 1900 9522
rect 1964 9042 1992 12038
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 2056 9178 2084 9862
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 1950 8800 2006 8809
rect 1950 8735 2006 8744
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1872 8022 1900 8434
rect 1860 8016 1912 8022
rect 1860 7958 1912 7964
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1596 6118 1624 6734
rect 1780 6458 1808 6802
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1676 6180 1728 6186
rect 1676 6122 1728 6128
rect 1584 6112 1636 6118
rect 1582 6080 1584 6089
rect 1636 6080 1638 6089
rect 1582 6015 1638 6024
rect 1688 5930 1716 6122
rect 1596 5902 1716 5930
rect 1780 5914 1808 6394
rect 1768 5908 1820 5914
rect 1596 4282 1624 5902
rect 1768 5850 1820 5856
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 1780 4622 1808 5102
rect 1858 4720 1914 4729
rect 1858 4655 1914 4664
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1676 4480 1728 4486
rect 1676 4422 1728 4428
rect 1584 4276 1636 4282
rect 1584 4218 1636 4224
rect 1688 4010 1716 4422
rect 1676 4004 1728 4010
rect 1676 3946 1728 3952
rect 1780 3602 1808 4558
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1872 3482 1900 4655
rect 1964 3777 1992 8735
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 2056 5574 2084 6258
rect 2148 5681 2176 12158
rect 2332 11558 2360 12242
rect 2424 11898 2452 18702
rect 2516 18290 2544 18702
rect 2504 18284 2556 18290
rect 2504 18226 2556 18232
rect 2504 18080 2556 18086
rect 2504 18022 2556 18028
rect 2516 17785 2544 18022
rect 2502 17776 2558 17785
rect 2502 17711 2558 17720
rect 2516 17241 2544 17711
rect 2502 17232 2558 17241
rect 2502 17167 2558 17176
rect 2504 17128 2556 17134
rect 2504 17070 2556 17076
rect 2516 13394 2544 17070
rect 2608 14618 2636 18935
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2976 18329 3004 18566
rect 2962 18320 3018 18329
rect 2962 18255 3018 18264
rect 2780 18148 2832 18154
rect 2780 18090 2832 18096
rect 2792 18034 2820 18090
rect 2700 18006 2820 18034
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 2700 17882 2728 18006
rect 2688 17876 2740 17882
rect 2688 17818 2740 17824
rect 2780 17740 2832 17746
rect 2780 17682 2832 17688
rect 2792 16998 2820 17682
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 2780 16992 2832 16998
rect 2780 16934 2832 16940
rect 2884 16794 2912 17614
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2700 16674 2728 16730
rect 2976 16726 3004 17614
rect 3056 17060 3108 17066
rect 3056 17002 3108 17008
rect 3068 16726 3096 17002
rect 2964 16720 3016 16726
rect 2700 16646 2820 16674
rect 2964 16662 3016 16668
rect 3056 16720 3108 16726
rect 3056 16662 3108 16668
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2700 15314 2728 16186
rect 2792 15706 2820 16646
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 2964 15972 3016 15978
rect 2964 15914 3016 15920
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2976 15638 3004 15914
rect 2964 15632 3016 15638
rect 2964 15574 3016 15580
rect 2976 15502 3004 15574
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2700 15286 2912 15314
rect 2686 15056 2742 15065
rect 2686 14991 2742 15000
rect 2700 14958 2728 14991
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2700 14550 2728 14894
rect 2688 14544 2740 14550
rect 2688 14486 2740 14492
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 13870 2820 14418
rect 2884 14074 2912 15286
rect 3068 15162 3096 15506
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 3160 14618 3188 16594
rect 3238 16280 3294 16289
rect 3238 16215 3294 16224
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3252 14498 3280 16215
rect 3160 14470 3280 14498
rect 3344 14482 3372 18022
rect 3528 15162 3556 19207
rect 3620 18426 3648 20198
rect 3988 19990 4016 21422
rect 4160 21344 4212 21350
rect 4160 21286 4212 21292
rect 4172 20913 4200 21286
rect 4448 21078 4476 23462
rect 5262 23216 5318 23225
rect 5262 23151 5318 23160
rect 4712 22432 4764 22438
rect 4712 22374 4764 22380
rect 4724 22273 4752 22374
rect 4710 22264 4766 22273
rect 4710 22199 4766 22208
rect 5276 21690 5304 23151
rect 5552 21962 5580 26522
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 7024 24177 7052 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 7010 24168 7066 24177
rect 7010 24103 7066 24112
rect 20166 24168 20222 24177
rect 20166 24103 20222 24112
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 7470 23760 7526 23769
rect 7470 23695 7526 23704
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 7484 22778 7512 23695
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 8298 23352 8354 23361
rect 10289 23344 10585 23364
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 8298 23287 8300 23296
rect 8352 23287 8354 23296
rect 8300 23258 8352 23264
rect 8116 23180 8168 23186
rect 8116 23122 8168 23128
rect 8128 22778 8156 23122
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 7472 22772 7524 22778
rect 7472 22714 7524 22720
rect 8116 22772 8168 22778
rect 8116 22714 8168 22720
rect 8116 22432 8168 22438
rect 8116 22374 8168 22380
rect 9588 22432 9640 22438
rect 9588 22374 9640 22380
rect 9954 22400 10010 22409
rect 6000 22092 6052 22098
rect 6000 22034 6052 22040
rect 7840 22092 7892 22098
rect 7840 22034 7892 22040
rect 5540 21956 5592 21962
rect 5540 21898 5592 21904
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6012 21690 6040 22034
rect 4528 21684 4580 21690
rect 4528 21626 4580 21632
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 6000 21684 6052 21690
rect 6000 21626 6052 21632
rect 4436 21072 4488 21078
rect 4436 21014 4488 21020
rect 4252 21004 4304 21010
rect 4252 20946 4304 20952
rect 4158 20904 4214 20913
rect 4158 20839 4214 20848
rect 4160 20256 4212 20262
rect 4264 20244 4292 20946
rect 4540 20466 4568 21626
rect 5080 21480 5132 21486
rect 5078 21448 5080 21457
rect 5132 21448 5134 21457
rect 5078 21383 5134 21392
rect 6012 21078 6040 21626
rect 7852 21350 7880 22034
rect 8128 21554 8156 22374
rect 8298 22264 8354 22273
rect 8298 22199 8354 22208
rect 8312 22030 8340 22199
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 8116 21548 8168 21554
rect 8116 21490 8168 21496
rect 7932 21480 7984 21486
rect 7932 21422 7984 21428
rect 7840 21344 7892 21350
rect 7838 21312 7840 21321
rect 7892 21312 7894 21321
rect 7838 21247 7894 21256
rect 6000 21072 6052 21078
rect 6000 21014 6052 21020
rect 6092 21004 6144 21010
rect 6092 20946 6144 20952
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5538 20496 5594 20505
rect 4528 20460 4580 20466
rect 5538 20431 5594 20440
rect 4528 20402 4580 20408
rect 5552 20398 5580 20431
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 5722 20360 5778 20369
rect 5448 20324 5500 20330
rect 5722 20295 5778 20304
rect 5448 20266 5500 20272
rect 4212 20216 4292 20244
rect 5080 20256 5132 20262
rect 5078 20224 5080 20233
rect 5356 20256 5408 20262
rect 5132 20224 5134 20233
rect 4160 20198 4212 20204
rect 4172 20058 4200 20198
rect 5356 20198 5408 20204
rect 5078 20159 5134 20168
rect 5170 20088 5226 20097
rect 4160 20052 4212 20058
rect 5170 20023 5226 20032
rect 4160 19994 4212 20000
rect 3976 19984 4028 19990
rect 3976 19926 4028 19932
rect 5080 19984 5132 19990
rect 5080 19926 5132 19932
rect 4712 19916 4764 19922
rect 4712 19858 4764 19864
rect 4160 19712 4212 19718
rect 4160 19654 4212 19660
rect 4068 18828 4120 18834
rect 4172 18816 4200 19654
rect 4724 19514 4752 19858
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 4120 18788 4200 18816
rect 4068 18770 4120 18776
rect 3700 18624 3752 18630
rect 3700 18566 3752 18572
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 3712 18329 3740 18566
rect 3698 18320 3754 18329
rect 3698 18255 3700 18264
rect 3752 18255 3754 18264
rect 3700 18226 3752 18232
rect 3712 18195 3740 18226
rect 4080 18193 4108 18770
rect 5092 18748 5120 19926
rect 5184 19514 5212 20023
rect 5368 19990 5396 20198
rect 5356 19984 5408 19990
rect 5356 19926 5408 19932
rect 5460 19854 5488 20266
rect 5736 20262 5764 20295
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 6104 20058 6132 20946
rect 7196 20936 7248 20942
rect 7196 20878 7248 20884
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6932 20398 6960 20742
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6092 20052 6144 20058
rect 6092 19994 6144 20000
rect 5356 19848 5408 19854
rect 5356 19790 5408 19796
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5368 19242 5396 19790
rect 5356 19236 5408 19242
rect 5356 19178 5408 19184
rect 5172 18760 5224 18766
rect 5092 18720 5172 18748
rect 5172 18702 5224 18708
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 4066 18184 4122 18193
rect 4066 18119 4122 18128
rect 4068 18080 4120 18086
rect 4264 18057 4292 18566
rect 5078 18456 5134 18465
rect 5078 18391 5134 18400
rect 4620 18080 4672 18086
rect 4068 18022 4120 18028
rect 4250 18048 4306 18057
rect 4080 17814 4108 18022
rect 4620 18022 4672 18028
rect 4250 17983 4306 17992
rect 4068 17808 4120 17814
rect 4068 17750 4120 17756
rect 3792 17672 3844 17678
rect 3792 17614 3844 17620
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 3804 17270 3832 17614
rect 3882 17504 3938 17513
rect 3882 17439 3938 17448
rect 3792 17264 3844 17270
rect 3792 17206 3844 17212
rect 3698 16824 3754 16833
rect 3698 16759 3754 16768
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3528 14822 3556 14962
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3422 14648 3478 14657
rect 3422 14583 3478 14592
rect 3332 14476 3384 14482
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 3068 13938 3096 14350
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 3056 13796 3108 13802
rect 3056 13738 3108 13744
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2608 12782 2636 13670
rect 3068 13530 3096 13738
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2596 12776 2648 12782
rect 2516 12736 2596 12764
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2332 10010 2360 11494
rect 2516 11286 2544 12736
rect 2596 12718 2648 12724
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 2608 11529 2636 11562
rect 2594 11520 2650 11529
rect 2594 11455 2650 11464
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2596 10600 2648 10606
rect 2596 10542 2648 10548
rect 2410 10160 2466 10169
rect 2410 10095 2412 10104
rect 2464 10095 2466 10104
rect 2412 10066 2464 10072
rect 2608 10062 2636 10542
rect 2596 10056 2648 10062
rect 2332 9982 2452 10010
rect 2596 9998 2648 10004
rect 2424 9568 2452 9982
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 2516 9761 2544 9862
rect 2502 9752 2558 9761
rect 2502 9687 2558 9696
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2332 9540 2452 9568
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 2240 7313 2268 7890
rect 2226 7304 2282 7313
rect 2226 7239 2282 7248
rect 2332 6934 2360 9540
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 2424 7818 2452 8230
rect 2516 8022 2544 8978
rect 2504 8016 2556 8022
rect 2504 7958 2556 7964
rect 2412 7812 2464 7818
rect 2412 7754 2464 7760
rect 2608 7546 2636 9658
rect 2884 9586 2912 12786
rect 3160 12345 3188 14470
rect 3332 14418 3384 14424
rect 3344 14226 3372 14418
rect 3252 14198 3372 14226
rect 3252 13802 3280 14198
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3240 13796 3292 13802
rect 3240 13738 3292 13744
rect 3240 13456 3292 13462
rect 3240 13398 3292 13404
rect 3146 12336 3202 12345
rect 3146 12271 3202 12280
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 2976 11801 3004 12038
rect 2962 11792 3018 11801
rect 2962 11727 3018 11736
rect 2976 11558 3004 11727
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2976 11218 3004 11494
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 3068 10810 3096 12174
rect 3252 11762 3280 13398
rect 3344 12782 3372 14010
rect 3436 13569 3464 14583
rect 3422 13560 3478 13569
rect 3422 13495 3478 13504
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 3344 12442 3372 12718
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3252 11370 3280 11698
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3160 11354 3280 11370
rect 3344 11354 3372 11630
rect 3148 11348 3280 11354
rect 3200 11342 3280 11348
rect 3332 11348 3384 11354
rect 3148 11290 3200 11296
rect 3332 11290 3384 11296
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3068 10606 3096 10746
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2976 9722 3004 9930
rect 3068 9722 3096 10542
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2884 9178 2912 9522
rect 3068 9178 3096 9658
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2700 8922 2728 9046
rect 2700 8894 2820 8922
rect 2792 8090 2820 8894
rect 2884 8634 2912 9114
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3068 8430 3096 8774
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2792 7698 2820 7890
rect 2792 7670 2912 7698
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2792 7342 2820 7482
rect 2884 7410 2912 7670
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2504 7200 2556 7206
rect 2504 7142 2556 7148
rect 2320 6928 2372 6934
rect 2320 6870 2372 6876
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2134 5672 2190 5681
rect 2134 5607 2190 5616
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2056 5098 2084 5510
rect 2044 5092 2096 5098
rect 2044 5034 2096 5040
rect 2148 5030 2176 5510
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2042 4176 2098 4185
rect 2042 4111 2044 4120
rect 2096 4111 2098 4120
rect 2044 4082 2096 4088
rect 1950 3768 2006 3777
rect 2056 3738 2084 4082
rect 1950 3703 2006 3712
rect 2044 3732 2096 3738
rect 1780 3454 1900 3482
rect 1492 3188 1544 3194
rect 1492 3130 1544 3136
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1780 480 1808 3454
rect 1964 3058 1992 3703
rect 2044 3674 2096 3680
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 1964 2650 1992 2994
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 2056 2310 2084 3538
rect 2148 2836 2176 4966
rect 2240 3194 2268 6802
rect 2516 6769 2544 7142
rect 2502 6760 2558 6769
rect 2502 6695 2558 6704
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2424 6322 2452 6598
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2424 5794 2452 6054
rect 2700 5914 2728 6190
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2424 5766 2544 5794
rect 2320 5636 2372 5642
rect 2320 5578 2372 5584
rect 2332 4758 2360 5578
rect 2320 4752 2372 4758
rect 2320 4694 2372 4700
rect 2332 4282 2360 4694
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2332 3738 2360 4218
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2240 2990 2268 3130
rect 2228 2984 2280 2990
rect 2228 2926 2280 2932
rect 2148 2808 2360 2836
rect 2134 2408 2190 2417
rect 2134 2343 2136 2352
rect 2188 2343 2190 2352
rect 2136 2314 2188 2320
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 2332 480 2360 2808
rect 2516 2689 2544 5766
rect 2502 2680 2558 2689
rect 2502 2615 2504 2624
rect 2556 2615 2558 2624
rect 2504 2586 2556 2592
rect 2516 2555 2544 2586
rect 202 0 258 480
rect 662 0 718 480
rect 1214 0 1270 480
rect 1766 0 1822 480
rect 2318 0 2374 480
rect 2792 377 2820 7278
rect 2884 7002 2912 7346
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2872 5704 2924 5710
rect 2976 5692 3004 8230
rect 3068 7274 3096 8366
rect 3160 7546 3188 11154
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 2924 5664 3004 5692
rect 2872 5646 2924 5652
rect 3252 5166 3280 5714
rect 3344 5545 3372 10950
rect 3436 9926 3464 12582
rect 3528 11898 3556 14758
rect 3620 13326 3648 14758
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 3712 12986 3740 16759
rect 3790 15192 3846 15201
rect 3790 15127 3846 15136
rect 3804 13977 3832 15127
rect 3790 13968 3846 13977
rect 3790 13903 3846 13912
rect 3896 13530 3924 17439
rect 3988 17134 4016 17614
rect 4080 17338 4108 17750
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 3988 16697 4016 17070
rect 4632 16998 4660 18022
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 3974 16688 4030 16697
rect 3974 16623 4030 16632
rect 3988 16522 4016 16623
rect 3976 16516 4028 16522
rect 3976 16458 4028 16464
rect 3988 16046 4016 16458
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3974 15736 4030 15745
rect 4080 15706 4108 16934
rect 4160 16720 4212 16726
rect 4160 16662 4212 16668
rect 4172 16522 4200 16662
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4160 16516 4212 16522
rect 4160 16458 4212 16464
rect 4172 16250 4200 16458
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4172 15706 4200 16186
rect 4448 16046 4476 16594
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 4436 16040 4488 16046
rect 4250 16008 4306 16017
rect 4436 15982 4488 15988
rect 4250 15943 4306 15952
rect 3974 15671 4030 15680
rect 4068 15700 4120 15706
rect 3988 14550 4016 15671
rect 4068 15642 4120 15648
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4068 15360 4120 15366
rect 4120 15308 4200 15314
rect 4068 15302 4200 15308
rect 4080 15286 4200 15302
rect 4172 15162 4200 15286
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4264 14618 4292 15943
rect 4540 15910 4568 16526
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4632 15065 4660 16934
rect 5092 16250 5120 18391
rect 5184 16697 5212 18702
rect 5368 18426 5396 19178
rect 5460 18970 5488 19790
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6012 19446 6040 19654
rect 6104 19514 6132 19994
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 6932 19446 6960 19654
rect 6000 19440 6052 19446
rect 6000 19382 6052 19388
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 7102 19408 7158 19417
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5644 18873 5672 19110
rect 5630 18864 5686 18873
rect 5540 18828 5592 18834
rect 5630 18799 5686 18808
rect 5540 18770 5592 18776
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5552 18290 5580 18770
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6748 18426 6776 19382
rect 6828 19372 6880 19378
rect 7102 19343 7158 19352
rect 6828 19314 6880 19320
rect 6736 18420 6788 18426
rect 6736 18362 6788 18368
rect 6090 18320 6146 18329
rect 5540 18284 5592 18290
rect 5540 18226 5592 18232
rect 5816 18284 5868 18290
rect 6090 18255 6146 18264
rect 6274 18320 6330 18329
rect 6274 18255 6276 18264
rect 5816 18226 5868 18232
rect 5828 17882 5856 18226
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 5816 17876 5868 17882
rect 5816 17818 5868 17824
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5460 17202 5488 17478
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6012 17377 6040 18022
rect 6104 17882 6132 18255
rect 6328 18255 6330 18264
rect 6276 18226 6328 18232
rect 6840 18034 6868 19314
rect 6840 18006 6960 18034
rect 6092 17876 6144 17882
rect 6092 17818 6144 17824
rect 5998 17368 6054 17377
rect 5998 17303 6054 17312
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 5828 16697 5856 17070
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5170 16688 5226 16697
rect 5170 16623 5226 16632
rect 5814 16688 5870 16697
rect 5814 16623 5816 16632
rect 5080 16244 5132 16250
rect 5080 16186 5132 16192
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 4618 15056 4674 15065
rect 4618 14991 4674 15000
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 3976 14544 4028 14550
rect 4028 14492 4108 14498
rect 3976 14486 4108 14492
rect 3988 14470 4108 14486
rect 3988 14421 4016 14470
rect 4080 14074 4108 14470
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 3976 14000 4028 14006
rect 3976 13942 4028 13948
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3884 13320 3936 13326
rect 3882 13288 3884 13297
rect 3936 13288 3938 13297
rect 3882 13223 3938 13232
rect 3700 12980 3752 12986
rect 3700 12922 3752 12928
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3896 11393 3924 12038
rect 3882 11384 3938 11393
rect 3882 11319 3938 11328
rect 3606 11112 3662 11121
rect 3606 11047 3662 11056
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3330 5536 3386 5545
rect 3330 5471 3386 5480
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 3148 5092 3200 5098
rect 3148 5034 3200 5040
rect 2870 4992 2926 5001
rect 2870 4927 2926 4936
rect 2884 480 2912 4927
rect 3160 4826 3188 5034
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3344 4282 3372 4966
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3344 4010 3372 4218
rect 3332 4004 3384 4010
rect 3252 3964 3332 3992
rect 3252 2650 3280 3964
rect 3332 3946 3384 3952
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3344 2990 3372 3470
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 2976 2417 3004 2450
rect 3252 2446 3280 2586
rect 3436 2553 3464 9318
rect 3514 7304 3570 7313
rect 3514 7239 3570 7248
rect 3528 7206 3556 7239
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3528 6662 3556 7142
rect 3620 6905 3648 11047
rect 3698 10024 3754 10033
rect 3698 9959 3754 9968
rect 3712 8634 3740 9959
rect 3882 9480 3938 9489
rect 3882 9415 3938 9424
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3698 8528 3754 8537
rect 3698 8463 3754 8472
rect 3606 6896 3662 6905
rect 3606 6831 3662 6840
rect 3712 6746 3740 8463
rect 3620 6718 3740 6746
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3528 3398 3556 6598
rect 3620 5012 3648 6718
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3712 5166 3740 5850
rect 3700 5160 3752 5166
rect 3698 5128 3700 5137
rect 3752 5128 3754 5137
rect 3698 5063 3754 5072
rect 3620 4984 3740 5012
rect 3606 4856 3662 4865
rect 3606 4791 3662 4800
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3528 3058 3556 3334
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3422 2544 3478 2553
rect 3422 2479 3478 2488
rect 3240 2440 3292 2446
rect 2962 2408 3018 2417
rect 3240 2382 3292 2388
rect 2962 2343 3018 2352
rect 3620 1873 3648 4791
rect 3712 4321 3740 4984
rect 3698 4312 3754 4321
rect 3698 4247 3754 4256
rect 3606 1864 3662 1873
rect 3606 1799 3662 1808
rect 3804 1601 3832 9318
rect 3896 7528 3924 9415
rect 3988 9042 4016 13942
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4080 12986 4108 13330
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 4356 12442 4384 12650
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4172 12345 4200 12378
rect 4158 12336 4214 12345
rect 4158 12271 4214 12280
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4356 12102 4384 12242
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4080 10266 4108 11086
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4172 10198 4200 11154
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4080 9654 4108 10066
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 4080 9178 4108 9590
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4066 9072 4122 9081
rect 3976 9036 4028 9042
rect 4066 9007 4122 9016
rect 3976 8978 4028 8984
rect 3988 8634 4016 8978
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4080 8537 4108 9007
rect 4066 8528 4122 8537
rect 4066 8463 4122 8472
rect 4172 7698 4200 9318
rect 4264 7818 4292 10746
rect 4356 9110 4384 12038
rect 4632 11234 4660 14991
rect 4712 14884 4764 14890
rect 4712 14826 4764 14832
rect 4724 14414 4752 14826
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4712 14408 4764 14414
rect 4710 14376 4712 14385
rect 4764 14376 4766 14385
rect 4710 14311 4766 14320
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4540 11206 4660 11234
rect 4434 10568 4490 10577
rect 4434 10503 4490 10512
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4356 8537 4384 8910
rect 4342 8528 4398 8537
rect 4448 8498 4476 10503
rect 4540 9586 4568 11206
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4632 10810 4660 11086
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4724 10470 4752 12582
rect 4816 12345 4844 13126
rect 4802 12336 4858 12345
rect 4802 12271 4858 12280
rect 4816 12102 4844 12271
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4724 8634 4752 8978
rect 4816 8838 4844 9998
rect 4908 9450 4936 14758
rect 5000 10305 5028 15846
rect 5184 15570 5212 16623
rect 5868 16623 5870 16632
rect 5816 16594 5868 16600
rect 5540 16584 5592 16590
rect 5828 16563 5856 16594
rect 5540 16526 5592 16532
rect 5356 16516 5408 16522
rect 5356 16458 5408 16464
rect 5368 15910 5396 16458
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5460 16114 5488 16390
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 5172 15564 5224 15570
rect 5172 15506 5224 15512
rect 5184 14770 5212 15506
rect 5092 14742 5212 14770
rect 5092 14482 5120 14742
rect 5170 14648 5226 14657
rect 5170 14583 5226 14592
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 5092 12481 5120 12582
rect 5078 12472 5134 12481
rect 5078 12407 5134 12416
rect 5184 12288 5212 14583
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5276 13870 5304 14418
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5368 13274 5396 15846
rect 5552 15722 5580 16526
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5552 15706 5672 15722
rect 5552 15700 5684 15706
rect 5552 15694 5632 15700
rect 5632 15642 5684 15648
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5552 15026 5580 15574
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5630 15056 5686 15065
rect 5540 15020 5592 15026
rect 5630 14991 5686 15000
rect 5540 14962 5592 14968
rect 5644 14906 5672 14991
rect 5552 14878 5672 14906
rect 5552 14822 5580 14878
rect 5540 14816 5592 14822
rect 5632 14816 5684 14822
rect 5540 14758 5592 14764
rect 5630 14784 5632 14793
rect 5684 14784 5686 14793
rect 5630 14719 5686 14728
rect 6012 14346 6040 16934
rect 6104 16726 6132 17818
rect 6368 17740 6420 17746
rect 6368 17682 6420 17688
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6196 17134 6224 17478
rect 6380 17202 6408 17682
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6184 17128 6236 17134
rect 6184 17070 6236 17076
rect 6932 16998 6960 18006
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 6932 16726 6960 16934
rect 6092 16720 6144 16726
rect 6092 16662 6144 16668
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 7116 16674 7144 19343
rect 7208 19310 7236 20878
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7392 19854 7420 20334
rect 7380 19848 7432 19854
rect 7380 19790 7432 19796
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7300 19378 7328 19654
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 7300 18970 7328 19314
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7392 18630 7420 18770
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7392 18154 7420 18566
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7380 18148 7432 18154
rect 7380 18090 7432 18096
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 17066 7236 17478
rect 7196 17060 7248 17066
rect 7196 17002 7248 17008
rect 7208 16794 7236 17002
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 6104 16250 6132 16662
rect 7116 16646 7236 16674
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5460 13530 5488 13738
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 5276 12442 5304 13262
rect 5368 13246 5488 13274
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5264 12300 5316 12306
rect 5184 12260 5264 12288
rect 5264 12242 5316 12248
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5184 11558 5212 12038
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5184 10538 5212 11494
rect 5276 11354 5304 12242
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 4986 10296 5042 10305
rect 4986 10231 5042 10240
rect 5184 9926 5212 10474
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5354 9888 5410 9897
rect 4896 9444 4948 9450
rect 4896 9386 4948 9392
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4342 8463 4398 8472
rect 4436 8492 4488 8498
rect 4356 8090 4384 8463
rect 4436 8434 4488 8440
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 4172 7670 4292 7698
rect 4160 7540 4212 7546
rect 3896 7500 4160 7528
rect 4160 7482 4212 7488
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 3896 6934 3924 7210
rect 4066 7168 4122 7177
rect 4066 7103 4122 7112
rect 3884 6928 3936 6934
rect 3884 6870 3936 6876
rect 4080 6474 4108 7103
rect 4080 6458 4200 6474
rect 4080 6452 4212 6458
rect 4080 6446 4160 6452
rect 4160 6394 4212 6400
rect 4160 5568 4212 5574
rect 3974 5536 4030 5545
rect 4160 5510 4212 5516
rect 3974 5471 4030 5480
rect 3882 5128 3938 5137
rect 3882 5063 3938 5072
rect 3790 1592 3846 1601
rect 3790 1527 3846 1536
rect 3896 1442 3924 5063
rect 3988 4865 4016 5471
rect 3974 4856 4030 4865
rect 4172 4842 4200 5510
rect 4080 4826 4200 4842
rect 3974 4791 4030 4800
rect 4068 4820 4200 4826
rect 4120 4814 4200 4820
rect 4068 4762 4120 4768
rect 3974 3768 4030 3777
rect 3974 3703 4030 3712
rect 3436 1414 3924 1442
rect 3436 480 3464 1414
rect 3988 480 4016 3703
rect 4080 2990 4108 4762
rect 4264 3233 4292 7670
rect 4356 6866 4384 8026
rect 4816 7206 4844 8774
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4356 6390 4384 6802
rect 4526 6760 4582 6769
rect 4526 6695 4582 6704
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4448 5030 4476 5646
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 4250 3224 4306 3233
rect 4356 3194 4384 3946
rect 4448 3777 4476 4966
rect 4434 3768 4490 3777
rect 4434 3703 4490 3712
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4250 3159 4306 3168
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4448 3058 4476 3334
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 4448 2514 4476 2994
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 4540 480 4568 6695
rect 4618 6624 4674 6633
rect 4618 6559 4674 6568
rect 4632 5914 4660 6559
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4632 5370 4660 5850
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4710 5400 4766 5409
rect 4620 5364 4672 5370
rect 4710 5335 4766 5344
rect 4620 5306 4672 5312
rect 4724 4690 4752 5335
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 4816 4622 4844 5646
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4632 3942 4660 4558
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4632 2990 4660 3878
rect 4724 3738 4752 4082
rect 4816 4078 4844 4218
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4632 2582 4660 2926
rect 4724 2922 4752 3674
rect 4816 3398 4844 4014
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 4620 2576 4672 2582
rect 4620 2518 4672 2524
rect 4908 2009 4936 9046
rect 5184 8906 5212 9862
rect 5354 9823 5410 9832
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 5184 8401 5212 8502
rect 5170 8392 5226 8401
rect 5170 8327 5226 8336
rect 5078 8120 5134 8129
rect 5078 8055 5134 8064
rect 5092 8022 5120 8055
rect 5276 8022 5304 9522
rect 5368 9466 5396 9823
rect 5460 9568 5488 13246
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 5552 12345 5580 12650
rect 6012 12646 6040 13330
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 5538 12336 5594 12345
rect 6104 12306 6132 16050
rect 6828 15904 6880 15910
rect 6880 15852 6960 15858
rect 6828 15846 6960 15852
rect 6840 15830 6960 15846
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 6380 14618 6408 14962
rect 6748 14657 6776 15642
rect 6734 14648 6790 14657
rect 6368 14612 6420 14618
rect 6932 14618 6960 15830
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6734 14583 6790 14592
rect 6920 14612 6972 14618
rect 6368 14554 6420 14560
rect 6920 14554 6972 14560
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6182 13832 6238 13841
rect 6182 13767 6238 13776
rect 5538 12271 5594 12280
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 11880 5580 12174
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6000 11892 6052 11898
rect 5552 11852 5672 11880
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5552 10810 5580 11630
rect 5644 11626 5672 11852
rect 6000 11834 6052 11840
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5644 11218 5672 11562
rect 6012 11286 6040 11834
rect 6104 11558 6132 12242
rect 6196 11801 6224 13767
rect 6276 13728 6328 13734
rect 6276 13670 6328 13676
rect 6288 13297 6316 13670
rect 6380 13462 6408 14214
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6368 13456 6420 13462
rect 6368 13398 6420 13404
rect 6458 13424 6514 13433
rect 6458 13359 6514 13368
rect 6274 13288 6330 13297
rect 6274 13223 6330 13232
rect 6366 12608 6422 12617
rect 6366 12543 6422 12552
rect 6182 11792 6238 11801
rect 6182 11727 6238 11736
rect 6380 11642 6408 12543
rect 6196 11614 6408 11642
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6090 11384 6146 11393
rect 6090 11319 6146 11328
rect 6000 11280 6052 11286
rect 6000 11222 6052 11228
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6012 10810 6040 11222
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 6012 10044 6040 10542
rect 6104 10266 6132 11319
rect 6196 10606 6224 11614
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6366 11520 6422 11529
rect 6288 11354 6316 11494
rect 6366 11455 6422 11464
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6380 11234 6408 11455
rect 6288 11206 6408 11234
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6196 10062 6224 10406
rect 6092 10056 6144 10062
rect 6012 10016 6092 10044
rect 6092 9998 6144 10004
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5998 9752 6054 9761
rect 5998 9687 6054 9696
rect 5540 9580 5592 9586
rect 5460 9540 5540 9568
rect 5540 9522 5592 9528
rect 5368 9438 5580 9466
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5368 8362 5396 8774
rect 5552 8548 5580 9438
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6012 8616 6040 9687
rect 6104 9382 6132 9998
rect 6196 9654 6224 9998
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6196 9081 6224 9318
rect 6182 9072 6238 9081
rect 6182 9007 6238 9016
rect 6012 8588 6224 8616
rect 5552 8520 5672 8548
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5092 7002 5120 7958
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5184 7041 5212 7142
rect 5170 7032 5226 7041
rect 5080 6996 5132 7002
rect 5170 6967 5226 6976
rect 5080 6938 5132 6944
rect 5078 5672 5134 5681
rect 5078 5607 5134 5616
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5000 4185 5028 5102
rect 4986 4176 5042 4185
rect 4986 4111 5042 4120
rect 4894 2000 4950 2009
rect 4894 1935 4950 1944
rect 5092 480 5120 5607
rect 5172 5024 5224 5030
rect 5276 5012 5304 7210
rect 5368 5370 5396 8298
rect 5552 8106 5580 8366
rect 5460 8090 5580 8106
rect 5448 8084 5580 8090
rect 5500 8078 5580 8084
rect 5448 8026 5500 8032
rect 5644 7857 5672 8520
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 5630 7848 5686 7857
rect 5630 7783 5686 7792
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 7206 5488 7686
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5460 6866 5488 7142
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 6012 6644 6040 8434
rect 6092 6656 6144 6662
rect 6012 6616 6092 6644
rect 5460 5778 5488 6598
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5552 5914 5580 6326
rect 6012 6322 6040 6616
rect 6092 6598 6144 6604
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6012 5914 6040 6258
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5224 4984 5304 5012
rect 5172 4966 5224 4972
rect 5184 4486 5212 4966
rect 5460 4622 5488 5714
rect 5552 5234 5580 5850
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5460 4282 5488 4558
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 5184 3738 5212 3946
rect 5448 3936 5500 3942
rect 5552 3924 5580 4694
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6012 4078 6040 5850
rect 6090 5808 6146 5817
rect 6090 5743 6146 5752
rect 6104 5166 6132 5743
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 6092 5024 6144 5030
rect 6090 4992 6092 5001
rect 6144 4992 6146 5001
rect 6090 4927 6146 4936
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 5500 3896 5580 3924
rect 5448 3878 5500 3884
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5460 3534 5488 3878
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5184 1601 5212 3334
rect 5460 3194 5488 3470
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 5736 2650 5764 2858
rect 5998 2680 6054 2689
rect 5724 2644 5776 2650
rect 5998 2615 6000 2624
rect 5724 2586 5776 2592
rect 6052 2615 6054 2624
rect 6000 2586 6052 2592
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5632 2032 5684 2038
rect 5632 1974 5684 1980
rect 5170 1592 5226 1601
rect 5170 1527 5226 1536
rect 5644 480 5672 1974
rect 6196 480 6224 8588
rect 6288 2038 6316 11206
rect 6368 10192 6420 10198
rect 6368 10134 6420 10140
rect 6380 9450 6408 10134
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6366 9344 6422 9353
rect 6366 9279 6422 9288
rect 6380 9042 6408 9279
rect 6472 9217 6500 13359
rect 6458 9208 6514 9217
rect 6564 9178 6592 13874
rect 6656 11898 6684 14010
rect 6932 13870 6960 14350
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6748 13258 6776 13738
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 6840 13025 6868 13670
rect 6826 13016 6882 13025
rect 6826 12951 6882 12960
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6748 12458 6776 12582
rect 6748 12442 6868 12458
rect 6748 12436 6880 12442
rect 6748 12430 6828 12436
rect 6828 12378 6880 12384
rect 6840 12347 6868 12378
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6932 11642 6960 13806
rect 7024 12442 7052 15302
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7116 12345 7144 12582
rect 7102 12336 7158 12345
rect 7102 12271 7158 12280
rect 6656 11614 6960 11642
rect 7010 11656 7066 11665
rect 6458 9143 6514 9152
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6366 6896 6422 6905
rect 6366 6831 6422 6840
rect 6380 4457 6408 6831
rect 6366 4448 6422 4457
rect 6366 4383 6422 4392
rect 6368 2440 6420 2446
rect 6366 2408 6368 2417
rect 6420 2408 6422 2417
rect 6366 2343 6422 2352
rect 6276 2032 6328 2038
rect 6276 1974 6328 1980
rect 6472 921 6500 8570
rect 6564 8129 6592 9114
rect 6550 8120 6606 8129
rect 6550 8055 6606 8064
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6564 5370 6592 5714
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6564 4729 6592 5034
rect 6550 4720 6606 4729
rect 6550 4655 6606 4664
rect 6656 3482 6684 11614
rect 7010 11591 7066 11600
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6932 10810 6960 11494
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6826 10160 6882 10169
rect 6826 10095 6882 10104
rect 6734 10024 6790 10033
rect 6734 9959 6736 9968
rect 6788 9959 6790 9968
rect 6736 9930 6788 9936
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6748 8090 6776 8978
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6840 7410 6868 10095
rect 6932 10033 6960 10474
rect 6918 10024 6974 10033
rect 6918 9959 6974 9968
rect 7024 9897 7052 11591
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7116 10044 7144 11290
rect 7208 10266 7236 16646
rect 7286 15736 7342 15745
rect 7286 15671 7288 15680
rect 7340 15671 7342 15680
rect 7288 15642 7340 15648
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 7300 14822 7328 15438
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7196 10056 7248 10062
rect 7116 10016 7196 10044
rect 7010 9888 7066 9897
rect 7010 9823 7066 9832
rect 7116 9489 7144 10016
rect 7196 9998 7248 10004
rect 7196 9512 7248 9518
rect 7102 9480 7158 9489
rect 7196 9454 7248 9460
rect 7102 9415 7158 9424
rect 7116 9382 7144 9415
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7116 8634 7144 9318
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6748 6610 6776 6802
rect 6932 6610 6960 8434
rect 7102 8392 7158 8401
rect 7102 8327 7158 8336
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 7024 7750 7052 8230
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6748 6582 6960 6610
rect 6748 6390 6776 6582
rect 6826 6488 6882 6497
rect 6826 6423 6828 6432
rect 6880 6423 6882 6432
rect 6828 6394 6880 6400
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 6748 4826 6776 6326
rect 7024 5137 7052 7686
rect 7116 6866 7144 8327
rect 7208 7886 7236 9454
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7208 7206 7236 7822
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7116 6186 7144 6802
rect 7104 6180 7156 6186
rect 7104 6122 7156 6128
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7010 5128 7066 5137
rect 7010 5063 7066 5072
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6840 4078 6868 4966
rect 7024 4321 7052 5063
rect 7116 4486 7144 5170
rect 7300 4604 7328 14758
rect 7392 13190 7420 18090
rect 7656 18080 7708 18086
rect 7654 18048 7656 18057
rect 7708 18048 7710 18057
rect 7654 17983 7710 17992
rect 7760 17610 7788 18226
rect 7748 17604 7800 17610
rect 7748 17546 7800 17552
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 7484 16046 7512 16662
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7668 14890 7696 15506
rect 7656 14884 7708 14890
rect 7656 14826 7708 14832
rect 7562 14784 7618 14793
rect 7562 14719 7618 14728
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7392 12646 7420 13126
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7380 12640 7432 12646
rect 7378 12608 7380 12617
rect 7432 12608 7434 12617
rect 7378 12543 7434 12552
rect 7484 12442 7512 12786
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7392 10810 7420 10950
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7392 9625 7420 10066
rect 7378 9616 7434 9625
rect 7378 9551 7434 9560
rect 7392 9382 7420 9551
rect 7484 9450 7512 12378
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 9110 7420 9318
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7484 7857 7512 7890
rect 7470 7848 7526 7857
rect 7470 7783 7526 7792
rect 7484 7546 7512 7783
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7378 6352 7434 6361
rect 7378 6287 7380 6296
rect 7432 6287 7434 6296
rect 7380 6258 7432 6264
rect 7392 5914 7420 6258
rect 7484 6254 7512 6598
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7300 4576 7420 4604
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7010 4312 7066 4321
rect 7010 4247 7066 4256
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6748 3602 6776 3878
rect 6840 3670 6868 4014
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6656 3454 6776 3482
rect 6458 912 6514 921
rect 6458 847 6514 856
rect 6748 480 6776 3454
rect 7024 2854 7052 3606
rect 7116 3466 7144 4422
rect 7300 4146 7328 4422
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7300 3738 7328 4082
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7194 3632 7250 3641
rect 7194 3567 7196 3576
rect 7248 3567 7250 3576
rect 7196 3538 7248 3544
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7116 2990 7144 3402
rect 7208 3194 7236 3538
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7012 2848 7064 2854
rect 7010 2816 7012 2825
rect 7064 2816 7066 2825
rect 7392 2802 7420 4576
rect 7472 3392 7524 3398
rect 7576 3380 7604 14719
rect 7668 14113 7696 14826
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 7654 14104 7710 14113
rect 7654 14039 7710 14048
rect 7760 13870 7788 14486
rect 7840 14408 7892 14414
rect 7840 14350 7892 14356
rect 7852 14074 7880 14350
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 7748 13864 7800 13870
rect 7840 13864 7892 13870
rect 7748 13806 7800 13812
rect 7838 13832 7840 13841
rect 7892 13832 7894 13841
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7668 12102 7696 13262
rect 7760 12288 7788 13806
rect 7838 13767 7894 13776
rect 7944 12442 7972 21422
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 8220 19922 8248 20198
rect 8208 19916 8260 19922
rect 8208 19858 8260 19864
rect 8220 19174 8248 19858
rect 9324 19718 9352 20198
rect 8668 19712 8720 19718
rect 8668 19654 8720 19660
rect 9036 19712 9088 19718
rect 9036 19654 9088 19660
rect 9312 19712 9364 19718
rect 9312 19654 9364 19660
rect 8680 19310 8708 19654
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8220 18766 8248 19110
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8208 18760 8260 18766
rect 8022 18728 8078 18737
rect 8260 18720 8340 18748
rect 8208 18702 8260 18708
rect 8022 18663 8078 18672
rect 8036 16794 8064 18663
rect 8312 17882 8340 18720
rect 8404 18222 8432 18770
rect 9048 18630 9076 19654
rect 9324 19242 9352 19654
rect 9312 19236 9364 19242
rect 9312 19178 9364 19184
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 8392 18216 8444 18222
rect 8390 18184 8392 18193
rect 8444 18184 8446 18193
rect 8390 18119 8446 18128
rect 8496 18034 8524 18566
rect 9232 18426 9260 18770
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 8404 18006 8524 18034
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8404 17762 8432 18006
rect 9232 17882 9260 18362
rect 9324 18222 9352 19178
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9508 18970 9536 19110
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 8220 17734 8432 17762
rect 8116 17264 8168 17270
rect 8116 17206 8168 17212
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 8036 15910 8064 16594
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 7760 12260 7972 12288
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7668 10985 7696 12038
rect 7760 11898 7788 12106
rect 7944 11937 7972 12260
rect 7930 11928 7986 11937
rect 7748 11892 7800 11898
rect 7930 11863 7986 11872
rect 7748 11834 7800 11840
rect 8036 11778 8064 15846
rect 8128 15162 8156 17206
rect 8220 17134 8248 17734
rect 9324 17270 9352 18158
rect 9416 17882 9444 18158
rect 9494 18048 9550 18057
rect 9494 17983 9550 17992
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9312 17264 9364 17270
rect 9312 17206 9364 17212
rect 8208 17128 8260 17134
rect 9312 17128 9364 17134
rect 8208 17070 8260 17076
rect 9232 17088 9312 17116
rect 8220 16726 8248 17070
rect 8208 16720 8260 16726
rect 8206 16688 8208 16697
rect 8260 16688 8262 16697
rect 8206 16623 8262 16632
rect 8220 15978 8248 16623
rect 8668 16584 8720 16590
rect 8668 16526 8720 16532
rect 8392 16516 8444 16522
rect 8392 16458 8444 16464
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 8404 15366 8432 16458
rect 8680 15706 8708 16526
rect 9232 16454 9260 17088
rect 9312 17070 9364 17076
rect 9220 16448 9272 16454
rect 9220 16390 9272 16396
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8392 15360 8444 15366
rect 8390 15328 8392 15337
rect 8444 15328 8446 15337
rect 8390 15263 8446 15272
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8666 14920 8722 14929
rect 8772 14906 8800 15846
rect 9232 15366 9260 16390
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 8722 14878 8800 14906
rect 8666 14855 8668 14864
rect 8720 14855 8722 14864
rect 8668 14826 8720 14832
rect 8680 14618 8708 14826
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 8758 14648 8814 14657
rect 8668 14612 8720 14618
rect 8758 14583 8760 14592
rect 8668 14554 8720 14560
rect 8812 14583 8814 14592
rect 8760 14554 8812 14560
rect 9140 14550 9168 14758
rect 8116 14544 8168 14550
rect 9128 14544 9180 14550
rect 8116 14486 8168 14492
rect 9126 14512 9128 14521
rect 9180 14512 9182 14521
rect 8128 13870 8156 14486
rect 9126 14447 9182 14456
rect 9140 14421 9168 14447
rect 8944 14340 8996 14346
rect 8944 14282 8996 14288
rect 8298 14104 8354 14113
rect 8298 14039 8354 14048
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 8116 13728 8168 13734
rect 8116 13670 8168 13676
rect 7852 11750 8064 11778
rect 7654 10976 7710 10985
rect 7654 10911 7710 10920
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7654 10432 7710 10441
rect 7654 10367 7710 10376
rect 7668 8090 7696 10367
rect 7760 10198 7788 10678
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7852 10130 7880 11750
rect 8128 11286 8156 13670
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8220 12646 8248 13262
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8116 11280 8168 11286
rect 8220 11257 8248 12582
rect 8312 11354 8340 14039
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8588 12918 8616 13330
rect 8576 12912 8628 12918
rect 8574 12880 8576 12889
rect 8628 12880 8630 12889
rect 8574 12815 8630 12824
rect 8392 12708 8444 12714
rect 8392 12650 8444 12656
rect 8668 12708 8720 12714
rect 8668 12650 8720 12656
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8116 11222 8168 11228
rect 8206 11248 8262 11257
rect 8022 11112 8078 11121
rect 8022 11047 8078 11056
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7944 10266 7972 10746
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 8036 9042 8064 11047
rect 8128 10674 8156 11222
rect 8206 11183 8262 11192
rect 8220 11098 8248 11183
rect 8220 11070 8340 11098
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8128 10266 8156 10610
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8116 10056 8168 10062
rect 8220 10044 8248 10950
rect 8168 10016 8248 10044
rect 8116 9998 8168 10004
rect 8128 9178 8156 9998
rect 8312 9353 8340 11070
rect 8404 10810 8432 12650
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8496 11626 8524 12174
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8496 11354 8524 11562
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8680 11121 8708 12650
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8772 12442 8800 12582
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8772 11898 8800 12378
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8852 11620 8904 11626
rect 8852 11562 8904 11568
rect 8666 11112 8722 11121
rect 8666 11047 8722 11056
rect 8864 10849 8892 11562
rect 8850 10840 8906 10849
rect 8392 10804 8444 10810
rect 8850 10775 8906 10784
rect 8392 10746 8444 10752
rect 8404 10538 8432 10746
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8390 10296 8446 10305
rect 8390 10231 8446 10240
rect 8298 9344 8354 9353
rect 8298 9279 8354 9288
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8298 8936 8354 8945
rect 8298 8871 8354 8880
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 7760 8430 7788 8774
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7746 6760 7802 6769
rect 7746 6695 7748 6704
rect 7800 6695 7802 6704
rect 7748 6666 7800 6672
rect 7852 5681 7880 8298
rect 7838 5672 7894 5681
rect 7838 5607 7894 5616
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 7944 4282 7972 5102
rect 8036 4729 8064 8774
rect 8312 8634 8340 8871
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8298 8528 8354 8537
rect 8298 8463 8300 8472
rect 8352 8463 8354 8472
rect 8300 8434 8352 8440
rect 8208 7200 8260 7206
rect 8260 7160 8340 7188
rect 8208 7142 8260 7148
rect 8206 7032 8262 7041
rect 8206 6967 8262 6976
rect 8220 6866 8248 6967
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8128 6458 8156 6802
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8128 5914 8156 6394
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8220 5778 8248 6802
rect 8312 6730 8340 7160
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8300 5636 8352 5642
rect 8220 5596 8300 5624
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8022 4720 8078 4729
rect 8022 4655 8078 4664
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 7944 4078 7972 4218
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8128 4010 8156 5034
rect 8220 4826 8248 5596
rect 8300 5578 8352 5584
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8312 4706 8340 4966
rect 8220 4678 8340 4706
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 8114 3768 8170 3777
rect 8114 3703 8116 3712
rect 8168 3703 8170 3712
rect 8116 3674 8168 3680
rect 7576 3352 7788 3380
rect 7472 3334 7524 3340
rect 7484 2990 7512 3334
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7010 2751 7066 2760
rect 7208 2774 7420 2802
rect 7208 2666 7236 2774
rect 7208 2638 7328 2666
rect 7300 480 7328 2638
rect 7484 2514 7512 2926
rect 7760 2666 7788 3352
rect 8220 3126 8248 4678
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8312 3738 8340 4558
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 7760 2638 7880 2666
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 7852 480 7880 2638
rect 8404 480 8432 10231
rect 8852 9376 8904 9382
rect 8850 9344 8852 9353
rect 8904 9344 8906 9353
rect 8850 9279 8906 9288
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8496 8362 8524 9046
rect 8850 8664 8906 8673
rect 8850 8599 8852 8608
rect 8904 8599 8906 8608
rect 8852 8570 8904 8576
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8496 5234 8524 8298
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8588 7342 8616 7686
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8588 6798 8616 7278
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8588 6458 8616 6734
rect 8772 6662 8800 7482
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8772 5914 8800 6598
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8772 5370 8800 5850
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8772 4826 8800 5306
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8588 3738 8616 4626
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8680 3398 8708 4558
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8680 2582 8708 3334
rect 8772 2922 8800 4762
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8956 480 8984 14282
rect 9232 13433 9260 15302
rect 9324 14618 9352 15506
rect 9508 15042 9536 17983
rect 9600 15178 9628 22374
rect 9954 22335 10010 22344
rect 9770 22128 9826 22137
rect 9770 22063 9826 22072
rect 9678 21312 9734 21321
rect 9678 21247 9734 21256
rect 9692 21146 9720 21247
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9784 18970 9812 22063
rect 9864 19984 9916 19990
rect 9864 19926 9916 19932
rect 9876 19378 9904 19926
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9876 19174 9904 19314
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9784 17270 9812 17614
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9784 16590 9812 17206
rect 9876 17134 9904 17682
rect 9968 17338 9996 22335
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 10690 21448 10746 21457
rect 10690 21383 10746 21392
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 10060 21146 10088 21286
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 10060 20602 10088 21082
rect 10704 20942 10732 21383
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 10692 20936 10744 20942
rect 10692 20878 10744 20884
rect 10152 20602 10180 20878
rect 10048 20596 10100 20602
rect 10048 20538 10100 20544
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10152 19514 10180 20538
rect 10704 20534 10732 20878
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 10692 20528 10744 20534
rect 10692 20470 10744 20476
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10704 20058 10732 20470
rect 12622 20360 12678 20369
rect 12622 20295 12678 20304
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 10060 17785 10088 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10980 19009 11008 19246
rect 10966 19000 11022 19009
rect 10966 18935 11022 18944
rect 11242 18864 11298 18873
rect 11242 18799 11298 18808
rect 10140 18760 10192 18766
rect 10138 18728 10140 18737
rect 10324 18760 10376 18766
rect 10192 18728 10194 18737
rect 10194 18686 10272 18714
rect 10324 18702 10376 18708
rect 10968 18760 11020 18766
rect 11020 18720 11100 18748
rect 10968 18702 11020 18708
rect 10138 18663 10194 18672
rect 10244 18426 10272 18686
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10336 18222 10364 18702
rect 10692 18352 10744 18358
rect 10690 18320 10692 18329
rect 10744 18320 10746 18329
rect 10690 18255 10746 18264
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 11072 17882 11100 18720
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 10046 17776 10102 17785
rect 10046 17711 10102 17720
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 11256 17202 11284 18799
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9876 16658 9904 17070
rect 10704 16998 10732 17138
rect 11336 17128 11388 17134
rect 11336 17070 11388 17076
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10692 16992 10744 16998
rect 10796 16969 10824 17002
rect 10692 16934 10744 16940
rect 10782 16960 10838 16969
rect 10152 16794 10180 16934
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9600 15162 9720 15178
rect 9600 15156 9732 15162
rect 9600 15150 9680 15156
rect 9680 15098 9732 15104
rect 9784 15065 9812 15846
rect 9968 15570 9996 16526
rect 10060 15706 10088 16594
rect 10152 16250 10180 16730
rect 10704 16658 10732 16934
rect 10782 16895 10838 16904
rect 11348 16794 11376 17070
rect 12084 16998 12112 18022
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 12438 16960 12494 16969
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11242 16688 11298 16697
rect 10692 16652 10744 16658
rect 11242 16623 11298 16632
rect 10692 16594 10744 16600
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10704 15638 10732 16050
rect 11256 15910 11284 16623
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 11072 15162 11100 15574
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 9770 15056 9826 15065
rect 9508 15014 9628 15042
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9324 13530 9352 14554
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9218 13424 9274 13433
rect 9218 13359 9274 13368
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 9324 12714 9352 13330
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9128 12232 9180 12238
rect 9126 12200 9128 12209
rect 9180 12200 9182 12209
rect 9126 12135 9182 12144
rect 9140 11218 9168 12135
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9232 11082 9260 11562
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9140 10130 9168 10406
rect 9416 10198 9444 10406
rect 9404 10192 9456 10198
rect 9404 10134 9456 10140
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9140 9178 9168 10066
rect 9416 9926 9444 10134
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9508 9722 9536 10610
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9048 7750 9076 8230
rect 9324 7750 9352 8842
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9508 8498 9536 8774
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9508 8401 9536 8434
rect 9494 8392 9550 8401
rect 9494 8327 9550 8336
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9048 7002 9076 7686
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9140 5914 9168 6598
rect 9324 6225 9352 7686
rect 9508 7585 9536 8026
rect 9494 7576 9550 7585
rect 9494 7511 9550 7520
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9416 6633 9444 7142
rect 9402 6624 9458 6633
rect 9402 6559 9458 6568
rect 9416 6254 9444 6559
rect 9404 6248 9456 6254
rect 9310 6216 9366 6225
rect 9404 6190 9456 6196
rect 9310 6151 9366 6160
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9416 5030 9444 5714
rect 9600 5624 9628 15014
rect 9770 14991 9826 15000
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10048 14884 10100 14890
rect 10048 14826 10100 14832
rect 9954 14104 10010 14113
rect 10060 14074 10088 14826
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14550 10732 14962
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10692 14544 10744 14550
rect 10692 14486 10744 14492
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 9954 14039 10010 14048
rect 10048 14068 10100 14074
rect 9968 13734 9996 14039
rect 10048 14010 10100 14016
rect 10152 13841 10180 14418
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10138 13832 10194 13841
rect 10138 13767 10194 13776
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9968 13530 9996 13670
rect 10046 13560 10102 13569
rect 9956 13524 10008 13530
rect 10046 13495 10102 13504
rect 9956 13466 10008 13472
rect 10060 12866 10088 13495
rect 10152 13394 10180 13767
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13462 10732 13874
rect 10796 13705 10824 14758
rect 10782 13696 10838 13705
rect 10782 13631 10838 13640
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10152 12986 10180 13330
rect 10704 12986 10732 13398
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 9772 12844 9824 12850
rect 10060 12838 10364 12866
rect 9772 12786 9824 12792
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 9692 12102 9720 12650
rect 9784 12306 9812 12786
rect 10336 12753 10364 12838
rect 10138 12744 10194 12753
rect 10048 12708 10100 12714
rect 10138 12679 10194 12688
rect 10322 12744 10378 12753
rect 10322 12679 10378 12688
rect 10048 12650 10100 12656
rect 10060 12442 10088 12650
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9784 11762 9812 12242
rect 10152 12073 10180 12679
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10138 12064 10194 12073
rect 10138 11999 10194 12008
rect 10046 11928 10102 11937
rect 10046 11863 10102 11872
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 10060 11218 10088 11863
rect 10140 11552 10192 11558
rect 10612 11540 10640 12310
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10704 11762 10732 12174
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10692 11552 10744 11558
rect 10612 11512 10692 11540
rect 10140 11494 10192 11500
rect 10692 11494 10744 11500
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9678 10976 9734 10985
rect 9678 10911 9734 10920
rect 9692 10810 9720 10911
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9784 9450 9812 11018
rect 9968 10470 9996 11086
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9692 8514 9720 8978
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9784 8634 9812 8910
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9692 8486 9812 8514
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9692 8090 9720 8366
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9692 7546 9720 8026
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9692 7342 9720 7482
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9508 5596 9628 5624
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 9416 4486 9444 4626
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9416 4282 9444 4422
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 9048 2990 9076 3946
rect 9416 3942 9444 4082
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9140 3369 9168 3878
rect 9416 3398 9444 3878
rect 9404 3392 9456 3398
rect 9126 3360 9182 3369
rect 9404 3334 9456 3340
rect 9126 3295 9182 3304
rect 9404 3120 9456 3126
rect 9402 3088 9404 3097
rect 9456 3088 9458 3097
rect 9402 3023 9458 3032
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 9048 2650 9076 2926
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9416 2310 9444 3023
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 9508 480 9536 5596
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9600 2530 9628 3470
rect 9692 2825 9720 6938
rect 9784 6458 9812 8486
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9784 5098 9812 6394
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9678 2816 9734 2825
rect 9678 2751 9734 2760
rect 9680 2576 9732 2582
rect 9600 2524 9680 2530
rect 9600 2518 9732 2524
rect 9600 2502 9720 2518
rect 9588 2440 9640 2446
rect 9784 2394 9812 3538
rect 9640 2388 9812 2394
rect 9588 2382 9812 2388
rect 9600 2366 9812 2382
rect 9784 2009 9812 2366
rect 9770 2000 9826 2009
rect 9770 1935 9826 1944
rect 9876 1426 9904 10406
rect 9968 4049 9996 10406
rect 10060 10266 10088 11154
rect 10152 11121 10180 11494
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10704 11150 10732 11494
rect 10692 11144 10744 11150
rect 10138 11112 10194 11121
rect 10692 11086 10744 11092
rect 10138 11047 10194 11056
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10704 10266 10732 11086
rect 10782 10840 10838 10849
rect 10782 10775 10838 10784
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10060 8498 10088 9318
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10138 9208 10194 9217
rect 10289 9200 10585 9220
rect 10138 9143 10140 9152
rect 10192 9143 10194 9152
rect 10140 9114 10192 9120
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10152 8430 10180 9114
rect 10704 9042 10732 9454
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 10704 8294 10732 8978
rect 10796 8378 10824 10775
rect 10888 8616 10916 14826
rect 11072 14618 11100 15098
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 11164 13734 11192 14486
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11164 13530 11192 13670
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11242 13288 11298 13297
rect 11242 13223 11298 13232
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11164 11626 11192 12038
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 11256 11354 11284 13223
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11058 11248 11114 11257
rect 11058 11183 11060 11192
rect 11112 11183 11114 11192
rect 11060 11154 11112 11160
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10980 10690 11008 11018
rect 10980 10674 11100 10690
rect 10980 10668 11112 10674
rect 10980 10662 11060 10668
rect 11060 10610 11112 10616
rect 11060 10464 11112 10470
rect 11152 10464 11204 10470
rect 11060 10406 11112 10412
rect 11150 10432 11152 10441
rect 11204 10432 11206 10441
rect 11072 10198 11100 10406
rect 11150 10367 11206 10376
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10980 9518 11008 9998
rect 11256 9722 11284 10066
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 11242 8664 11298 8673
rect 10888 8588 11100 8616
rect 11242 8599 11298 8608
rect 10966 8528 11022 8537
rect 10966 8463 10968 8472
rect 11020 8463 11022 8472
rect 10968 8434 11020 8440
rect 10796 8350 11008 8378
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 7954 10732 8230
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10784 7880 10836 7886
rect 10980 7834 11008 8350
rect 10784 7822 10836 7828
rect 10796 7342 10824 7822
rect 10888 7806 11008 7834
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10152 6934 10180 7142
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10140 6928 10192 6934
rect 10796 6905 10824 7142
rect 10140 6870 10192 6876
rect 10782 6896 10838 6905
rect 10324 6860 10376 6866
rect 10782 6831 10838 6840
rect 10324 6802 10376 6808
rect 10336 6458 10364 6802
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10336 6361 10364 6394
rect 10322 6352 10378 6361
rect 10322 6287 10378 6296
rect 10796 6118 10824 6598
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9954 4040 10010 4049
rect 9954 3975 10010 3984
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9968 3126 9996 3334
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 9968 2417 9996 2450
rect 9954 2408 10010 2417
rect 9954 2343 10010 2352
rect 9864 1420 9916 1426
rect 9864 1362 9916 1368
rect 10060 480 10088 5850
rect 10232 5704 10284 5710
rect 10152 5664 10232 5692
rect 10152 5030 10180 5664
rect 10232 5646 10284 5652
rect 10796 5574 10824 6054
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10796 5166 10824 5510
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10152 4706 10180 4966
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10152 4678 10272 4706
rect 10244 4622 10272 4678
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10152 3738 10180 4558
rect 10244 4010 10272 4558
rect 10704 4185 10732 4966
rect 10796 4486 10824 5102
rect 10888 5001 10916 7806
rect 11072 5914 11100 8588
rect 11256 7342 11284 8599
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10874 4992 10930 5001
rect 10874 4927 10930 4936
rect 10980 4842 11008 5578
rect 10980 4826 11100 4842
rect 10980 4820 11112 4826
rect 10980 4814 11060 4820
rect 11060 4762 11112 4768
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10796 4282 10824 4422
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10690 4176 10746 4185
rect 10690 4111 10746 4120
rect 10704 4078 10732 4111
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10232 4004 10284 4010
rect 10232 3946 10284 3952
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10704 3738 10732 4014
rect 10140 3732 10192 3738
rect 10692 3732 10744 3738
rect 10192 3692 10272 3720
rect 10140 3674 10192 3680
rect 10140 3528 10192 3534
rect 10138 3496 10140 3505
rect 10192 3496 10194 3505
rect 10138 3431 10194 3440
rect 10244 3194 10272 3692
rect 10692 3674 10744 3680
rect 10796 3602 10824 4218
rect 10874 3768 10930 3777
rect 11072 3738 11100 4762
rect 11164 4593 11192 6054
rect 11348 5370 11376 15914
rect 12084 15910 12112 16934
rect 12438 16895 12494 16904
rect 12452 16114 12480 16895
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 11808 14074 11836 15846
rect 12084 15570 12112 15846
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12084 15366 12112 15506
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11900 14929 11928 14962
rect 11886 14920 11942 14929
rect 11886 14855 11942 14864
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11900 14618 11928 14758
rect 12084 14618 12112 15302
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12268 14414 12296 14758
rect 12636 14618 12664 20295
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12820 15366 12848 19110
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 13726 19000 13782 19009
rect 19622 18992 19918 19012
rect 13726 18935 13782 18944
rect 13740 17898 13768 18935
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14094 18184 14150 18193
rect 14094 18119 14150 18128
rect 13740 17870 13952 17898
rect 13174 17368 13230 17377
rect 13174 17303 13230 17312
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12820 14958 12848 15302
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12900 14544 12952 14550
rect 12900 14486 12952 14492
rect 12990 14512 13046 14521
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12806 14376 12862 14385
rect 12268 14074 12296 14350
rect 12806 14311 12862 14320
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11610 12336 11666 12345
rect 11610 12271 11612 12280
rect 11664 12271 11666 12280
rect 11612 12242 11664 12248
rect 11624 11354 11652 12242
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11624 10470 11652 11154
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11624 10169 11652 10406
rect 11610 10160 11666 10169
rect 11610 10095 11666 10104
rect 11716 9636 11744 13738
rect 11888 13728 11940 13734
rect 12440 13728 12492 13734
rect 11888 13670 11940 13676
rect 12438 13696 12440 13705
rect 12492 13696 12494 13705
rect 11900 13530 11928 13670
rect 12438 13631 12494 13640
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11900 12918 11928 13466
rect 12162 13424 12218 13433
rect 12162 13359 12218 13368
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11992 12986 12020 13126
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11900 12714 11928 12854
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11900 12594 11928 12650
rect 11808 12566 11928 12594
rect 11808 12209 11836 12566
rect 11992 12238 12020 12922
rect 12176 12782 12204 13359
rect 12438 13152 12494 13161
rect 12494 13110 12572 13138
rect 12438 13087 12494 13096
rect 12438 12880 12494 12889
rect 12438 12815 12494 12824
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 11980 12232 12032 12238
rect 11794 12200 11850 12209
rect 11980 12174 12032 12180
rect 11794 12135 11850 12144
rect 11992 11898 12020 12174
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12256 10736 12308 10742
rect 12256 10678 12308 10684
rect 12268 10606 12296 10678
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12360 10266 12388 10610
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 11624 9608 11744 9636
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11532 8430 11560 8978
rect 11520 8424 11572 8430
rect 11518 8392 11520 8401
rect 11572 8392 11574 8401
rect 11518 8327 11574 8336
rect 11624 6746 11652 9608
rect 12360 9586 12388 10202
rect 12452 9654 12480 12815
rect 12544 10810 12572 13110
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12728 11694 12756 12242
rect 12716 11688 12768 11694
rect 12714 11656 12716 11665
rect 12768 11656 12770 11665
rect 12714 11591 12770 11600
rect 12820 11354 12848 14311
rect 12912 13870 12940 14486
rect 12990 14447 13046 14456
rect 13004 14414 13032 14447
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 13004 14074 13032 14350
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12912 13025 12940 13806
rect 12898 13016 12954 13025
rect 12898 12951 12954 12960
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 13004 11558 13032 12718
rect 13188 12186 13216 17303
rect 13818 15328 13874 15337
rect 13818 15263 13874 15272
rect 13832 12356 13860 15263
rect 13648 12328 13860 12356
rect 13188 12158 13400 12186
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12820 10606 12848 10950
rect 13096 10674 13124 11086
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12808 10600 12860 10606
rect 12806 10568 12808 10577
rect 12860 10568 12862 10577
rect 12806 10503 12862 10512
rect 13096 10146 13124 10610
rect 13188 10266 13216 11154
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13096 10118 13216 10146
rect 13188 10062 13216 10118
rect 13176 10056 13228 10062
rect 13174 10024 13176 10033
rect 13228 10024 13230 10033
rect 13174 9959 13230 9968
rect 12530 9888 12586 9897
rect 12530 9823 12586 9832
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12164 9512 12216 9518
rect 12162 9480 12164 9489
rect 12216 9480 12218 9489
rect 12162 9415 12218 9424
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12452 9110 12480 9318
rect 12440 9104 12492 9110
rect 12438 9072 12440 9081
rect 12492 9072 12494 9081
rect 12438 9007 12494 9016
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12176 8022 12204 8774
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 12176 7546 12204 7958
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 11794 7440 11850 7449
rect 11794 7375 11850 7384
rect 11532 6718 11652 6746
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11440 6458 11468 6598
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11150 4584 11206 4593
rect 11150 4519 11206 4528
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11150 4040 11206 4049
rect 11150 3975 11206 3984
rect 10874 3703 10930 3712
rect 11060 3732 11112 3738
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10888 3058 10916 3703
rect 11060 3674 11112 3680
rect 10966 3632 11022 3641
rect 10966 3567 11022 3576
rect 10980 3369 11008 3567
rect 10966 3360 11022 3369
rect 10966 3295 11022 3304
rect 10966 3224 11022 3233
rect 10966 3159 11022 3168
rect 10980 3058 11008 3159
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 10140 2848 10192 2854
rect 10138 2816 10140 2825
rect 10192 2816 10194 2825
rect 10690 2816 10746 2825
rect 10138 2751 10194 2760
rect 10289 2748 10585 2768
rect 10690 2751 10746 2760
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10704 2378 10732 2751
rect 10888 2650 10916 2994
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 10692 2372 10744 2378
rect 10692 2314 10744 2320
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10980 1737 11008 2246
rect 10966 1728 11022 1737
rect 10966 1663 11022 1672
rect 10600 1420 10652 1426
rect 10600 1362 10652 1368
rect 10612 480 10640 1362
rect 11164 480 11192 3975
rect 11256 1465 11284 4422
rect 11532 4026 11560 6718
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11624 5710 11652 6598
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11808 5302 11836 7375
rect 12268 6866 12296 8366
rect 12544 7936 12572 9823
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12820 9178 12848 9522
rect 13280 9466 13308 12038
rect 12992 9444 13044 9450
rect 12992 9386 13044 9392
rect 13096 9438 13308 9466
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12360 7908 12572 7936
rect 12360 7562 12388 7908
rect 12530 7848 12586 7857
rect 12530 7783 12532 7792
rect 12584 7783 12586 7792
rect 12532 7754 12584 7760
rect 12360 7534 12480 7562
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11900 5846 11928 6394
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 12268 5778 12296 6802
rect 12452 5914 12480 7534
rect 12636 6066 12664 8502
rect 13004 8498 13032 9386
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13004 8090 13032 8434
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12990 7984 13046 7993
rect 12990 7919 12992 7928
rect 13044 7919 13046 7928
rect 12992 7890 13044 7896
rect 12900 7744 12952 7750
rect 12714 7712 12770 7721
rect 12900 7686 12952 7692
rect 12714 7647 12770 7656
rect 12544 6038 12664 6066
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12544 5817 12572 6038
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12530 5808 12586 5817
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 12348 5772 12400 5778
rect 12400 5732 12480 5760
rect 12530 5743 12586 5752
rect 12348 5714 12400 5720
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11336 4004 11388 4010
rect 11532 3998 11652 4026
rect 11900 4010 11928 4558
rect 11336 3946 11388 3952
rect 11348 3097 11376 3946
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11532 3670 11560 3878
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11532 3126 11560 3606
rect 11520 3120 11572 3126
rect 11334 3088 11390 3097
rect 11334 3023 11390 3032
rect 11518 3088 11520 3097
rect 11572 3088 11574 3097
rect 11518 3023 11574 3032
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 11440 2650 11468 2926
rect 11428 2644 11480 2650
rect 11428 2586 11480 2592
rect 11242 1456 11298 1465
rect 11242 1391 11298 1400
rect 11624 610 11652 3998
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11612 604 11664 610
rect 11612 546 11664 552
rect 11704 604 11756 610
rect 11704 546 11756 552
rect 11716 480 11744 546
rect 12268 480 12296 5306
rect 12452 5234 12480 5732
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12440 4480 12492 4486
rect 12438 4448 12440 4457
rect 12492 4448 12494 4457
rect 12438 4383 12494 4392
rect 12452 4078 12480 4383
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12360 2990 12388 3538
rect 12452 3194 12480 3878
rect 12544 3738 12572 4082
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12544 2990 12572 3674
rect 12636 3602 12664 5850
rect 12728 4758 12756 7647
rect 12912 6866 12940 7686
rect 13004 7546 13032 7890
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12820 6322 12848 6734
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12806 6216 12862 6225
rect 12806 6151 12862 6160
rect 12820 4826 12848 6151
rect 12912 6118 12940 6802
rect 12990 6624 13046 6633
rect 12990 6559 13046 6568
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12716 4752 12768 4758
rect 12716 4694 12768 4700
rect 12728 3738 12756 4694
rect 12806 4448 12862 4457
rect 12806 4383 12862 4392
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12360 2802 12388 2926
rect 12360 2774 12480 2802
rect 12452 2514 12480 2774
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12820 480 12848 4383
rect 12912 3777 12940 4966
rect 13004 4622 13032 6559
rect 13096 6458 13124 9438
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13188 8294 13216 9318
rect 13280 8974 13308 9318
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13188 7206 13216 7822
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 13096 5914 13124 6190
rect 13188 6089 13216 7142
rect 13174 6080 13230 6089
rect 13174 6015 13230 6024
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13280 5370 13308 8910
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 12898 3768 12954 3777
rect 13004 3738 13032 4558
rect 12898 3703 12954 3712
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 13280 3233 13308 4762
rect 13266 3224 13322 3233
rect 13266 3159 13322 3168
rect 13372 480 13400 12158
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13464 10470 13492 11154
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13464 9761 13492 10406
rect 13450 9752 13506 9761
rect 13450 9687 13506 9696
rect 13648 9625 13676 12328
rect 13728 11552 13780 11558
rect 13780 11500 13860 11506
rect 13728 11494 13860 11500
rect 13740 11478 13860 11494
rect 13832 10810 13860 11478
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13740 9654 13768 9862
rect 13728 9648 13780 9654
rect 13634 9616 13690 9625
rect 13728 9590 13780 9596
rect 13634 9551 13690 9560
rect 13740 9178 13768 9590
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13464 8294 13492 9046
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13648 8634 13676 8910
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13464 7410 13492 8230
rect 13556 8022 13584 8298
rect 13544 8016 13596 8022
rect 13544 7958 13596 7964
rect 13556 7410 13584 7958
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13556 7002 13584 7346
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13464 4826 13492 6394
rect 13556 5914 13584 6938
rect 13648 6254 13676 8570
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13464 3942 13492 4626
rect 13740 4434 13768 8774
rect 13924 8634 13952 17870
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 14108 8514 14136 18119
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 14554 12064 14610 12073
rect 14554 11999 14610 12008
rect 14278 10432 14334 10441
rect 14278 10367 14334 10376
rect 13924 8486 14136 8514
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13832 5098 13860 7686
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13740 4406 13860 4434
rect 13726 4312 13782 4321
rect 13726 4247 13782 4256
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13464 3641 13492 3878
rect 13740 3738 13768 4247
rect 13832 4010 13860 4406
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13450 3632 13506 3641
rect 13450 3567 13506 3576
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13648 2514 13676 3334
rect 13740 3194 13768 3674
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13832 2582 13860 2790
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 13636 2508 13688 2514
rect 13636 2450 13688 2456
rect 13924 480 13952 8486
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14016 5370 14044 8366
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14108 7274 14136 7686
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 14108 6662 14136 7210
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14004 5364 14056 5370
rect 14004 5306 14056 5312
rect 14016 5166 14044 5306
rect 14108 5234 14136 6598
rect 14186 6488 14242 6497
rect 14186 6423 14242 6432
rect 14200 5778 14228 6423
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14200 5370 14228 5714
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 14108 4826 14136 5170
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 14200 2922 14228 3334
rect 14188 2916 14240 2922
rect 14188 2858 14240 2864
rect 14200 2650 14228 2858
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14292 2038 14320 10367
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14384 5352 14412 8570
rect 14462 8392 14518 8401
rect 14462 8327 14518 8336
rect 14476 7546 14504 8327
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14568 6254 14596 11999
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 17132 8560 17184 8566
rect 17130 8528 17132 8537
rect 17184 8528 17186 8537
rect 17130 8463 17186 8472
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15672 7274 15700 8230
rect 15764 8022 15792 8366
rect 20180 8265 20208 24103
rect 21008 23866 21036 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 20996 23860 21048 23866
rect 20996 23802 21048 23808
rect 23478 23352 23534 23361
rect 23478 23287 23534 23296
rect 23492 21457 23520 23287
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 23478 21448 23534 21457
rect 23478 21383 23534 21392
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 23478 15600 23534 15609
rect 23478 15535 23534 15544
rect 23492 14482 23520 15535
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 23480 14476 23532 14482
rect 23480 14418 23532 14424
rect 23492 14074 23520 14418
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 24860 14000 24912 14006
rect 23662 13968 23718 13977
rect 23662 13903 23718 13912
rect 23846 13968 23902 13977
rect 24860 13942 24912 13948
rect 23846 13903 23902 13912
rect 23676 13870 23704 13903
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 22284 13388 22336 13394
rect 22284 13330 22336 13336
rect 22296 12782 22324 13330
rect 23480 13184 23532 13190
rect 23480 13126 23532 13132
rect 22284 12776 22336 12782
rect 22282 12744 22284 12753
rect 22336 12744 22338 12753
rect 22282 12679 22338 12688
rect 21732 12300 21784 12306
rect 21732 12242 21784 12248
rect 21744 11830 21772 12242
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21732 11824 21784 11830
rect 21730 11792 21732 11801
rect 21784 11792 21786 11801
rect 21730 11727 21786 11736
rect 21928 11121 21956 12038
rect 21914 11112 21970 11121
rect 21914 11047 21970 11056
rect 20166 8256 20222 8265
rect 19622 8188 19918 8208
rect 20166 8191 20222 8200
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15856 7546 15884 7822
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16500 7290 16528 7346
rect 16500 7274 16620 7290
rect 15660 7268 15712 7274
rect 15660 7210 15712 7216
rect 16488 7268 16620 7274
rect 16540 7262 16620 7268
rect 16488 7210 16540 7216
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 16396 7200 16448 7206
rect 16500 7179 16528 7210
rect 16396 7142 16448 7148
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14844 6458 14872 6802
rect 15672 6798 15700 6938
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15672 6458 15700 6734
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15764 6322 15792 6802
rect 15948 6361 15976 7142
rect 16408 6934 16436 7142
rect 16396 6928 16448 6934
rect 16396 6870 16448 6876
rect 16592 6662 16620 7262
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 17866 6896 17922 6905
rect 17866 6831 17868 6840
rect 17920 6831 17922 6840
rect 17868 6802 17920 6808
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 17880 6458 17908 6802
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 19062 6760 19118 6769
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 15934 6352 15990 6361
rect 15752 6316 15804 6322
rect 15934 6287 15990 6296
rect 16120 6316 16172 6322
rect 15752 6258 15804 6264
rect 16120 6258 16172 6264
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14830 6216 14886 6225
rect 14568 5846 14596 6190
rect 14830 6151 14886 6160
rect 14740 6112 14792 6118
rect 14738 6080 14740 6089
rect 14792 6080 14794 6089
rect 14738 6015 14794 6024
rect 14556 5840 14608 5846
rect 14556 5782 14608 5788
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14646 5400 14702 5409
rect 14384 5324 14596 5352
rect 14646 5335 14702 5344
rect 14464 5092 14516 5098
rect 14464 5034 14516 5040
rect 14476 4826 14504 5034
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14568 4706 14596 5324
rect 14660 4758 14688 5335
rect 14752 5273 14780 5646
rect 14738 5264 14794 5273
rect 14738 5199 14794 5208
rect 14738 5128 14794 5137
rect 14738 5063 14794 5072
rect 14384 4678 14596 4706
rect 14648 4752 14700 4758
rect 14648 4694 14700 4700
rect 14280 2032 14332 2038
rect 14280 1974 14332 1980
rect 14384 480 14412 4678
rect 14752 3670 14780 5063
rect 14844 5030 14872 6151
rect 16132 6118 16160 6258
rect 16580 6248 16632 6254
rect 16578 6216 16580 6225
rect 16632 6216 16634 6225
rect 16578 6151 16634 6160
rect 16854 6216 16910 6225
rect 16854 6151 16856 6160
rect 16908 6151 16910 6160
rect 16856 6122 16908 6128
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 16132 5914 16160 6054
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 16212 5704 16264 5710
rect 15658 5672 15714 5681
rect 15658 5607 15714 5616
rect 15842 5672 15898 5681
rect 16212 5646 16264 5652
rect 15842 5607 15898 5616
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 15488 4486 15516 5510
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15488 4078 15516 4422
rect 15672 4282 15700 5607
rect 15660 4276 15712 4282
rect 15660 4218 15712 4224
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15108 4004 15160 4010
rect 15108 3946 15160 3952
rect 14740 3664 14792 3670
rect 15120 3641 15148 3946
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 14740 3606 14792 3612
rect 15106 3632 15162 3641
rect 14464 3596 14516 3602
rect 15106 3567 15162 3576
rect 14464 3538 14516 3544
rect 14476 3194 14504 3538
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 15304 2446 15332 3878
rect 15488 3398 15516 4014
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15488 2990 15516 3334
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15856 2650 15884 5607
rect 16028 5092 16080 5098
rect 16028 5034 16080 5040
rect 16040 3738 16068 5034
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16132 4593 16160 4966
rect 16118 4584 16174 4593
rect 16118 4519 16174 4528
rect 16224 3738 16252 5646
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 16500 5114 16528 5510
rect 16592 5234 16620 5714
rect 18064 5681 18092 6054
rect 18156 5778 18184 6734
rect 19062 6695 19118 6704
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 18050 5672 18106 5681
rect 18050 5607 18106 5616
rect 18156 5370 18184 5714
rect 18788 5568 18840 5574
rect 18788 5510 18840 5516
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 18052 5160 18104 5166
rect 16500 5086 16620 5114
rect 18052 5102 18104 5108
rect 16592 5030 16620 5086
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16316 3942 16344 4626
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16592 3738 16620 4966
rect 17420 4826 17448 4966
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17958 4312 18014 4321
rect 17958 4247 18014 4256
rect 17406 4176 17462 4185
rect 17406 4111 17408 4120
rect 17460 4111 17462 4120
rect 17408 4082 17460 4088
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16224 3194 16252 3674
rect 16396 3664 16448 3670
rect 16396 3606 16448 3612
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 15474 2544 15530 2553
rect 15474 2479 15530 2488
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 15488 2378 15516 2479
rect 16040 2446 16068 2790
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14924 2032 14976 2038
rect 14924 1974 14976 1980
rect 14936 480 14964 1974
rect 15580 1170 15608 2314
rect 15488 1142 15608 1170
rect 15488 480 15516 1142
rect 16132 1034 16160 3062
rect 16408 3058 16436 3606
rect 16684 3534 16712 3878
rect 17590 3768 17646 3777
rect 17866 3768 17922 3777
rect 17646 3726 17816 3754
rect 17590 3703 17646 3712
rect 17788 3534 17816 3726
rect 17866 3703 17868 3712
rect 17920 3703 17922 3712
rect 17868 3674 17920 3680
rect 16672 3528 16724 3534
rect 17776 3528 17828 3534
rect 16672 3470 16724 3476
rect 16946 3496 17002 3505
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16578 2816 16634 2825
rect 16578 2751 16634 2760
rect 16040 1006 16160 1034
rect 16040 480 16068 1006
rect 16592 480 16620 2751
rect 16684 2650 16712 3470
rect 16946 3431 16948 3440
rect 17000 3431 17002 3440
rect 17774 3496 17776 3505
rect 17828 3496 17830 3505
rect 17774 3431 17830 3440
rect 16948 3402 17000 3408
rect 16960 2990 16988 3402
rect 17682 3224 17738 3233
rect 17682 3159 17738 3168
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 17130 2952 17186 2961
rect 17130 2887 17186 2896
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 17144 480 17172 2887
rect 17696 480 17724 3159
rect 17788 2650 17816 3431
rect 17880 3194 17908 3674
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 17972 2802 18000 4247
rect 18064 3194 18092 5102
rect 18328 5092 18380 5098
rect 18328 5034 18380 5040
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 18248 4457 18276 4626
rect 18234 4448 18290 4457
rect 18234 4383 18290 4392
rect 18248 4282 18276 4383
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 18340 4049 18368 5034
rect 18420 4752 18472 4758
rect 18420 4694 18472 4700
rect 18326 4040 18382 4049
rect 18144 4004 18196 4010
rect 18432 4010 18460 4694
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18524 4185 18552 4558
rect 18510 4176 18566 4185
rect 18510 4111 18566 4120
rect 18326 3975 18382 3984
rect 18420 4004 18472 4010
rect 18144 3946 18196 3952
rect 18420 3946 18472 3952
rect 18156 3534 18184 3946
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18340 3738 18368 3878
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18156 3194 18184 3470
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18340 3058 18368 3674
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18616 3097 18644 3334
rect 18602 3088 18658 3097
rect 18328 3052 18380 3058
rect 18602 3023 18604 3032
rect 18328 2994 18380 3000
rect 18656 3023 18658 3032
rect 18604 2994 18656 3000
rect 18156 2854 18184 2885
rect 18144 2848 18196 2854
rect 17972 2796 18144 2802
rect 17972 2790 18196 2796
rect 17972 2774 18184 2790
rect 18156 2650 18184 2774
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 17866 2136 17922 2145
rect 17866 2071 17922 2080
rect 17880 1737 17908 2071
rect 17866 1728 17922 1737
rect 17866 1663 17922 1672
rect 18050 1728 18106 1737
rect 18050 1663 18106 1672
rect 18064 1465 18092 1663
rect 18340 1601 18368 2450
rect 18512 2440 18564 2446
rect 18510 2408 18512 2417
rect 18564 2408 18566 2417
rect 18510 2343 18566 2352
rect 18326 1592 18382 1601
rect 18326 1527 18382 1536
rect 18050 1456 18106 1465
rect 18050 1391 18106 1400
rect 18234 1456 18290 1465
rect 18234 1391 18290 1400
rect 18248 480 18276 1391
rect 18800 480 18828 5510
rect 19076 3602 19104 6695
rect 19522 6352 19578 6361
rect 19522 6287 19578 6296
rect 19536 6254 19564 6287
rect 19524 6248 19576 6254
rect 19524 6190 19576 6196
rect 22466 6216 22522 6225
rect 20536 6180 20588 6186
rect 22466 6151 22522 6160
rect 20536 6122 20588 6128
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 20258 5808 20314 5817
rect 20258 5743 20314 5752
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 19076 3058 19104 3538
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19352 480 19380 4966
rect 19444 3670 19472 5102
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19524 4684 19576 4690
rect 19524 4626 19576 4632
rect 19536 4593 19564 4626
rect 19522 4584 19578 4593
rect 19522 4519 19578 4528
rect 19536 4282 19564 4519
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 19524 4072 19576 4078
rect 19524 4014 19576 4020
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19536 2553 19564 4014
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19522 2544 19578 2553
rect 19522 2479 19578 2488
rect 19616 2508 19668 2514
rect 19616 2450 19668 2456
rect 19628 1737 19656 2450
rect 19614 1728 19670 1737
rect 19614 1663 19670 1672
rect 19996 1034 20024 3878
rect 20272 2990 20300 5743
rect 20548 5166 20576 6122
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20640 5030 20668 5714
rect 20996 5568 21048 5574
rect 20996 5510 21048 5516
rect 20628 5024 20680 5030
rect 20680 4972 20760 4978
rect 20628 4966 20760 4972
rect 20640 4950 20760 4966
rect 20260 2984 20312 2990
rect 20260 2926 20312 2932
rect 20442 2816 20498 2825
rect 20442 2751 20498 2760
rect 19904 1006 20024 1034
rect 19904 480 19932 1006
rect 20456 480 20484 2751
rect 20732 2582 20760 4950
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 20916 4282 20944 4626
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 20902 4176 20958 4185
rect 20902 4111 20958 4120
rect 20916 4078 20944 4111
rect 20904 4072 20956 4078
rect 20904 4014 20956 4020
rect 20902 3632 20958 3641
rect 20902 3567 20904 3576
rect 20956 3567 20958 3576
rect 20904 3538 20956 3544
rect 20916 2650 20944 3538
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 20720 2576 20772 2582
rect 20720 2518 20772 2524
rect 21008 480 21036 5510
rect 21362 5264 21418 5273
rect 21362 5199 21418 5208
rect 21088 3392 21140 3398
rect 21088 3334 21140 3340
rect 21100 3233 21128 3334
rect 21086 3224 21142 3233
rect 21376 3194 21404 5199
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 21086 3159 21142 3168
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 21376 2990 21404 3130
rect 21364 2984 21416 2990
rect 21364 2926 21416 2932
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 21192 2145 21220 2450
rect 21178 2136 21234 2145
rect 21178 2071 21234 2080
rect 21560 480 21588 4422
rect 22006 4040 22062 4049
rect 22006 3975 22062 3984
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21836 3058 21864 3878
rect 22020 3602 22048 3975
rect 22008 3596 22060 3602
rect 22008 3538 22060 3544
rect 22020 3194 22048 3538
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 21730 2952 21786 2961
rect 21730 2887 21786 2896
rect 21744 2854 21772 2887
rect 21732 2848 21784 2854
rect 21732 2790 21784 2796
rect 22112 480 22140 4422
rect 22204 4146 22232 4558
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 22204 2825 22232 3334
rect 22190 2816 22246 2825
rect 22190 2751 22246 2760
rect 22480 2514 22508 6151
rect 22560 5024 22612 5030
rect 22560 4966 22612 4972
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 22572 1306 22600 4966
rect 23204 4004 23256 4010
rect 23204 3946 23256 3952
rect 22652 2304 22704 2310
rect 22652 2246 22704 2252
rect 22664 1465 22692 2246
rect 22650 1456 22706 1465
rect 22650 1391 22706 1400
rect 22572 1278 22692 1306
rect 22664 480 22692 1278
rect 23216 480 23244 3946
rect 23492 2038 23520 13126
rect 23860 11665 23888 13903
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 23846 11656 23902 11665
rect 23846 11591 23902 11600
rect 23570 11112 23626 11121
rect 23570 11047 23626 11056
rect 23480 2032 23532 2038
rect 23480 1974 23532 1980
rect 23584 610 23612 11047
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24766 8256 24822 8265
rect 24766 8191 24822 8200
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 23940 3596 23992 3602
rect 23940 3538 23992 3544
rect 23952 2854 23980 3538
rect 24124 3392 24176 3398
rect 24124 3334 24176 3340
rect 24136 3097 24164 3334
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24780 3194 24808 8191
rect 24768 3188 24820 3194
rect 24768 3130 24820 3136
rect 24122 3088 24178 3097
rect 24122 3023 24178 3032
rect 23940 2848 23992 2854
rect 23940 2790 23992 2796
rect 24766 2816 24822 2825
rect 23952 2009 23980 2790
rect 24766 2751 24822 2760
rect 24780 2650 24808 2751
rect 24768 2644 24820 2650
rect 24768 2586 24820 2592
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24308 2032 24360 2038
rect 23938 2000 23994 2009
rect 24308 1974 24360 1980
rect 23938 1935 23994 1944
rect 23572 604 23624 610
rect 23572 546 23624 552
rect 23756 604 23808 610
rect 23756 546 23808 552
rect 23768 480 23796 546
rect 24320 480 24348 1974
rect 24872 480 24900 13942
rect 24964 610 24992 14214
rect 26514 3632 26570 3641
rect 26514 3567 26570 3576
rect 25962 3088 26018 3097
rect 25962 3023 26018 3032
rect 25226 2952 25282 2961
rect 25226 2887 25228 2896
rect 25280 2887 25282 2896
rect 25228 2858 25280 2864
rect 24952 604 25004 610
rect 24952 546 25004 552
rect 25412 604 25464 610
rect 25412 546 25464 552
rect 25424 480 25452 546
rect 25976 480 26004 3023
rect 26528 480 26556 3567
rect 27066 2952 27122 2961
rect 27066 2887 27122 2896
rect 27080 480 27108 2887
rect 27618 2816 27674 2825
rect 27618 2751 27674 2760
rect 27632 480 27660 2751
rect 2778 368 2834 377
rect 2778 303 2834 312
rect 2870 0 2926 480
rect 3422 0 3478 480
rect 3974 0 4030 480
rect 4526 0 4582 480
rect 5078 0 5134 480
rect 5630 0 5686 480
rect 6182 0 6238 480
rect 6734 0 6790 480
rect 7286 0 7342 480
rect 7838 0 7894 480
rect 8390 0 8446 480
rect 8942 0 8998 480
rect 9494 0 9550 480
rect 10046 0 10102 480
rect 10598 0 10654 480
rect 11150 0 11206 480
rect 11702 0 11758 480
rect 12254 0 12310 480
rect 12806 0 12862 480
rect 13358 0 13414 480
rect 13910 0 13966 480
rect 14370 0 14426 480
rect 14922 0 14978 480
rect 15474 0 15530 480
rect 16026 0 16082 480
rect 16578 0 16634 480
rect 17130 0 17186 480
rect 17682 0 17738 480
rect 18234 0 18290 480
rect 18786 0 18842 480
rect 19338 0 19394 480
rect 19890 0 19946 480
rect 20442 0 20498 480
rect 20994 0 21050 480
rect 21546 0 21602 480
rect 22098 0 22154 480
rect 22650 0 22706 480
rect 23202 0 23258 480
rect 23754 0 23810 480
rect 24306 0 24362 480
rect 24858 0 24914 480
rect 25410 0 25466 480
rect 25962 0 26018 480
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 2410 27648 2466 27704
rect 1582 24792 1638 24848
rect 1582 21392 1638 21448
rect 1950 21392 2006 21448
rect 1950 20460 2006 20496
rect 1950 20440 1952 20460
rect 1952 20440 2004 20460
rect 2004 20440 2006 20460
rect 1398 18400 1454 18456
rect 1582 19252 1584 19272
rect 1584 19252 1636 19272
rect 1636 19252 1638 19272
rect 1582 19216 1638 19252
rect 1582 18264 1638 18320
rect 1674 18128 1730 18184
rect 1490 15988 1492 16008
rect 1492 15988 1544 16008
rect 1544 15988 1546 16008
rect 1490 15952 1546 15988
rect 1306 12280 1362 12336
rect 1490 9696 1546 9752
rect 662 2760 718 2816
rect 2134 20032 2190 20088
rect 2134 19352 2190 19408
rect 4066 27104 4122 27160
rect 4066 26580 4122 26616
rect 4066 26560 4068 26580
rect 4068 26560 4120 26580
rect 4120 26560 4122 26580
rect 3790 26016 3846 26072
rect 2686 25336 2742 25392
rect 4066 24248 4122 24304
rect 2502 22380 2504 22400
rect 2504 22380 2556 22400
rect 2556 22380 2558 22400
rect 2502 22344 2558 22380
rect 4066 23296 4122 23352
rect 4250 22480 4306 22536
rect 2870 22072 2926 22128
rect 3146 21936 3202 21992
rect 2870 19624 2926 19680
rect 3514 19216 3570 19272
rect 3054 19080 3110 19136
rect 2594 18944 2650 19000
rect 2870 18944 2926 19000
rect 2226 18536 2282 18592
rect 1674 12416 1730 12472
rect 1950 8744 2006 8800
rect 1582 6060 1584 6080
rect 1584 6060 1636 6080
rect 1636 6060 1638 6080
rect 1582 6024 1638 6060
rect 1858 4664 1914 4720
rect 2502 17720 2558 17776
rect 2502 17176 2558 17232
rect 2962 18264 3018 18320
rect 2686 15000 2742 15056
rect 3238 16224 3294 16280
rect 5262 23160 5318 23216
rect 4710 22208 4766 22264
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 7010 24112 7066 24168
rect 20166 24112 20222 24168
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 7470 23704 7526 23760
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 8298 23316 8354 23352
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 8298 23296 8300 23316
rect 8300 23296 8352 23316
rect 8352 23296 8354 23316
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 4158 20848 4214 20904
rect 5078 21428 5080 21448
rect 5080 21428 5132 21448
rect 5132 21428 5134 21448
rect 5078 21392 5134 21428
rect 8298 22208 8354 22264
rect 7838 21292 7840 21312
rect 7840 21292 7892 21312
rect 7892 21292 7894 21312
rect 7838 21256 7894 21292
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5538 20440 5594 20496
rect 5722 20304 5778 20360
rect 5078 20204 5080 20224
rect 5080 20204 5132 20224
rect 5132 20204 5134 20224
rect 5078 20168 5134 20204
rect 5170 20032 5226 20088
rect 3698 18284 3754 18320
rect 3698 18264 3700 18284
rect 3700 18264 3752 18284
rect 3752 18264 3754 18284
rect 4066 18128 4122 18184
rect 5078 18400 5134 18456
rect 4250 17992 4306 18048
rect 3882 17448 3938 17504
rect 3698 16768 3754 16824
rect 3422 14592 3478 14648
rect 2594 11464 2650 11520
rect 2410 10124 2466 10160
rect 2410 10104 2412 10124
rect 2412 10104 2464 10124
rect 2464 10104 2466 10124
rect 2502 9696 2558 9752
rect 2226 7248 2282 7304
rect 3146 12280 3202 12336
rect 2962 11736 3018 11792
rect 3422 13504 3478 13560
rect 2134 5616 2190 5672
rect 2042 4140 2098 4176
rect 2042 4120 2044 4140
rect 2044 4120 2096 4140
rect 2096 4120 2098 4140
rect 1950 3712 2006 3768
rect 2502 6704 2558 6760
rect 2134 2372 2190 2408
rect 2134 2352 2136 2372
rect 2136 2352 2188 2372
rect 2188 2352 2190 2372
rect 2502 2644 2558 2680
rect 2502 2624 2504 2644
rect 2504 2624 2556 2644
rect 2556 2624 2558 2644
rect 3790 15136 3846 15192
rect 3790 13912 3846 13968
rect 3974 16632 4030 16688
rect 3974 15680 4030 15736
rect 4250 15952 4306 16008
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5630 18808 5686 18864
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 7102 19352 7158 19408
rect 6090 18264 6146 18320
rect 6274 18284 6330 18320
rect 6274 18264 6276 18284
rect 6276 18264 6328 18284
rect 6328 18264 6330 18284
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5998 17312 6054 17368
rect 5170 16632 5226 16688
rect 5814 16652 5870 16688
rect 5814 16632 5816 16652
rect 5816 16632 5868 16652
rect 5868 16632 5870 16652
rect 4618 15000 4674 15056
rect 3882 13268 3884 13288
rect 3884 13268 3936 13288
rect 3936 13268 3938 13288
rect 3882 13232 3938 13268
rect 3882 11328 3938 11384
rect 3606 11056 3662 11112
rect 3330 5480 3386 5536
rect 2870 4936 2926 4992
rect 3514 7248 3570 7304
rect 3698 9968 3754 10024
rect 3882 9424 3938 9480
rect 3698 8472 3754 8528
rect 3606 6840 3662 6896
rect 3698 5108 3700 5128
rect 3700 5108 3752 5128
rect 3752 5108 3754 5128
rect 3698 5072 3754 5108
rect 3606 4800 3662 4856
rect 3422 2488 3478 2544
rect 2962 2352 3018 2408
rect 3698 4256 3754 4312
rect 3606 1808 3662 1864
rect 4158 12280 4214 12336
rect 4066 9016 4122 9072
rect 4066 8472 4122 8528
rect 4710 14356 4712 14376
rect 4712 14356 4764 14376
rect 4764 14356 4766 14376
rect 4710 14320 4766 14356
rect 4434 10512 4490 10568
rect 4342 8472 4398 8528
rect 4802 12280 4858 12336
rect 5170 14592 5226 14648
rect 5078 12416 5134 12472
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5630 15000 5686 15056
rect 5630 14764 5632 14784
rect 5632 14764 5684 14784
rect 5684 14764 5686 14784
rect 5630 14728 5686 14764
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 4986 10240 5042 10296
rect 4066 7112 4122 7168
rect 3974 5480 4030 5536
rect 3882 5072 3938 5128
rect 3790 1536 3846 1592
rect 3974 4800 4030 4856
rect 3974 3712 4030 3768
rect 4526 6704 4582 6760
rect 4250 3168 4306 3224
rect 4434 3712 4490 3768
rect 4618 6568 4674 6624
rect 4710 5344 4766 5400
rect 5354 9832 5410 9888
rect 5170 8336 5226 8392
rect 5078 8064 5134 8120
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5538 12280 5594 12336
rect 6734 14592 6790 14648
rect 6182 13776 6238 13832
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6458 13368 6514 13424
rect 6274 13232 6330 13288
rect 6366 12552 6422 12608
rect 6182 11736 6238 11792
rect 6090 11328 6146 11384
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 6366 11464 6422 11520
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5998 9696 6054 9752
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 6182 9016 6238 9072
rect 5170 6976 5226 7032
rect 5078 5616 5134 5672
rect 4986 4120 5042 4176
rect 4894 1944 4950 2000
rect 5630 7792 5686 7848
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 6090 5752 6146 5808
rect 6090 4972 6092 4992
rect 6092 4972 6144 4992
rect 6144 4972 6146 4992
rect 6090 4936 6146 4972
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5998 2644 6054 2680
rect 5998 2624 6000 2644
rect 6000 2624 6052 2644
rect 6052 2624 6054 2644
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 5170 1536 5226 1592
rect 6366 9288 6422 9344
rect 6458 9152 6514 9208
rect 6826 12960 6882 13016
rect 7102 12280 7158 12336
rect 6366 6840 6422 6896
rect 6366 4392 6422 4448
rect 6366 2388 6368 2408
rect 6368 2388 6420 2408
rect 6420 2388 6422 2408
rect 6366 2352 6422 2388
rect 6550 8064 6606 8120
rect 6550 4664 6606 4720
rect 7010 11600 7066 11656
rect 6826 10104 6882 10160
rect 6734 9988 6790 10024
rect 6734 9968 6736 9988
rect 6736 9968 6788 9988
rect 6788 9968 6790 9988
rect 6918 9968 6974 10024
rect 7286 15700 7342 15736
rect 7286 15680 7288 15700
rect 7288 15680 7340 15700
rect 7340 15680 7342 15700
rect 7010 9832 7066 9888
rect 7102 9424 7158 9480
rect 7102 8336 7158 8392
rect 6826 6452 6882 6488
rect 6826 6432 6828 6452
rect 6828 6432 6880 6452
rect 6880 6432 6882 6452
rect 7010 5072 7066 5128
rect 7654 18028 7656 18048
rect 7656 18028 7708 18048
rect 7708 18028 7710 18048
rect 7654 17992 7710 18028
rect 7562 14728 7618 14784
rect 7378 12588 7380 12608
rect 7380 12588 7432 12608
rect 7432 12588 7434 12608
rect 7378 12552 7434 12588
rect 7378 9560 7434 9616
rect 7470 7792 7526 7848
rect 7378 6316 7434 6352
rect 7378 6296 7380 6316
rect 7380 6296 7432 6316
rect 7432 6296 7434 6316
rect 7010 4256 7066 4312
rect 6458 856 6514 912
rect 7194 3596 7250 3632
rect 7194 3576 7196 3596
rect 7196 3576 7248 3596
rect 7248 3576 7250 3596
rect 7010 2796 7012 2816
rect 7012 2796 7064 2816
rect 7064 2796 7066 2816
rect 7654 14048 7710 14104
rect 7838 13812 7840 13832
rect 7840 13812 7892 13832
rect 7892 13812 7894 13832
rect 7838 13776 7894 13812
rect 8022 18672 8078 18728
rect 8390 18164 8392 18184
rect 8392 18164 8444 18184
rect 8444 18164 8446 18184
rect 8390 18128 8446 18164
rect 7930 11872 7986 11928
rect 9494 17992 9550 18048
rect 8206 16668 8208 16688
rect 8208 16668 8260 16688
rect 8260 16668 8262 16688
rect 8206 16632 8262 16668
rect 8390 15308 8392 15328
rect 8392 15308 8444 15328
rect 8444 15308 8446 15328
rect 8390 15272 8446 15308
rect 8666 14884 8722 14920
rect 8666 14864 8668 14884
rect 8668 14864 8720 14884
rect 8720 14864 8722 14884
rect 8758 14612 8814 14648
rect 8758 14592 8760 14612
rect 8760 14592 8812 14612
rect 8812 14592 8814 14612
rect 9126 14492 9128 14512
rect 9128 14492 9180 14512
rect 9180 14492 9182 14512
rect 9126 14456 9182 14492
rect 8298 14048 8354 14104
rect 7654 10920 7710 10976
rect 7654 10376 7710 10432
rect 8574 12860 8576 12880
rect 8576 12860 8628 12880
rect 8628 12860 8630 12880
rect 8574 12824 8630 12860
rect 8022 11056 8078 11112
rect 8206 11192 8262 11248
rect 8666 11056 8722 11112
rect 8850 10784 8906 10840
rect 8390 10240 8446 10296
rect 8298 9288 8354 9344
rect 8298 8880 8354 8936
rect 7746 6724 7802 6760
rect 7746 6704 7748 6724
rect 7748 6704 7800 6724
rect 7800 6704 7802 6724
rect 7838 5616 7894 5672
rect 8298 8492 8354 8528
rect 8298 8472 8300 8492
rect 8300 8472 8352 8492
rect 8352 8472 8354 8492
rect 8206 6976 8262 7032
rect 8022 4664 8078 4720
rect 8114 3732 8170 3768
rect 8114 3712 8116 3732
rect 8116 3712 8168 3732
rect 8168 3712 8170 3732
rect 7010 2760 7066 2796
rect 8850 9324 8852 9344
rect 8852 9324 8904 9344
rect 8904 9324 8906 9344
rect 8850 9288 8906 9324
rect 8850 8628 8906 8664
rect 8850 8608 8852 8628
rect 8852 8608 8904 8628
rect 8904 8608 8906 8628
rect 9954 22344 10010 22400
rect 9770 22072 9826 22128
rect 9678 21256 9734 21312
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 10690 21392 10746 21448
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 12622 20304 12678 20360
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10966 18944 11022 19000
rect 11242 18808 11298 18864
rect 10138 18708 10140 18728
rect 10140 18708 10192 18728
rect 10192 18708 10194 18728
rect 10138 18672 10194 18708
rect 10690 18300 10692 18320
rect 10692 18300 10744 18320
rect 10744 18300 10746 18320
rect 10690 18264 10746 18300
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10046 17720 10102 17776
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10782 16904 10838 16960
rect 11242 16632 11298 16688
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 9218 13368 9274 13424
rect 9126 12180 9128 12200
rect 9128 12180 9180 12200
rect 9180 12180 9182 12200
rect 9126 12144 9182 12180
rect 9494 8336 9550 8392
rect 9494 7520 9550 7576
rect 9402 6568 9458 6624
rect 9310 6160 9366 6216
rect 9770 15000 9826 15056
rect 9954 14048 10010 14104
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10138 13776 10194 13832
rect 10046 13504 10102 13560
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10782 13640 10838 13696
rect 10138 12688 10194 12744
rect 10322 12688 10378 12744
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10138 12008 10194 12064
rect 10046 11872 10102 11928
rect 9678 10920 9734 10976
rect 9126 3304 9182 3360
rect 9402 3068 9404 3088
rect 9404 3068 9456 3088
rect 9456 3068 9458 3088
rect 9402 3032 9458 3068
rect 9678 2760 9734 2816
rect 9770 1944 9826 2000
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10138 11056 10194 11112
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10782 10784 10838 10840
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10138 9172 10194 9208
rect 10138 9152 10140 9172
rect 10140 9152 10192 9172
rect 10192 9152 10194 9172
rect 11242 13232 11298 13288
rect 11058 11212 11114 11248
rect 11058 11192 11060 11212
rect 11060 11192 11112 11212
rect 11112 11192 11114 11212
rect 11150 10412 11152 10432
rect 11152 10412 11204 10432
rect 11204 10412 11206 10432
rect 11150 10376 11206 10412
rect 11242 8608 11298 8664
rect 10966 8492 11022 8528
rect 10966 8472 10968 8492
rect 10968 8472 11020 8492
rect 11020 8472 11022 8492
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10782 6840 10838 6896
rect 10322 6296 10378 6352
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 9954 3984 10010 4040
rect 9954 2352 10010 2408
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10874 4936 10930 4992
rect 10690 4120 10746 4176
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10138 3476 10140 3496
rect 10140 3476 10192 3496
rect 10192 3476 10194 3496
rect 10138 3440 10194 3476
rect 10874 3712 10930 3768
rect 12438 16904 12494 16960
rect 11886 14864 11942 14920
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 13726 18944 13782 19000
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14094 18128 14150 18184
rect 13174 17312 13230 17368
rect 12806 14320 12862 14376
rect 11610 12300 11666 12336
rect 11610 12280 11612 12300
rect 11612 12280 11664 12300
rect 11664 12280 11666 12300
rect 11610 10104 11666 10160
rect 12438 13676 12440 13696
rect 12440 13676 12492 13696
rect 12492 13676 12494 13696
rect 12438 13640 12494 13676
rect 12162 13368 12218 13424
rect 12438 13096 12494 13152
rect 12438 12824 12494 12880
rect 11794 12144 11850 12200
rect 11518 8372 11520 8392
rect 11520 8372 11572 8392
rect 11572 8372 11574 8392
rect 11518 8336 11574 8372
rect 12714 11636 12716 11656
rect 12716 11636 12768 11656
rect 12768 11636 12770 11656
rect 12714 11600 12770 11636
rect 12990 14456 13046 14512
rect 12898 12960 12954 13016
rect 13818 15272 13874 15328
rect 12806 10548 12808 10568
rect 12808 10548 12860 10568
rect 12860 10548 12862 10568
rect 12806 10512 12862 10548
rect 13174 10004 13176 10024
rect 13176 10004 13228 10024
rect 13228 10004 13230 10024
rect 13174 9968 13230 10004
rect 12530 9832 12586 9888
rect 12162 9460 12164 9480
rect 12164 9460 12216 9480
rect 12216 9460 12218 9480
rect 12162 9424 12218 9460
rect 12438 9052 12440 9072
rect 12440 9052 12492 9072
rect 12492 9052 12494 9072
rect 12438 9016 12494 9052
rect 11794 7384 11850 7440
rect 11150 4528 11206 4584
rect 11150 3984 11206 4040
rect 10966 3576 11022 3632
rect 10966 3304 11022 3360
rect 10966 3168 11022 3224
rect 10138 2796 10140 2816
rect 10140 2796 10192 2816
rect 10192 2796 10194 2816
rect 10138 2760 10194 2796
rect 10690 2760 10746 2816
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10966 1672 11022 1728
rect 12530 7812 12586 7848
rect 12530 7792 12532 7812
rect 12532 7792 12584 7812
rect 12584 7792 12586 7812
rect 12990 7948 13046 7984
rect 12990 7928 12992 7948
rect 12992 7928 13044 7948
rect 13044 7928 13046 7948
rect 12714 7656 12770 7712
rect 12530 5752 12586 5808
rect 11334 3032 11390 3088
rect 11518 3068 11520 3088
rect 11520 3068 11572 3088
rect 11572 3068 11574 3088
rect 11518 3032 11574 3068
rect 11242 1400 11298 1456
rect 12438 4428 12440 4448
rect 12440 4428 12492 4448
rect 12492 4428 12494 4448
rect 12438 4392 12494 4428
rect 12806 6160 12862 6216
rect 12990 6568 13046 6624
rect 12806 4392 12862 4448
rect 13174 6024 13230 6080
rect 12898 3712 12954 3768
rect 13266 3168 13322 3224
rect 13450 9696 13506 9752
rect 13634 9560 13690 9616
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 14554 12008 14610 12064
rect 14278 10376 14334 10432
rect 13726 4256 13782 4312
rect 13450 3576 13506 3632
rect 14186 6432 14242 6488
rect 14462 8336 14518 8392
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 17130 8508 17132 8528
rect 17132 8508 17184 8528
rect 17184 8508 17186 8528
rect 17130 8472 17186 8508
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 23478 23296 23534 23352
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 23478 21392 23534 21448
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 23478 15544 23534 15600
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 23662 13912 23718 13968
rect 23846 13912 23902 13968
rect 22282 12724 22284 12744
rect 22284 12724 22336 12744
rect 22336 12724 22338 12744
rect 22282 12688 22338 12724
rect 21730 11772 21732 11792
rect 21732 11772 21784 11792
rect 21784 11772 21786 11792
rect 21730 11736 21786 11772
rect 21914 11056 21970 11112
rect 20166 8200 20222 8256
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 17866 6860 17922 6896
rect 17866 6840 17868 6860
rect 17868 6840 17920 6860
rect 17920 6840 17922 6860
rect 15934 6296 15990 6352
rect 14830 6160 14886 6216
rect 14738 6060 14740 6080
rect 14740 6060 14792 6080
rect 14792 6060 14794 6080
rect 14738 6024 14794 6060
rect 14646 5344 14702 5400
rect 14738 5208 14794 5264
rect 14738 5072 14794 5128
rect 16578 6196 16580 6216
rect 16580 6196 16632 6216
rect 16632 6196 16634 6216
rect 16578 6160 16634 6196
rect 16854 6180 16910 6216
rect 16854 6160 16856 6180
rect 16856 6160 16908 6180
rect 16908 6160 16910 6180
rect 15658 5616 15714 5672
rect 15842 5616 15898 5672
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15106 3576 15162 3632
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 16118 4528 16174 4584
rect 19062 6704 19118 6760
rect 18050 5616 18106 5672
rect 17958 4256 18014 4312
rect 17406 4140 17462 4176
rect 17406 4120 17408 4140
rect 17408 4120 17460 4140
rect 17460 4120 17462 4140
rect 15474 2488 15530 2544
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 17590 3712 17646 3768
rect 17866 3732 17922 3768
rect 17866 3712 17868 3732
rect 17868 3712 17920 3732
rect 17920 3712 17922 3732
rect 16578 2760 16634 2816
rect 16946 3460 17002 3496
rect 16946 3440 16948 3460
rect 16948 3440 17000 3460
rect 17000 3440 17002 3460
rect 17774 3476 17776 3496
rect 17776 3476 17828 3496
rect 17828 3476 17830 3496
rect 17774 3440 17830 3476
rect 17682 3168 17738 3224
rect 17130 2896 17186 2952
rect 18234 4392 18290 4448
rect 18326 3984 18382 4040
rect 18510 4120 18566 4176
rect 18602 3052 18658 3088
rect 18602 3032 18604 3052
rect 18604 3032 18656 3052
rect 18656 3032 18658 3052
rect 17866 2080 17922 2136
rect 17866 1672 17922 1728
rect 18050 1672 18106 1728
rect 18510 2388 18512 2408
rect 18512 2388 18564 2408
rect 18564 2388 18566 2408
rect 18510 2352 18566 2388
rect 18326 1536 18382 1592
rect 18050 1400 18106 1456
rect 18234 1400 18290 1456
rect 19522 6296 19578 6352
rect 22466 6160 22522 6216
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 20258 5752 20314 5808
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19522 4528 19578 4584
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 19522 2488 19578 2544
rect 19614 1672 19670 1728
rect 20442 2760 20498 2816
rect 20902 4120 20958 4176
rect 20902 3596 20958 3632
rect 20902 3576 20904 3596
rect 20904 3576 20956 3596
rect 20956 3576 20958 3596
rect 21362 5208 21418 5264
rect 21086 3168 21142 3224
rect 21178 2080 21234 2136
rect 22006 3984 22062 4040
rect 21730 2896 21786 2952
rect 22190 2760 22246 2816
rect 22650 1400 22706 1456
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 23846 11600 23902 11656
rect 23570 11056 23626 11112
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24766 8200 24822 8256
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24122 3032 24178 3088
rect 24766 2760 24822 2816
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 23938 1944 23994 2000
rect 26514 3576 26570 3632
rect 25962 3032 26018 3088
rect 25226 2916 25282 2952
rect 25226 2896 25228 2916
rect 25228 2896 25280 2916
rect 25280 2896 25282 2916
rect 27066 2896 27122 2952
rect 27618 2760 27674 2816
rect 2778 312 2834 368
<< metal3 >>
rect 0 27706 480 27736
rect 2405 27706 2471 27709
rect 0 27704 2471 27706
rect 0 27648 2410 27704
rect 2466 27648 2471 27704
rect 0 27646 2471 27648
rect 0 27616 480 27646
rect 2405 27643 2471 27646
rect 0 27162 480 27192
rect 4061 27162 4127 27165
rect 0 27160 4127 27162
rect 0 27104 4066 27160
rect 4122 27104 4127 27160
rect 0 27102 4127 27104
rect 0 27072 480 27102
rect 4061 27099 4127 27102
rect 0 26618 480 26648
rect 4061 26618 4127 26621
rect 0 26616 4127 26618
rect 0 26560 4066 26616
rect 4122 26560 4127 26616
rect 0 26558 4127 26560
rect 0 26528 480 26558
rect 4061 26555 4127 26558
rect 0 26074 480 26104
rect 3785 26074 3851 26077
rect 0 26072 3851 26074
rect 0 26016 3790 26072
rect 3846 26016 3851 26072
rect 0 26014 3851 26016
rect 0 25984 480 26014
rect 3785 26011 3851 26014
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25394 480 25424
rect 2681 25394 2747 25397
rect 0 25392 2747 25394
rect 0 25336 2686 25392
rect 2742 25336 2747 25392
rect 0 25334 2747 25336
rect 0 25304 480 25334
rect 2681 25331 2747 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24850 480 24880
rect 1577 24850 1643 24853
rect 0 24848 1643 24850
rect 0 24792 1582 24848
rect 1638 24792 1643 24848
rect 0 24790 1643 24792
rect 0 24760 480 24790
rect 1577 24787 1643 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 0 24306 480 24336
rect 4061 24306 4127 24309
rect 0 24304 4127 24306
rect 0 24248 4066 24304
rect 4122 24248 4127 24304
rect 0 24246 4127 24248
rect 0 24216 480 24246
rect 4061 24243 4127 24246
rect 7005 24170 7071 24173
rect 20161 24170 20227 24173
rect 7005 24168 20227 24170
rect 7005 24112 7010 24168
rect 7066 24112 20166 24168
rect 20222 24112 20227 24168
rect 7005 24110 20227 24112
rect 7005 24107 7071 24110
rect 20161 24107 20227 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 0 23762 480 23792
rect 7465 23762 7531 23765
rect 0 23760 7531 23762
rect 0 23704 7470 23760
rect 7526 23704 7531 23760
rect 0 23702 7531 23704
rect 0 23672 480 23702
rect 7465 23699 7531 23702
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 4061 23354 4127 23357
rect 8293 23354 8359 23357
rect 4061 23352 8359 23354
rect 4061 23296 4066 23352
rect 4122 23296 8298 23352
rect 8354 23296 8359 23352
rect 4061 23294 8359 23296
rect 4061 23291 4127 23294
rect 8293 23291 8359 23294
rect 23473 23354 23539 23357
rect 27520 23354 28000 23384
rect 23473 23352 28000 23354
rect 23473 23296 23478 23352
rect 23534 23296 28000 23352
rect 23473 23294 28000 23296
rect 23473 23291 23539 23294
rect 27520 23264 28000 23294
rect 0 23218 480 23248
rect 5257 23218 5323 23221
rect 0 23216 5323 23218
rect 0 23160 5262 23216
rect 5318 23160 5323 23216
rect 0 23158 5323 23160
rect 0 23128 480 23158
rect 5257 23155 5323 23158
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 0 22538 480 22568
rect 4245 22538 4311 22541
rect 0 22536 4311 22538
rect 0 22480 4250 22536
rect 4306 22480 4311 22536
rect 0 22478 4311 22480
rect 0 22448 480 22478
rect 4245 22475 4311 22478
rect 2497 22402 2563 22405
rect 9949 22402 10015 22405
rect 2497 22400 10015 22402
rect 2497 22344 2502 22400
rect 2558 22344 9954 22400
rect 10010 22344 10015 22400
rect 2497 22342 10015 22344
rect 2497 22339 2563 22342
rect 9949 22339 10015 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 4705 22266 4771 22269
rect 8293 22266 8359 22269
rect 4705 22264 8359 22266
rect 4705 22208 4710 22264
rect 4766 22208 8298 22264
rect 8354 22208 8359 22264
rect 4705 22206 8359 22208
rect 4705 22203 4771 22206
rect 8293 22203 8359 22206
rect 2865 22130 2931 22133
rect 9765 22130 9831 22133
rect 2865 22128 9831 22130
rect 2865 22072 2870 22128
rect 2926 22072 9770 22128
rect 9826 22072 9831 22128
rect 2865 22070 9831 22072
rect 2865 22067 2931 22070
rect 9765 22067 9831 22070
rect 0 21994 480 22024
rect 3141 21994 3207 21997
rect 0 21992 3207 21994
rect 0 21936 3146 21992
rect 3202 21936 3207 21992
rect 0 21934 3207 21936
rect 0 21904 480 21934
rect 3141 21931 3207 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 0 21450 480 21480
rect 1577 21450 1643 21453
rect 0 21448 1643 21450
rect 0 21392 1582 21448
rect 1638 21392 1643 21448
rect 0 21390 1643 21392
rect 0 21360 480 21390
rect 1577 21387 1643 21390
rect 1945 21450 2011 21453
rect 5073 21450 5139 21453
rect 1945 21448 5139 21450
rect 1945 21392 1950 21448
rect 2006 21392 5078 21448
rect 5134 21392 5139 21448
rect 1945 21390 5139 21392
rect 1945 21387 2011 21390
rect 5073 21387 5139 21390
rect 10685 21450 10751 21453
rect 23473 21450 23539 21453
rect 10685 21448 23539 21450
rect 10685 21392 10690 21448
rect 10746 21392 23478 21448
rect 23534 21392 23539 21448
rect 10685 21390 23539 21392
rect 10685 21387 10751 21390
rect 23473 21387 23539 21390
rect 7833 21314 7899 21317
rect 9673 21314 9739 21317
rect 7833 21312 9739 21314
rect 7833 21256 7838 21312
rect 7894 21256 9678 21312
rect 9734 21256 9739 21312
rect 7833 21254 9739 21256
rect 7833 21251 7899 21254
rect 9673 21251 9739 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 0 20906 480 20936
rect 4153 20906 4219 20909
rect 0 20904 4219 20906
rect 0 20848 4158 20904
rect 4214 20848 4219 20904
rect 0 20846 4219 20848
rect 0 20816 480 20846
rect 4153 20843 4219 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 1945 20498 2011 20501
rect 5533 20498 5599 20501
rect 1945 20496 5599 20498
rect 1945 20440 1950 20496
rect 2006 20440 5538 20496
rect 5594 20440 5599 20496
rect 1945 20438 5599 20440
rect 1945 20435 2011 20438
rect 5533 20435 5599 20438
rect 0 20362 480 20392
rect 5717 20362 5783 20365
rect 12617 20362 12683 20365
rect 0 20360 5783 20362
rect 0 20304 5722 20360
rect 5778 20304 5783 20360
rect 0 20302 5783 20304
rect 0 20272 480 20302
rect 5717 20299 5783 20302
rect 5950 20360 12683 20362
rect 5950 20304 12622 20360
rect 12678 20304 12683 20360
rect 5950 20302 12683 20304
rect 5073 20226 5139 20229
rect 5950 20226 6010 20302
rect 12617 20299 12683 20302
rect 5073 20224 6010 20226
rect 5073 20168 5078 20224
rect 5134 20168 6010 20224
rect 5073 20166 6010 20168
rect 5073 20163 5139 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 2129 20090 2195 20093
rect 5165 20090 5231 20093
rect 2129 20088 5231 20090
rect 2129 20032 2134 20088
rect 2190 20032 5170 20088
rect 5226 20032 5231 20088
rect 2129 20030 5231 20032
rect 2129 20027 2195 20030
rect 5165 20027 5231 20030
rect 0 19682 480 19712
rect 2865 19682 2931 19685
rect 0 19680 2931 19682
rect 0 19624 2870 19680
rect 2926 19624 2931 19680
rect 0 19622 2931 19624
rect 0 19592 480 19622
rect 2865 19619 2931 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 2129 19410 2195 19413
rect 7097 19410 7163 19413
rect 2129 19408 7163 19410
rect 2129 19352 2134 19408
rect 2190 19352 7102 19408
rect 7158 19352 7163 19408
rect 2129 19350 7163 19352
rect 2129 19347 2195 19350
rect 7097 19347 7163 19350
rect 1577 19274 1643 19277
rect 3509 19274 3575 19277
rect 1577 19272 3575 19274
rect 1577 19216 1582 19272
rect 1638 19216 3514 19272
rect 3570 19216 3575 19272
rect 1577 19214 3575 19216
rect 1577 19211 1643 19214
rect 3509 19211 3575 19214
rect 0 19138 480 19168
rect 3049 19138 3115 19141
rect 0 19136 3115 19138
rect 0 19080 3054 19136
rect 3110 19080 3115 19136
rect 0 19078 3115 19080
rect 0 19048 480 19078
rect 3049 19075 3115 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 2589 19002 2655 19005
rect 2865 19002 2931 19005
rect 2589 19000 2931 19002
rect 2589 18944 2594 19000
rect 2650 18944 2870 19000
rect 2926 18944 2931 19000
rect 2589 18942 2931 18944
rect 2589 18939 2655 18942
rect 2865 18939 2931 18942
rect 10961 19002 11027 19005
rect 13721 19002 13787 19005
rect 10961 19000 13787 19002
rect 10961 18944 10966 19000
rect 11022 18944 13726 19000
rect 13782 18944 13787 19000
rect 10961 18942 13787 18944
rect 10961 18939 11027 18942
rect 13721 18939 13787 18942
rect 5625 18866 5691 18869
rect 11237 18866 11303 18869
rect 5625 18864 11303 18866
rect 5625 18808 5630 18864
rect 5686 18808 11242 18864
rect 11298 18808 11303 18864
rect 5625 18806 11303 18808
rect 5625 18803 5691 18806
rect 11237 18803 11303 18806
rect 8017 18730 8083 18733
rect 10133 18730 10199 18733
rect 8017 18728 10199 18730
rect 8017 18672 8022 18728
rect 8078 18672 10138 18728
rect 10194 18672 10199 18728
rect 8017 18670 10199 18672
rect 8017 18667 8083 18670
rect 10133 18667 10199 18670
rect 0 18594 480 18624
rect 2221 18594 2287 18597
rect 0 18592 2287 18594
rect 0 18536 2226 18592
rect 2282 18536 2287 18592
rect 0 18534 2287 18536
rect 0 18504 480 18534
rect 2221 18531 2287 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 1393 18458 1459 18461
rect 5073 18458 5139 18461
rect 1393 18456 5139 18458
rect 1393 18400 1398 18456
rect 1454 18400 5078 18456
rect 5134 18400 5139 18456
rect 1393 18398 5139 18400
rect 1393 18395 1459 18398
rect 5073 18395 5139 18398
rect 1577 18322 1643 18325
rect 2957 18322 3023 18325
rect 1577 18320 3023 18322
rect 1577 18264 1582 18320
rect 1638 18264 2962 18320
rect 3018 18264 3023 18320
rect 1577 18262 3023 18264
rect 1577 18259 1643 18262
rect 2957 18259 3023 18262
rect 3693 18322 3759 18325
rect 6085 18322 6151 18325
rect 3693 18320 6151 18322
rect 3693 18264 3698 18320
rect 3754 18264 6090 18320
rect 6146 18264 6151 18320
rect 3693 18262 6151 18264
rect 3693 18259 3759 18262
rect 6085 18259 6151 18262
rect 6269 18322 6335 18325
rect 10685 18322 10751 18325
rect 6269 18320 10751 18322
rect 6269 18264 6274 18320
rect 6330 18264 10690 18320
rect 10746 18264 10751 18320
rect 6269 18262 10751 18264
rect 6269 18259 6335 18262
rect 10685 18259 10751 18262
rect 1669 18186 1735 18189
rect 4061 18186 4127 18189
rect 1669 18184 4127 18186
rect 1669 18128 1674 18184
rect 1730 18128 4066 18184
rect 4122 18128 4127 18184
rect 1669 18126 4127 18128
rect 1669 18123 1735 18126
rect 4061 18123 4127 18126
rect 8385 18186 8451 18189
rect 14089 18186 14155 18189
rect 8385 18184 14155 18186
rect 8385 18128 8390 18184
rect 8446 18128 14094 18184
rect 14150 18128 14155 18184
rect 8385 18126 14155 18128
rect 8385 18123 8451 18126
rect 14089 18123 14155 18126
rect 0 18050 480 18080
rect 4245 18050 4311 18053
rect 0 18048 4311 18050
rect 0 17992 4250 18048
rect 4306 17992 4311 18048
rect 0 17990 4311 17992
rect 0 17960 480 17990
rect 4245 17987 4311 17990
rect 7649 18050 7715 18053
rect 9489 18050 9555 18053
rect 7649 18048 9555 18050
rect 7649 17992 7654 18048
rect 7710 17992 9494 18048
rect 9550 17992 9555 18048
rect 7649 17990 9555 17992
rect 7649 17987 7715 17990
rect 9489 17987 9555 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 2497 17778 2563 17781
rect 10041 17778 10107 17781
rect 2497 17776 10107 17778
rect 2497 17720 2502 17776
rect 2558 17720 10046 17776
rect 10102 17720 10107 17776
rect 2497 17718 10107 17720
rect 2497 17715 2563 17718
rect 10041 17715 10107 17718
rect 0 17506 480 17536
rect 3877 17506 3943 17509
rect 0 17504 3943 17506
rect 0 17448 3882 17504
rect 3938 17448 3943 17504
rect 0 17446 3943 17448
rect 0 17416 480 17446
rect 3877 17443 3943 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 5993 17370 6059 17373
rect 13169 17370 13235 17373
rect 5993 17368 13235 17370
rect 5993 17312 5998 17368
rect 6054 17312 13174 17368
rect 13230 17312 13235 17368
rect 5993 17310 13235 17312
rect 5993 17307 6059 17310
rect 13169 17307 13235 17310
rect 2497 17236 2563 17237
rect 2446 17172 2452 17236
rect 2516 17234 2563 17236
rect 2516 17232 2608 17234
rect 2558 17176 2608 17232
rect 2516 17174 2608 17176
rect 2516 17172 2563 17174
rect 2497 17171 2563 17172
rect 10777 16962 10843 16965
rect 12433 16962 12499 16965
rect 10777 16960 12499 16962
rect 10777 16904 10782 16960
rect 10838 16904 12438 16960
rect 12494 16904 12499 16960
rect 10777 16902 12499 16904
rect 10777 16899 10843 16902
rect 12433 16899 12499 16902
rect 10277 16896 10597 16897
rect 0 16826 480 16856
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 3693 16826 3759 16829
rect 0 16824 3759 16826
rect 0 16768 3698 16824
rect 3754 16768 3759 16824
rect 0 16766 3759 16768
rect 0 16736 480 16766
rect 3693 16763 3759 16766
rect 3969 16690 4035 16693
rect 5165 16690 5231 16693
rect 5809 16690 5875 16693
rect 3969 16688 5875 16690
rect 3969 16632 3974 16688
rect 4030 16632 5170 16688
rect 5226 16632 5814 16688
rect 5870 16632 5875 16688
rect 3969 16630 5875 16632
rect 3969 16627 4035 16630
rect 5165 16627 5231 16630
rect 5809 16627 5875 16630
rect 8201 16690 8267 16693
rect 11237 16690 11303 16693
rect 8201 16688 11303 16690
rect 8201 16632 8206 16688
rect 8262 16632 11242 16688
rect 11298 16632 11303 16688
rect 8201 16630 11303 16632
rect 8201 16627 8267 16630
rect 11237 16627 11303 16630
rect 5610 16352 5930 16353
rect 0 16282 480 16312
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 3233 16282 3299 16285
rect 0 16280 3299 16282
rect 0 16224 3238 16280
rect 3294 16224 3299 16280
rect 0 16222 3299 16224
rect 0 16192 480 16222
rect 3233 16219 3299 16222
rect 1485 16010 1551 16013
rect 4245 16010 4311 16013
rect 1485 16008 4311 16010
rect 1485 15952 1490 16008
rect 1546 15952 4250 16008
rect 4306 15952 4311 16008
rect 1485 15950 4311 15952
rect 1485 15947 1551 15950
rect 4245 15947 4311 15950
rect 10277 15808 10597 15809
rect 0 15738 480 15768
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 3969 15738 4035 15741
rect 7281 15738 7347 15741
rect 0 15678 2698 15738
rect 0 15648 480 15678
rect 2638 15602 2698 15678
rect 3969 15736 7347 15738
rect 3969 15680 3974 15736
rect 4030 15680 7286 15736
rect 7342 15680 7347 15736
rect 3969 15678 7347 15680
rect 3969 15675 4035 15678
rect 7281 15675 7347 15678
rect 23473 15602 23539 15605
rect 2638 15568 2744 15602
rect 2822 15600 23539 15602
rect 2822 15568 23478 15600
rect 2638 15544 23478 15568
rect 23534 15544 23539 15600
rect 2638 15542 23539 15544
rect 2684 15508 2882 15542
rect 23473 15539 23539 15542
rect 8385 15330 8451 15333
rect 13813 15330 13879 15333
rect 8385 15328 13879 15330
rect 8385 15272 8390 15328
rect 8446 15272 13818 15328
rect 13874 15272 13879 15328
rect 8385 15270 13879 15272
rect 8385 15267 8451 15270
rect 13813 15267 13879 15270
rect 5610 15264 5930 15265
rect 0 15194 480 15224
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 3785 15194 3851 15197
rect 0 15192 3851 15194
rect 0 15136 3790 15192
rect 3846 15136 3851 15192
rect 0 15134 3851 15136
rect 0 15104 480 15134
rect 3785 15131 3851 15134
rect 2681 15058 2747 15061
rect 4613 15058 4679 15061
rect 2681 15056 4679 15058
rect 2681 15000 2686 15056
rect 2742 15000 4618 15056
rect 4674 15000 4679 15056
rect 2681 14998 4679 15000
rect 2681 14995 2747 14998
rect 4613 14995 4679 14998
rect 5625 15058 5691 15061
rect 9765 15058 9831 15061
rect 5625 15056 9831 15058
rect 5625 15000 5630 15056
rect 5686 15000 9770 15056
rect 9826 15000 9831 15056
rect 5625 14998 9831 15000
rect 5625 14995 5691 14998
rect 9765 14995 9831 14998
rect 8661 14922 8727 14925
rect 11881 14922 11947 14925
rect 8661 14920 11947 14922
rect 8661 14864 8666 14920
rect 8722 14864 11886 14920
rect 11942 14864 11947 14920
rect 8661 14862 11947 14864
rect 8661 14859 8727 14862
rect 11881 14859 11947 14862
rect 5625 14786 5691 14789
rect 7557 14786 7623 14789
rect 5625 14784 7623 14786
rect 5625 14728 5630 14784
rect 5686 14728 7562 14784
rect 7618 14728 7623 14784
rect 5625 14726 7623 14728
rect 5625 14723 5691 14726
rect 7557 14723 7623 14726
rect 10277 14720 10597 14721
rect 0 14650 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 3417 14650 3483 14653
rect 0 14648 3483 14650
rect 0 14592 3422 14648
rect 3478 14592 3483 14648
rect 0 14590 3483 14592
rect 0 14560 480 14590
rect 3417 14587 3483 14590
rect 5165 14650 5231 14653
rect 6729 14650 6795 14653
rect 8753 14650 8819 14653
rect 5165 14648 8819 14650
rect 5165 14592 5170 14648
rect 5226 14592 6734 14648
rect 6790 14592 8758 14648
rect 8814 14592 8819 14648
rect 5165 14590 8819 14592
rect 5165 14587 5231 14590
rect 6729 14587 6795 14590
rect 8753 14587 8819 14590
rect 9121 14514 9187 14517
rect 12985 14514 13051 14517
rect 9121 14512 13051 14514
rect 9121 14456 9126 14512
rect 9182 14456 12990 14512
rect 13046 14456 13051 14512
rect 9121 14454 13051 14456
rect 9121 14451 9187 14454
rect 12985 14451 13051 14454
rect 4705 14378 4771 14381
rect 12801 14378 12867 14381
rect 4705 14376 12867 14378
rect 4705 14320 4710 14376
rect 4766 14320 12806 14376
rect 12862 14320 12867 14376
rect 4705 14318 12867 14320
rect 4705 14315 4771 14318
rect 12801 14315 12867 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 7649 14106 7715 14109
rect 8293 14106 8359 14109
rect 9949 14106 10015 14109
rect 7649 14104 10015 14106
rect 7649 14048 7654 14104
rect 7710 14048 8298 14104
rect 8354 14048 9954 14104
rect 10010 14048 10015 14104
rect 7649 14046 10015 14048
rect 7649 14043 7715 14046
rect 8293 14043 8359 14046
rect 9949 14043 10015 14046
rect 0 13970 480 14000
rect 3785 13970 3851 13973
rect 23657 13970 23723 13973
rect 0 13910 2744 13970
rect 0 13880 480 13910
rect 2684 13834 2744 13910
rect 3785 13968 23723 13970
rect 3785 13912 3790 13968
rect 3846 13912 23662 13968
rect 23718 13912 23723 13968
rect 3785 13910 23723 13912
rect 3785 13907 3851 13910
rect 23657 13907 23723 13910
rect 23841 13970 23907 13973
rect 27520 13970 28000 14000
rect 23841 13968 28000 13970
rect 23841 13912 23846 13968
rect 23902 13912 28000 13968
rect 23841 13910 28000 13912
rect 23841 13907 23907 13910
rect 27520 13880 28000 13910
rect 6177 13834 6243 13837
rect 2684 13832 6243 13834
rect 2684 13776 6182 13832
rect 6238 13776 6243 13832
rect 2684 13774 6243 13776
rect 6177 13771 6243 13774
rect 7833 13834 7899 13837
rect 10133 13834 10199 13837
rect 7833 13832 10199 13834
rect 7833 13776 7838 13832
rect 7894 13776 10138 13832
rect 10194 13776 10199 13832
rect 7833 13774 10199 13776
rect 7833 13771 7899 13774
rect 10133 13771 10199 13774
rect 10777 13698 10843 13701
rect 12433 13698 12499 13701
rect 10777 13696 12499 13698
rect 10777 13640 10782 13696
rect 10838 13640 12438 13696
rect 12494 13640 12499 13696
rect 10777 13638 12499 13640
rect 10777 13635 10843 13638
rect 12433 13635 12499 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 3417 13562 3483 13565
rect 10041 13562 10107 13565
rect 3417 13560 10107 13562
rect 3417 13504 3422 13560
rect 3478 13504 10046 13560
rect 10102 13504 10107 13560
rect 3417 13502 10107 13504
rect 3417 13499 3483 13502
rect 10041 13499 10107 13502
rect 0 13426 480 13456
rect 6453 13426 6519 13429
rect 0 13424 6519 13426
rect 0 13368 6458 13424
rect 6514 13368 6519 13424
rect 0 13366 6519 13368
rect 0 13336 480 13366
rect 6453 13363 6519 13366
rect 9213 13426 9279 13429
rect 12157 13426 12223 13429
rect 9213 13424 12223 13426
rect 9213 13368 9218 13424
rect 9274 13368 12162 13424
rect 12218 13368 12223 13424
rect 9213 13366 12223 13368
rect 9213 13363 9279 13366
rect 12157 13363 12223 13366
rect 3877 13290 3943 13293
rect 6269 13290 6335 13293
rect 11237 13290 11303 13293
rect 3877 13288 6194 13290
rect 3877 13232 3882 13288
rect 3938 13232 6194 13288
rect 3877 13230 6194 13232
rect 3877 13227 3943 13230
rect 6134 13154 6194 13230
rect 6269 13288 11303 13290
rect 6269 13232 6274 13288
rect 6330 13232 11242 13288
rect 11298 13232 11303 13288
rect 6269 13230 11303 13232
rect 6269 13227 6335 13230
rect 11237 13227 11303 13230
rect 12433 13154 12499 13157
rect 6134 13152 12499 13154
rect 6134 13096 12438 13152
rect 12494 13096 12499 13152
rect 6134 13094 12499 13096
rect 12433 13091 12499 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 6821 13018 6887 13021
rect 12893 13018 12959 13021
rect 6821 13016 12959 13018
rect 6821 12960 6826 13016
rect 6882 12960 12898 13016
rect 12954 12960 12959 13016
rect 6821 12958 12959 12960
rect 6821 12955 6887 12958
rect 12893 12955 12959 12958
rect 0 12882 480 12912
rect 8569 12882 8635 12885
rect 12433 12882 12499 12885
rect 0 12822 2744 12882
rect 0 12792 480 12822
rect 2684 12780 2744 12822
rect 8569 12880 12499 12882
rect 8569 12824 8574 12880
rect 8630 12824 12438 12880
rect 12494 12824 12499 12880
rect 8569 12822 12499 12824
rect 8569 12819 8635 12822
rect 12433 12819 12499 12822
rect 2684 12746 2882 12780
rect 10133 12746 10199 12749
rect 2684 12744 10199 12746
rect 2684 12720 10138 12744
rect 2822 12688 10138 12720
rect 10194 12688 10199 12744
rect 2822 12686 10199 12688
rect 10133 12683 10199 12686
rect 10317 12746 10383 12749
rect 22277 12746 22343 12749
rect 10317 12744 22343 12746
rect 10317 12688 10322 12744
rect 10378 12688 22282 12744
rect 22338 12688 22343 12744
rect 10317 12686 22343 12688
rect 10317 12683 10383 12686
rect 22277 12683 22343 12686
rect 6361 12610 6427 12613
rect 7373 12610 7439 12613
rect 6361 12608 7439 12610
rect 6361 12552 6366 12608
rect 6422 12552 7378 12608
rect 7434 12552 7439 12608
rect 6361 12550 7439 12552
rect 6361 12547 6427 12550
rect 7373 12547 7439 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 1669 12474 1735 12477
rect 5073 12474 5139 12477
rect 1669 12472 5139 12474
rect 1669 12416 1674 12472
rect 1730 12416 5078 12472
rect 5134 12416 5139 12472
rect 1669 12414 5139 12416
rect 1669 12411 1735 12414
rect 5073 12411 5139 12414
rect 0 12338 480 12368
rect 1301 12338 1367 12341
rect 0 12336 1367 12338
rect 0 12280 1306 12336
rect 1362 12280 1367 12336
rect 0 12278 1367 12280
rect 0 12248 480 12278
rect 1301 12275 1367 12278
rect 3141 12338 3207 12341
rect 4153 12338 4219 12341
rect 3141 12336 4219 12338
rect 3141 12280 3146 12336
rect 3202 12280 4158 12336
rect 4214 12280 4219 12336
rect 3141 12278 4219 12280
rect 3141 12275 3207 12278
rect 4153 12275 4219 12278
rect 4797 12338 4863 12341
rect 5533 12338 5599 12341
rect 4797 12336 5599 12338
rect 4797 12280 4802 12336
rect 4858 12280 5538 12336
rect 5594 12280 5599 12336
rect 4797 12278 5599 12280
rect 4797 12275 4863 12278
rect 5533 12275 5599 12278
rect 7097 12338 7163 12341
rect 11605 12338 11671 12341
rect 7097 12336 11671 12338
rect 7097 12280 7102 12336
rect 7158 12280 11610 12336
rect 11666 12280 11671 12336
rect 7097 12278 11671 12280
rect 7097 12275 7163 12278
rect 11605 12275 11671 12278
rect 9121 12202 9187 12205
rect 11789 12202 11855 12205
rect 9121 12200 11855 12202
rect 9121 12144 9126 12200
rect 9182 12144 11794 12200
rect 11850 12144 11855 12200
rect 9121 12142 11855 12144
rect 9121 12139 9187 12142
rect 11789 12139 11855 12142
rect 10133 12066 10199 12069
rect 14549 12066 14615 12069
rect 10133 12064 14615 12066
rect 10133 12008 10138 12064
rect 10194 12008 14554 12064
rect 14610 12008 14615 12064
rect 10133 12006 14615 12008
rect 10133 12003 10199 12006
rect 14549 12003 14615 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 7925 11930 7991 11933
rect 10041 11930 10107 11933
rect 5996 11928 10107 11930
rect 5996 11872 7930 11928
rect 7986 11872 10046 11928
rect 10102 11872 10107 11928
rect 5996 11870 10107 11872
rect 0 11794 480 11824
rect 2957 11794 3023 11797
rect 5996 11794 6056 11870
rect 7925 11867 7991 11870
rect 10041 11867 10107 11870
rect 0 11734 2882 11794
rect 0 11704 480 11734
rect 2822 11658 2882 11734
rect 2957 11792 6056 11794
rect 2957 11736 2962 11792
rect 3018 11736 6056 11792
rect 2957 11734 6056 11736
rect 6177 11794 6243 11797
rect 21725 11794 21791 11797
rect 6177 11792 21791 11794
rect 6177 11736 6182 11792
rect 6238 11736 21730 11792
rect 21786 11736 21791 11792
rect 6177 11734 21791 11736
rect 2957 11731 3023 11734
rect 6177 11731 6243 11734
rect 21725 11731 21791 11734
rect 7005 11658 7071 11661
rect 2822 11656 7071 11658
rect 2822 11600 7010 11656
rect 7066 11600 7071 11656
rect 2822 11598 7071 11600
rect 7005 11595 7071 11598
rect 12709 11658 12775 11661
rect 23841 11658 23907 11661
rect 12709 11656 23907 11658
rect 12709 11600 12714 11656
rect 12770 11600 23846 11656
rect 23902 11600 23907 11656
rect 12709 11598 23907 11600
rect 12709 11595 12775 11598
rect 23841 11595 23907 11598
rect 2589 11522 2655 11525
rect 6361 11522 6427 11525
rect 2589 11520 6427 11522
rect 2589 11464 2594 11520
rect 2650 11464 6366 11520
rect 6422 11464 6427 11520
rect 2589 11462 6427 11464
rect 2589 11459 2655 11462
rect 6361 11459 6427 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 3877 11386 3943 11389
rect 6085 11386 6151 11389
rect 3877 11384 6151 11386
rect 3877 11328 3882 11384
rect 3938 11328 6090 11384
rect 6146 11328 6151 11384
rect 3877 11326 6151 11328
rect 3877 11323 3943 11326
rect 6085 11323 6151 11326
rect 8201 11250 8267 11253
rect 11053 11250 11119 11253
rect 8201 11248 11119 11250
rect 8201 11192 8206 11248
rect 8262 11192 11058 11248
rect 11114 11192 11119 11248
rect 8201 11190 11119 11192
rect 8201 11187 8267 11190
rect 11053 11187 11119 11190
rect 0 11114 480 11144
rect 3601 11114 3667 11117
rect 0 11112 3667 11114
rect 0 11056 3606 11112
rect 3662 11056 3667 11112
rect 0 11054 3667 11056
rect 0 11024 480 11054
rect 3601 11051 3667 11054
rect 8017 11114 8083 11117
rect 8661 11114 8727 11117
rect 10133 11114 10199 11117
rect 8017 11112 10199 11114
rect 8017 11056 8022 11112
rect 8078 11056 8666 11112
rect 8722 11056 10138 11112
rect 10194 11056 10199 11112
rect 8017 11054 10199 11056
rect 8017 11051 8083 11054
rect 8661 11051 8727 11054
rect 10133 11051 10199 11054
rect 21909 11114 21975 11117
rect 23565 11114 23631 11117
rect 21909 11112 23631 11114
rect 21909 11056 21914 11112
rect 21970 11056 23570 11112
rect 23626 11056 23631 11112
rect 21909 11054 23631 11056
rect 21909 11051 21975 11054
rect 23565 11051 23631 11054
rect 7649 10978 7715 10981
rect 9673 10978 9739 10981
rect 7649 10976 9739 10978
rect 7649 10920 7654 10976
rect 7710 10920 9678 10976
rect 9734 10920 9739 10976
rect 7649 10918 9739 10920
rect 7649 10915 7715 10918
rect 9673 10915 9739 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 8845 10842 8911 10845
rect 10777 10842 10843 10845
rect 8845 10840 10843 10842
rect 8845 10784 8850 10840
rect 8906 10784 10782 10840
rect 10838 10784 10843 10840
rect 8845 10782 10843 10784
rect 8845 10779 8911 10782
rect 10777 10779 10843 10782
rect 0 10570 480 10600
rect 4429 10570 4495 10573
rect 12801 10570 12867 10573
rect 0 10510 1410 10570
rect 0 10480 480 10510
rect 1350 10434 1410 10510
rect 4429 10568 12867 10570
rect 4429 10512 4434 10568
rect 4490 10512 12806 10568
rect 12862 10512 12867 10568
rect 4429 10510 12867 10512
rect 4429 10507 4495 10510
rect 12801 10507 12867 10510
rect 7649 10434 7715 10437
rect 1350 10432 7715 10434
rect 1350 10376 7654 10432
rect 7710 10376 7715 10432
rect 1350 10374 7715 10376
rect 7649 10371 7715 10374
rect 11145 10434 11211 10437
rect 14273 10434 14339 10437
rect 11145 10432 14339 10434
rect 11145 10376 11150 10432
rect 11206 10376 14278 10432
rect 14334 10376 14339 10432
rect 11145 10374 14339 10376
rect 11145 10371 11211 10374
rect 14273 10371 14339 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 4981 10298 5047 10301
rect 8385 10298 8451 10301
rect 4981 10296 8451 10298
rect 4981 10240 4986 10296
rect 5042 10240 8390 10296
rect 8446 10240 8451 10296
rect 4981 10238 8451 10240
rect 4981 10235 5047 10238
rect 8385 10235 8451 10238
rect 2405 10162 2471 10165
rect 6821 10162 6887 10165
rect 11605 10162 11671 10165
rect 2405 10160 3618 10162
rect 2405 10104 2410 10160
rect 2466 10104 3618 10160
rect 2405 10102 3618 10104
rect 2405 10099 2471 10102
rect 0 10026 480 10056
rect 3558 10026 3618 10102
rect 6821 10160 11671 10162
rect 6821 10104 6826 10160
rect 6882 10104 11610 10160
rect 11666 10104 11671 10160
rect 6821 10102 11671 10104
rect 6821 10099 6887 10102
rect 11605 10099 11671 10102
rect 3693 10026 3759 10029
rect 6729 10026 6795 10029
rect 0 9966 3480 10026
rect 3558 10024 6795 10026
rect 3558 9968 3698 10024
rect 3754 9968 6734 10024
rect 6790 9968 6795 10024
rect 3558 9966 6795 9968
rect 0 9936 480 9966
rect 3420 9890 3480 9966
rect 3693 9963 3759 9966
rect 6729 9963 6795 9966
rect 6913 10026 6979 10029
rect 13169 10026 13235 10029
rect 6913 10024 13235 10026
rect 6913 9968 6918 10024
rect 6974 9968 13174 10024
rect 13230 9968 13235 10024
rect 6913 9966 13235 9968
rect 6913 9963 6979 9966
rect 13169 9963 13235 9966
rect 5349 9890 5415 9893
rect 3420 9888 5415 9890
rect 3420 9832 5354 9888
rect 5410 9832 5415 9888
rect 3420 9830 5415 9832
rect 5349 9827 5415 9830
rect 7005 9890 7071 9893
rect 12525 9890 12591 9893
rect 7005 9888 12591 9890
rect 7005 9832 7010 9888
rect 7066 9832 12530 9888
rect 12586 9832 12591 9888
rect 7005 9830 12591 9832
rect 7005 9827 7071 9830
rect 12525 9827 12591 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 1485 9754 1551 9757
rect 2497 9754 2563 9757
rect 1485 9752 2563 9754
rect 1485 9696 1490 9752
rect 1546 9696 2502 9752
rect 2558 9696 2563 9752
rect 1485 9694 2563 9696
rect 1485 9691 1551 9694
rect 2497 9691 2563 9694
rect 5993 9754 6059 9757
rect 13445 9754 13511 9757
rect 5993 9752 13511 9754
rect 5993 9696 5998 9752
rect 6054 9696 13450 9752
rect 13506 9696 13511 9752
rect 5993 9694 13511 9696
rect 5993 9691 6059 9694
rect 13445 9691 13511 9694
rect 7373 9618 7439 9621
rect 7373 9616 9506 9618
rect 7373 9560 7378 9616
rect 7434 9584 9506 9616
rect 9622 9584 9628 9620
rect 7434 9560 9628 9584
rect 7373 9558 9628 9560
rect 7373 9555 7439 9558
rect 9446 9556 9628 9558
rect 9692 9556 9698 9620
rect 12934 9556 12940 9620
rect 13004 9618 13010 9620
rect 13629 9618 13695 9621
rect 13004 9616 13695 9618
rect 13004 9560 13634 9616
rect 13690 9560 13695 9616
rect 13004 9558 13695 9560
rect 13004 9556 13010 9558
rect 9446 9524 9690 9556
rect 13629 9555 13695 9558
rect 0 9482 480 9512
rect 3877 9482 3943 9485
rect 0 9480 3943 9482
rect 0 9424 3882 9480
rect 3938 9424 3943 9480
rect 0 9422 3943 9424
rect 0 9392 480 9422
rect 3877 9419 3943 9422
rect 7097 9482 7163 9485
rect 12157 9482 12223 9485
rect 7097 9480 9184 9482
rect 7097 9424 7102 9480
rect 7158 9448 9184 9480
rect 9768 9480 12223 9482
rect 9768 9448 12162 9480
rect 7158 9424 12162 9448
rect 12218 9424 12223 9480
rect 7097 9422 12223 9424
rect 7097 9419 7163 9422
rect 9124 9388 9828 9422
rect 12157 9419 12223 9422
rect 6361 9346 6427 9349
rect 8293 9346 8359 9349
rect 8845 9346 8911 9349
rect 6361 9344 8911 9346
rect 6361 9288 6366 9344
rect 6422 9288 8298 9344
rect 8354 9288 8850 9344
rect 8906 9288 8911 9344
rect 6361 9286 8911 9288
rect 6361 9283 6427 9286
rect 8293 9283 8359 9286
rect 8845 9283 8911 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 6453 9210 6519 9213
rect 10133 9210 10199 9213
rect 6453 9208 10199 9210
rect 6453 9152 6458 9208
rect 6514 9152 10138 9208
rect 10194 9152 10199 9208
rect 6453 9150 10199 9152
rect 6453 9147 6519 9150
rect 10133 9147 10199 9150
rect 4061 9074 4127 9077
rect 6177 9074 6243 9077
rect 4061 9072 6243 9074
rect 4061 9016 4066 9072
rect 4122 9016 6182 9072
rect 6238 9016 6243 9072
rect 4061 9014 6243 9016
rect 4061 9011 4127 9014
rect 6177 9011 6243 9014
rect 9622 9012 9628 9076
rect 9692 9074 9698 9076
rect 12433 9074 12499 9077
rect 9692 9072 12499 9074
rect 9692 9016 12438 9072
rect 12494 9016 12499 9072
rect 9692 9014 12499 9016
rect 9692 9012 9698 9014
rect 12433 9011 12499 9014
rect 0 8938 480 8968
rect 8293 8938 8359 8941
rect 0 8936 8359 8938
rect 0 8880 8298 8936
rect 8354 8880 8359 8936
rect 0 8878 8359 8880
rect 0 8848 480 8878
rect 8293 8875 8359 8878
rect 1945 8802 2011 8805
rect 2446 8802 2452 8804
rect 1945 8800 2452 8802
rect 1945 8744 1950 8800
rect 2006 8744 2452 8800
rect 1945 8742 2452 8744
rect 1945 8739 2011 8742
rect 2446 8740 2452 8742
rect 2516 8740 2522 8804
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 8845 8666 8911 8669
rect 11237 8666 11303 8669
rect 8845 8664 11303 8666
rect 8845 8608 8850 8664
rect 8906 8608 11242 8664
rect 11298 8608 11303 8664
rect 8845 8606 11303 8608
rect 8845 8603 8911 8606
rect 11237 8603 11303 8606
rect 3693 8530 3759 8533
rect 4061 8530 4127 8533
rect 3693 8528 4127 8530
rect 3693 8472 3698 8528
rect 3754 8472 4066 8528
rect 4122 8472 4127 8528
rect 3693 8470 4127 8472
rect 3693 8467 3759 8470
rect 4061 8467 4127 8470
rect 4337 8530 4403 8533
rect 8293 8530 8359 8533
rect 4337 8528 8359 8530
rect 4337 8472 4342 8528
rect 4398 8472 8298 8528
rect 8354 8472 8359 8528
rect 4337 8470 8359 8472
rect 4337 8467 4403 8470
rect 8293 8467 8359 8470
rect 10961 8530 11027 8533
rect 17125 8530 17191 8533
rect 10961 8528 17191 8530
rect 10961 8472 10966 8528
rect 11022 8472 17130 8528
rect 17186 8472 17191 8528
rect 10961 8470 17191 8472
rect 10961 8467 11027 8470
rect 17125 8467 17191 8470
rect 5165 8394 5231 8397
rect 7097 8394 7163 8397
rect 5165 8392 7163 8394
rect 5165 8336 5170 8392
rect 5226 8336 7102 8392
rect 7158 8336 7163 8392
rect 5165 8334 7163 8336
rect 5165 8331 5231 8334
rect 7097 8331 7163 8334
rect 9489 8394 9555 8397
rect 11513 8394 11579 8397
rect 14457 8394 14523 8397
rect 9489 8392 14523 8394
rect 9489 8336 9494 8392
rect 9550 8336 11518 8392
rect 11574 8336 14462 8392
rect 14518 8336 14523 8392
rect 9489 8334 14523 8336
rect 9489 8331 9555 8334
rect 11513 8331 11579 8334
rect 14457 8331 14523 8334
rect 0 8258 480 8288
rect 20161 8258 20227 8261
rect 24761 8258 24827 8261
rect 0 8198 4906 8258
rect 0 8168 480 8198
rect 4846 7986 4906 8198
rect 20161 8256 24827 8258
rect 20161 8200 20166 8256
rect 20222 8200 24766 8256
rect 24822 8200 24827 8256
rect 20161 8198 24827 8200
rect 20161 8195 20227 8198
rect 24761 8195 24827 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 5073 8122 5139 8125
rect 6545 8122 6611 8125
rect 5073 8120 6611 8122
rect 5073 8064 5078 8120
rect 5134 8064 6550 8120
rect 6606 8064 6611 8120
rect 5073 8062 6611 8064
rect 5073 8059 5139 8062
rect 6545 8059 6611 8062
rect 12985 7986 13051 7989
rect 4846 7984 13051 7986
rect 4846 7928 12990 7984
rect 13046 7928 13051 7984
rect 4846 7926 13051 7928
rect 12985 7923 13051 7926
rect 5625 7850 5691 7853
rect 7465 7850 7531 7853
rect 12525 7850 12591 7853
rect 5625 7848 6056 7850
rect 5625 7792 5630 7848
rect 5686 7792 6056 7848
rect 5625 7790 6056 7792
rect 5625 7787 5691 7790
rect 0 7714 480 7744
rect 5996 7714 6056 7790
rect 7465 7848 12591 7850
rect 7465 7792 7470 7848
rect 7526 7792 12530 7848
rect 12586 7792 12591 7848
rect 7465 7790 12591 7792
rect 7465 7787 7531 7790
rect 12525 7787 12591 7790
rect 12709 7714 12775 7717
rect 0 7654 4906 7714
rect 5996 7712 12775 7714
rect 5996 7656 12714 7712
rect 12770 7656 12775 7712
rect 5996 7654 12775 7656
rect 0 7624 480 7654
rect 4846 7442 4906 7654
rect 12709 7651 12775 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 9489 7576 9555 7581
rect 9489 7520 9494 7576
rect 9550 7544 9555 7576
rect 9622 7544 9628 7580
rect 9550 7520 9628 7544
rect 9489 7516 9628 7520
rect 9692 7516 9698 7580
rect 9489 7515 9690 7516
rect 9492 7484 9690 7515
rect 11789 7442 11855 7445
rect 4846 7408 9368 7442
rect 9768 7440 11855 7442
rect 9768 7408 11794 7440
rect 4846 7384 11794 7408
rect 11850 7384 11855 7440
rect 4846 7382 11855 7384
rect 9308 7348 9828 7382
rect 11789 7379 11855 7382
rect 2221 7306 2287 7309
rect 3509 7306 3575 7309
rect 2221 7304 3575 7306
rect 2221 7248 2226 7304
rect 2282 7248 3514 7304
rect 3570 7248 3575 7304
rect 2221 7246 3575 7248
rect 2221 7243 2287 7246
rect 3509 7243 3575 7246
rect 0 7170 480 7200
rect 4061 7170 4127 7173
rect 0 7168 4127 7170
rect 0 7112 4066 7168
rect 4122 7112 4127 7168
rect 0 7110 4127 7112
rect 0 7080 480 7110
rect 4061 7107 4127 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 5165 7034 5231 7037
rect 8201 7034 8267 7037
rect 5165 7032 8267 7034
rect 5165 6976 5170 7032
rect 5226 6976 8206 7032
rect 8262 6976 8267 7032
rect 5165 6974 8267 6976
rect 5165 6971 5231 6974
rect 8201 6971 8267 6974
rect 3601 6898 3667 6901
rect 6361 6898 6427 6901
rect 3601 6896 6427 6898
rect 3601 6840 3606 6896
rect 3662 6840 6366 6896
rect 6422 6840 6427 6896
rect 3601 6838 6427 6840
rect 3601 6835 3667 6838
rect 6361 6835 6427 6838
rect 10777 6898 10843 6901
rect 17861 6898 17927 6901
rect 10777 6896 17927 6898
rect 10777 6840 10782 6896
rect 10838 6840 17866 6896
rect 17922 6840 17927 6896
rect 10777 6838 17927 6840
rect 10777 6835 10843 6838
rect 17861 6835 17927 6838
rect 2497 6762 2563 6765
rect 4521 6762 4587 6765
rect 2497 6760 4587 6762
rect 2497 6704 2502 6760
rect 2558 6704 4526 6760
rect 4582 6704 4587 6760
rect 2497 6702 4587 6704
rect 2497 6699 2563 6702
rect 4521 6699 4587 6702
rect 7741 6762 7807 6765
rect 19057 6762 19123 6765
rect 7741 6760 19123 6762
rect 7741 6704 7746 6760
rect 7802 6704 19062 6760
rect 19118 6704 19123 6760
rect 7741 6702 19123 6704
rect 7741 6699 7807 6702
rect 19057 6699 19123 6702
rect 0 6626 480 6656
rect 4613 6626 4679 6629
rect 0 6624 4679 6626
rect 0 6568 4618 6624
rect 4674 6568 4679 6624
rect 0 6566 4679 6568
rect 0 6536 480 6566
rect 4613 6563 4679 6566
rect 9397 6626 9463 6629
rect 12985 6626 13051 6629
rect 9397 6624 13051 6626
rect 9397 6568 9402 6624
rect 9458 6568 12990 6624
rect 13046 6568 13051 6624
rect 9397 6566 13051 6568
rect 9397 6563 9463 6566
rect 12985 6563 13051 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 6821 6490 6887 6493
rect 14181 6490 14247 6493
rect 6821 6488 14247 6490
rect 6821 6432 6826 6488
rect 6882 6432 14186 6488
rect 14242 6432 14247 6488
rect 6821 6430 14247 6432
rect 6821 6427 6887 6430
rect 14181 6427 14247 6430
rect 7373 6354 7439 6357
rect 10317 6354 10383 6357
rect 7373 6352 10383 6354
rect 7373 6296 7378 6352
rect 7434 6296 10322 6352
rect 10378 6296 10383 6352
rect 7373 6294 10383 6296
rect 7373 6291 7439 6294
rect 10317 6291 10383 6294
rect 15929 6354 15995 6357
rect 19517 6354 19583 6357
rect 15929 6352 19583 6354
rect 15929 6296 15934 6352
rect 15990 6296 19522 6352
rect 19578 6296 19583 6352
rect 15929 6294 19583 6296
rect 15929 6291 15995 6294
rect 19517 6291 19583 6294
rect 9305 6218 9371 6221
rect 12801 6218 12867 6221
rect 9305 6216 12867 6218
rect 9305 6160 9310 6216
rect 9366 6160 12806 6216
rect 12862 6160 12867 6216
rect 9305 6158 12867 6160
rect 9305 6155 9371 6158
rect 12801 6155 12867 6158
rect 14825 6218 14891 6221
rect 16573 6218 16639 6221
rect 14825 6216 16639 6218
rect 14825 6160 14830 6216
rect 14886 6160 16578 6216
rect 16634 6160 16639 6216
rect 14825 6158 16639 6160
rect 14825 6155 14891 6158
rect 16573 6155 16639 6158
rect 16849 6218 16915 6221
rect 22461 6218 22527 6221
rect 16849 6216 22527 6218
rect 16849 6160 16854 6216
rect 16910 6160 22466 6216
rect 22522 6160 22527 6216
rect 16849 6158 22527 6160
rect 16849 6155 16915 6158
rect 22461 6155 22527 6158
rect 0 6082 480 6112
rect 1577 6082 1643 6085
rect 13169 6082 13235 6085
rect 14733 6082 14799 6085
rect 0 6080 1643 6082
rect 0 6024 1582 6080
rect 1638 6024 1643 6080
rect 0 6022 1643 6024
rect 0 5992 480 6022
rect 1577 6019 1643 6022
rect 10734 6080 14799 6082
rect 10734 6024 13174 6080
rect 13230 6024 14738 6080
rect 14794 6024 14799 6080
rect 10734 6022 14799 6024
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 6085 5810 6151 5813
rect 10734 5810 10794 6022
rect 13169 6019 13235 6022
rect 14733 6019 14799 6022
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 6085 5808 10794 5810
rect 6085 5752 6090 5808
rect 6146 5752 10794 5808
rect 6085 5750 10794 5752
rect 12525 5810 12591 5813
rect 20253 5810 20319 5813
rect 12525 5808 20319 5810
rect 12525 5752 12530 5808
rect 12586 5752 20258 5808
rect 20314 5752 20319 5808
rect 12525 5750 20319 5752
rect 6085 5747 6151 5750
rect 12525 5747 12591 5750
rect 20253 5747 20319 5750
rect 2129 5674 2195 5677
rect 5073 5674 5139 5677
rect 2129 5672 5139 5674
rect 2129 5616 2134 5672
rect 2190 5616 5078 5672
rect 5134 5616 5139 5672
rect 2129 5614 5139 5616
rect 2129 5611 2195 5614
rect 5073 5611 5139 5614
rect 7833 5674 7899 5677
rect 15653 5674 15719 5677
rect 7833 5672 15719 5674
rect 7833 5616 7838 5672
rect 7894 5616 15658 5672
rect 15714 5616 15719 5672
rect 7833 5614 15719 5616
rect 7833 5611 7899 5614
rect 15653 5611 15719 5614
rect 15837 5674 15903 5677
rect 18045 5674 18111 5677
rect 15837 5672 18111 5674
rect 15837 5616 15842 5672
rect 15898 5616 18050 5672
rect 18106 5616 18111 5672
rect 15837 5614 18111 5616
rect 15837 5611 15903 5614
rect 18045 5611 18111 5614
rect 3325 5538 3391 5541
rect 3969 5538 4035 5541
rect 3325 5536 4035 5538
rect 3325 5480 3330 5536
rect 3386 5480 3974 5536
rect 4030 5480 4035 5536
rect 3325 5478 4035 5480
rect 3325 5475 3391 5478
rect 3969 5475 4035 5478
rect 5610 5472 5930 5473
rect 0 5402 480 5432
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 4705 5402 4771 5405
rect 0 5400 4771 5402
rect 0 5344 4710 5400
rect 4766 5344 4771 5400
rect 0 5342 4771 5344
rect 0 5312 480 5342
rect 4705 5339 4771 5342
rect 9622 5340 9628 5404
rect 9692 5402 9698 5404
rect 14641 5402 14707 5405
rect 9692 5400 14707 5402
rect 9692 5344 14646 5400
rect 14702 5344 14707 5400
rect 9692 5342 14707 5344
rect 9692 5340 9698 5342
rect 14641 5339 14707 5342
rect 14733 5266 14799 5269
rect 21357 5266 21423 5269
rect 14733 5264 21423 5266
rect 14733 5208 14738 5264
rect 14794 5208 21362 5264
rect 21418 5208 21423 5264
rect 14733 5206 21423 5208
rect 14733 5203 14799 5206
rect 21357 5203 21423 5206
rect 3693 5130 3759 5133
rect 3877 5130 3943 5133
rect 7005 5130 7071 5133
rect 14733 5130 14799 5133
rect 3693 5128 7071 5130
rect 3693 5072 3698 5128
rect 3754 5072 3882 5128
rect 3938 5072 7010 5128
rect 7066 5072 7071 5128
rect 3693 5070 7071 5072
rect 3693 5067 3759 5070
rect 3877 5067 3943 5070
rect 7005 5067 7071 5070
rect 7238 5128 14799 5130
rect 7238 5072 14738 5128
rect 14794 5072 14799 5128
rect 7238 5070 14799 5072
rect 2865 4994 2931 4997
rect 6085 4994 6151 4997
rect 2865 4992 6151 4994
rect 2865 4936 2870 4992
rect 2926 4936 6090 4992
rect 6146 4936 6151 4992
rect 2865 4934 6151 4936
rect 2865 4931 2931 4934
rect 6085 4931 6151 4934
rect 0 4858 480 4888
rect 3601 4858 3667 4861
rect 0 4856 3667 4858
rect 0 4800 3606 4856
rect 3662 4800 3667 4856
rect 0 4798 3667 4800
rect 0 4768 480 4798
rect 3601 4795 3667 4798
rect 3969 4858 4035 4861
rect 7238 4858 7298 5070
rect 14733 5067 14799 5070
rect 10869 4994 10935 4997
rect 10869 4992 17234 4994
rect 10869 4936 10874 4992
rect 10930 4936 17234 4992
rect 10869 4934 17234 4936
rect 10869 4931 10935 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 3969 4856 7298 4858
rect 3969 4800 3974 4856
rect 4030 4800 7298 4856
rect 3969 4798 7298 4800
rect 3969 4795 4035 4798
rect 1853 4722 1919 4725
rect 6545 4722 6611 4725
rect 1853 4720 6611 4722
rect 1853 4664 1858 4720
rect 1914 4664 6550 4720
rect 6606 4664 6611 4720
rect 1853 4662 6611 4664
rect 1853 4659 1919 4662
rect 6545 4659 6611 4662
rect 8017 4722 8083 4725
rect 17174 4722 17234 4934
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 27520 4722 28000 4752
rect 8017 4720 15946 4722
rect 8017 4664 8022 4720
rect 8078 4664 15946 4720
rect 8017 4662 15946 4664
rect 17174 4662 28000 4722
rect 8017 4659 8083 4662
rect 11145 4586 11211 4589
rect 11145 4584 15762 4586
rect 11145 4528 11150 4584
rect 11206 4528 15762 4584
rect 11145 4526 15762 4528
rect 11145 4523 11211 4526
rect 6361 4450 6427 4453
rect 12433 4450 12499 4453
rect 6361 4448 12499 4450
rect 6361 4392 6366 4448
rect 6422 4392 12438 4448
rect 12494 4392 12499 4448
rect 6361 4390 12499 4392
rect 6361 4387 6427 4390
rect 12433 4387 12499 4390
rect 12801 4450 12867 4453
rect 12934 4450 12940 4452
rect 12801 4448 12940 4450
rect 12801 4392 12806 4448
rect 12862 4392 12940 4448
rect 12801 4390 12940 4392
rect 12801 4387 12867 4390
rect 12934 4388 12940 4390
rect 13004 4388 13010 4452
rect 5610 4384 5930 4385
rect 0 4314 480 4344
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 3693 4314 3759 4317
rect 0 4312 3759 4314
rect 0 4256 3698 4312
rect 3754 4256 3759 4312
rect 0 4254 3759 4256
rect 0 4224 480 4254
rect 3693 4251 3759 4254
rect 7005 4314 7071 4317
rect 13721 4314 13787 4317
rect 7005 4312 13787 4314
rect 7005 4256 7010 4312
rect 7066 4256 13726 4312
rect 13782 4256 13787 4312
rect 7005 4254 13787 4256
rect 15702 4314 15762 4526
rect 15886 4450 15946 4662
rect 27520 4632 28000 4662
rect 16113 4586 16179 4589
rect 19517 4586 19583 4589
rect 16113 4584 19583 4586
rect 16113 4528 16118 4584
rect 16174 4528 19522 4584
rect 19578 4528 19583 4584
rect 16113 4526 19583 4528
rect 16113 4523 16179 4526
rect 19517 4523 19583 4526
rect 18229 4450 18295 4453
rect 15886 4448 18295 4450
rect 15886 4392 18234 4448
rect 18290 4392 18295 4448
rect 15886 4390 18295 4392
rect 18229 4387 18295 4390
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 17953 4314 18019 4317
rect 15702 4312 18019 4314
rect 15702 4256 17958 4312
rect 18014 4256 18019 4312
rect 15702 4254 18019 4256
rect 7005 4251 7071 4254
rect 13721 4251 13787 4254
rect 17953 4251 18019 4254
rect 2037 4178 2103 4181
rect 4981 4178 5047 4181
rect 2037 4176 5047 4178
rect 2037 4120 2042 4176
rect 2098 4120 4986 4176
rect 5042 4120 5047 4176
rect 2037 4118 5047 4120
rect 2037 4115 2103 4118
rect 4981 4115 5047 4118
rect 10685 4178 10751 4181
rect 17401 4178 17467 4181
rect 10685 4176 17467 4178
rect 10685 4120 10690 4176
rect 10746 4120 17406 4176
rect 17462 4120 17467 4176
rect 10685 4118 17467 4120
rect 10685 4115 10751 4118
rect 17401 4115 17467 4118
rect 18505 4178 18571 4181
rect 20897 4178 20963 4181
rect 18505 4176 20963 4178
rect 18505 4120 18510 4176
rect 18566 4120 20902 4176
rect 20958 4120 20963 4176
rect 18505 4118 20963 4120
rect 18505 4115 18571 4118
rect 20897 4115 20963 4118
rect 9949 4042 10015 4045
rect 11145 4042 11211 4045
rect 9949 4040 11211 4042
rect 9949 3984 9954 4040
rect 10010 3984 11150 4040
rect 11206 3984 11211 4040
rect 9949 3982 11211 3984
rect 9949 3979 10015 3982
rect 11145 3979 11211 3982
rect 18321 4042 18387 4045
rect 22001 4042 22067 4045
rect 18321 4040 22067 4042
rect 18321 3984 18326 4040
rect 18382 3984 22006 4040
rect 22062 3984 22067 4040
rect 18321 3982 22067 3984
rect 18321 3979 18387 3982
rect 22001 3979 22067 3982
rect 10277 3840 10597 3841
rect 0 3770 480 3800
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 1945 3770 2011 3773
rect 0 3768 2011 3770
rect 0 3712 1950 3768
rect 2006 3712 2011 3768
rect 0 3710 2011 3712
rect 0 3680 480 3710
rect 1945 3707 2011 3710
rect 3969 3770 4035 3773
rect 4429 3770 4495 3773
rect 8109 3772 8175 3773
rect 8109 3770 8156 3772
rect 3969 3768 8156 3770
rect 3969 3712 3974 3768
rect 4030 3712 4434 3768
rect 4490 3712 8114 3768
rect 3969 3710 8156 3712
rect 3969 3707 4035 3710
rect 4429 3707 4495 3710
rect 8109 3708 8156 3710
rect 8220 3708 8226 3772
rect 10869 3770 10935 3773
rect 12893 3770 12959 3773
rect 17585 3770 17651 3773
rect 10734 3768 17651 3770
rect 10734 3712 10874 3768
rect 10930 3712 12898 3768
rect 12954 3712 17590 3768
rect 17646 3712 17651 3768
rect 10734 3710 17651 3712
rect 8109 3707 8175 3708
rect 7189 3634 7255 3637
rect 10734 3634 10794 3710
rect 10869 3707 10935 3710
rect 12893 3707 12959 3710
rect 17585 3707 17651 3710
rect 17718 3708 17724 3772
rect 17788 3770 17794 3772
rect 17861 3770 17927 3773
rect 17788 3768 17927 3770
rect 17788 3712 17866 3768
rect 17922 3712 17927 3768
rect 17788 3710 17927 3712
rect 17788 3708 17794 3710
rect 17861 3707 17927 3710
rect 7189 3632 10794 3634
rect 7189 3576 7194 3632
rect 7250 3576 10794 3632
rect 7189 3574 10794 3576
rect 10961 3634 11027 3637
rect 13445 3634 13511 3637
rect 10961 3632 13511 3634
rect 10961 3576 10966 3632
rect 11022 3576 13450 3632
rect 13506 3576 13511 3632
rect 10961 3574 13511 3576
rect 7189 3571 7255 3574
rect 10961 3571 11027 3574
rect 13445 3571 13511 3574
rect 15101 3634 15167 3637
rect 20897 3634 20963 3637
rect 26509 3634 26575 3637
rect 15101 3632 20963 3634
rect 15101 3576 15106 3632
rect 15162 3576 20902 3632
rect 20958 3576 20963 3632
rect 15101 3574 20963 3576
rect 15101 3571 15167 3574
rect 20897 3571 20963 3574
rect 21038 3632 26575 3634
rect 21038 3576 26514 3632
rect 26570 3576 26575 3632
rect 21038 3574 26575 3576
rect 10133 3498 10199 3501
rect 16941 3498 17007 3501
rect 10133 3496 17007 3498
rect 10133 3440 10138 3496
rect 10194 3440 16946 3496
rect 17002 3440 17007 3496
rect 10133 3438 17007 3440
rect 10133 3435 10199 3438
rect 16941 3435 17007 3438
rect 17769 3498 17835 3501
rect 21038 3498 21098 3574
rect 26509 3571 26575 3574
rect 17769 3496 21098 3498
rect 17769 3440 17774 3496
rect 17830 3440 21098 3496
rect 17769 3438 21098 3440
rect 17769 3435 17835 3438
rect 9121 3362 9187 3365
rect 10961 3362 11027 3365
rect 9121 3360 11027 3362
rect 9121 3304 9126 3360
rect 9182 3304 10966 3360
rect 11022 3304 11027 3360
rect 9121 3302 11027 3304
rect 9121 3299 9187 3302
rect 10961 3299 11027 3302
rect 5610 3296 5930 3297
rect 0 3226 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 4245 3226 4311 3229
rect 0 3224 4311 3226
rect 0 3168 4250 3224
rect 4306 3168 4311 3224
rect 0 3166 4311 3168
rect 0 3136 480 3166
rect 4245 3163 4311 3166
rect 10961 3226 11027 3229
rect 13261 3226 13327 3229
rect 10961 3224 13327 3226
rect 10961 3168 10966 3224
rect 11022 3168 13266 3224
rect 13322 3168 13327 3224
rect 10961 3166 13327 3168
rect 10961 3163 11027 3166
rect 13261 3163 13327 3166
rect 17677 3226 17743 3229
rect 21081 3226 21147 3229
rect 17677 3224 21147 3226
rect 17677 3168 17682 3224
rect 17738 3168 21086 3224
rect 21142 3168 21147 3224
rect 17677 3166 21147 3168
rect 17677 3163 17743 3166
rect 21081 3163 21147 3166
rect 9397 3090 9463 3093
rect 11329 3090 11395 3093
rect 9397 3088 11395 3090
rect 9397 3032 9402 3088
rect 9458 3032 11334 3088
rect 11390 3032 11395 3088
rect 9397 3030 11395 3032
rect 9397 3027 9463 3030
rect 11329 3027 11395 3030
rect 11513 3090 11579 3093
rect 18597 3090 18663 3093
rect 11513 3088 18663 3090
rect 11513 3032 11518 3088
rect 11574 3032 18602 3088
rect 18658 3032 18663 3088
rect 11513 3030 18663 3032
rect 11513 3027 11579 3030
rect 18597 3027 18663 3030
rect 24117 3090 24183 3093
rect 25957 3090 26023 3093
rect 24117 3088 26023 3090
rect 24117 3032 24122 3088
rect 24178 3032 25962 3088
rect 26018 3032 26023 3088
rect 24117 3030 26023 3032
rect 24117 3027 24183 3030
rect 25957 3027 26023 3030
rect 17125 2954 17191 2957
rect 21725 2954 21791 2957
rect 17125 2952 21791 2954
rect 17125 2896 17130 2952
rect 17186 2896 21730 2952
rect 21786 2896 21791 2952
rect 17125 2894 21791 2896
rect 17125 2891 17191 2894
rect 21725 2891 21791 2894
rect 25221 2954 25287 2957
rect 27061 2954 27127 2957
rect 25221 2952 27127 2954
rect 25221 2896 25226 2952
rect 25282 2896 27066 2952
rect 27122 2896 27127 2952
rect 25221 2894 27127 2896
rect 25221 2891 25287 2894
rect 27061 2891 27127 2894
rect 657 2818 723 2821
rect 7005 2818 7071 2821
rect 9673 2818 9739 2821
rect 10133 2818 10199 2821
rect 657 2816 10199 2818
rect 657 2760 662 2816
rect 718 2760 7010 2816
rect 7066 2760 9678 2816
rect 9734 2760 10138 2816
rect 10194 2760 10199 2816
rect 657 2758 10199 2760
rect 657 2755 723 2758
rect 7005 2755 7071 2758
rect 9673 2755 9739 2758
rect 10133 2755 10199 2758
rect 10685 2818 10751 2821
rect 16573 2818 16639 2821
rect 10685 2816 16639 2818
rect 10685 2760 10690 2816
rect 10746 2760 16578 2816
rect 16634 2760 16639 2816
rect 10685 2758 16639 2760
rect 10685 2755 10751 2758
rect 16573 2755 16639 2758
rect 20437 2818 20503 2821
rect 22185 2818 22251 2821
rect 20437 2816 22251 2818
rect 20437 2760 20442 2816
rect 20498 2760 22190 2816
rect 22246 2760 22251 2816
rect 20437 2758 22251 2760
rect 20437 2755 20503 2758
rect 22185 2755 22251 2758
rect 24761 2818 24827 2821
rect 27613 2818 27679 2821
rect 24761 2816 27679 2818
rect 24761 2760 24766 2816
rect 24822 2760 27618 2816
rect 27674 2760 27679 2816
rect 24761 2758 27679 2760
rect 24761 2755 24827 2758
rect 27613 2755 27679 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 2497 2682 2563 2685
rect 5993 2682 6059 2685
rect 2497 2680 6059 2682
rect 2497 2624 2502 2680
rect 2558 2624 5998 2680
rect 6054 2624 6059 2680
rect 2497 2622 6059 2624
rect 2497 2619 2563 2622
rect 5993 2619 6059 2622
rect 0 2546 480 2576
rect 3417 2546 3483 2549
rect 0 2544 3483 2546
rect 0 2488 3422 2544
rect 3478 2488 3483 2544
rect 0 2486 3483 2488
rect 0 2456 480 2486
rect 3417 2483 3483 2486
rect 15469 2546 15535 2549
rect 19517 2546 19583 2549
rect 15469 2544 19583 2546
rect 15469 2488 15474 2544
rect 15530 2488 19522 2544
rect 19578 2488 19583 2544
rect 15469 2486 19583 2488
rect 15469 2483 15535 2486
rect 19517 2483 19583 2486
rect 2129 2410 2195 2413
rect 2957 2410 3023 2413
rect 6361 2410 6427 2413
rect 2129 2408 2882 2410
rect 2129 2352 2134 2408
rect 2190 2352 2882 2408
rect 2129 2350 2882 2352
rect 2129 2347 2195 2350
rect 2822 2138 2882 2350
rect 2957 2408 6427 2410
rect 2957 2352 2962 2408
rect 3018 2352 6366 2408
rect 6422 2352 6427 2408
rect 2957 2350 6427 2352
rect 2957 2347 3023 2350
rect 6361 2347 6427 2350
rect 9949 2410 10015 2413
rect 18505 2410 18571 2413
rect 9949 2408 18571 2410
rect 9949 2352 9954 2408
rect 10010 2352 18510 2408
rect 18566 2352 18571 2408
rect 9949 2350 18571 2352
rect 9949 2347 10015 2350
rect 18505 2347 18571 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 17861 2138 17927 2141
rect 21173 2138 21239 2141
rect 2822 2078 5274 2138
rect 0 2002 480 2032
rect 4889 2002 4955 2005
rect 0 2000 4955 2002
rect 0 1944 4894 2000
rect 4950 1944 4955 2000
rect 0 1942 4955 1944
rect 5214 2002 5274 2078
rect 17861 2136 21239 2138
rect 17861 2080 17866 2136
rect 17922 2080 21178 2136
rect 21234 2080 21239 2136
rect 17861 2078 21239 2080
rect 17861 2075 17927 2078
rect 21173 2075 21239 2078
rect 9765 2002 9831 2005
rect 23933 2002 23999 2005
rect 5214 2000 9831 2002
rect 5214 1944 9770 2000
rect 9826 1944 9831 2000
rect 5214 1942 9831 1944
rect 0 1912 480 1942
rect 4889 1939 4955 1942
rect 9765 1939 9831 1942
rect 9998 2000 23999 2002
rect 9998 1944 23938 2000
rect 23994 1944 23999 2000
rect 9998 1942 23999 1944
rect 3601 1866 3667 1869
rect 9998 1866 10058 1942
rect 23933 1939 23999 1942
rect 3601 1864 10058 1866
rect 3601 1808 3606 1864
rect 3662 1808 10058 1864
rect 3601 1806 10058 1808
rect 3601 1803 3667 1806
rect 10961 1730 11027 1733
rect 17861 1730 17927 1733
rect 10961 1728 17927 1730
rect 10961 1672 10966 1728
rect 11022 1672 17866 1728
rect 17922 1672 17927 1728
rect 10961 1670 17927 1672
rect 10961 1667 11027 1670
rect 17861 1667 17927 1670
rect 18045 1730 18111 1733
rect 19609 1730 19675 1733
rect 18045 1728 19675 1730
rect 18045 1672 18050 1728
rect 18106 1672 19614 1728
rect 19670 1672 19675 1728
rect 18045 1670 19675 1672
rect 18045 1667 18111 1670
rect 19609 1667 19675 1670
rect 3785 1594 3851 1597
rect 3190 1592 3851 1594
rect 3190 1536 3790 1592
rect 3846 1536 3851 1592
rect 3190 1534 3851 1536
rect 0 1458 480 1488
rect 3190 1458 3250 1534
rect 3785 1531 3851 1534
rect 5165 1594 5231 1597
rect 18321 1594 18387 1597
rect 5165 1592 18387 1594
rect 5165 1536 5170 1592
rect 5226 1536 18326 1592
rect 18382 1536 18387 1592
rect 5165 1534 18387 1536
rect 5165 1531 5231 1534
rect 18321 1531 18387 1534
rect 0 1398 3250 1458
rect 11237 1458 11303 1461
rect 18045 1458 18111 1461
rect 11237 1456 18111 1458
rect 11237 1400 11242 1456
rect 11298 1400 18050 1456
rect 18106 1400 18111 1456
rect 11237 1398 18111 1400
rect 0 1368 480 1398
rect 11237 1395 11303 1398
rect 18045 1395 18111 1398
rect 18229 1458 18295 1461
rect 22645 1458 22711 1461
rect 18229 1456 22711 1458
rect 18229 1400 18234 1456
rect 18290 1400 22650 1456
rect 22706 1400 22711 1456
rect 18229 1398 22711 1400
rect 18229 1395 18295 1398
rect 22645 1395 22711 1398
rect 0 914 480 944
rect 6453 914 6519 917
rect 0 912 6519 914
rect 0 856 6458 912
rect 6514 856 6519 912
rect 0 854 6519 856
rect 0 824 480 854
rect 6453 851 6519 854
rect 0 370 480 400
rect 2773 370 2839 373
rect 0 368 2839 370
rect 0 312 2778 368
rect 2834 312 2839 368
rect 0 310 2839 312
rect 0 280 480 310
rect 2773 307 2839 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 2452 17232 2516 17236
rect 2452 17176 2502 17232
rect 2502 17176 2516 17232
rect 2452 17172 2516 17176
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 9628 9556 9692 9620
rect 12940 9556 13004 9620
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 9628 9012 9692 9076
rect 2452 8740 2516 8804
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 9628 7516 9692 7580
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 9628 5340 9692 5404
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 12940 4388 13004 4452
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 8156 3768 8220 3772
rect 8156 3712 8170 3768
rect 8170 3712 8220 3768
rect 8156 3708 8220 3712
rect 17724 3708 17788 3772
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 2451 17236 2517 17237
rect 2451 17172 2452 17236
rect 2516 17172 2517 17236
rect 2451 17171 2517 17172
rect 2454 8805 2514 17171
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 2451 8804 2517 8805
rect 2451 8740 2452 8804
rect 2516 8740 2517 8804
rect 2451 8739 2517 8740
rect 5610 8736 5931 9760
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 9627 9620 9693 9621
rect 9627 9556 9628 9620
rect 9692 9556 9693 9620
rect 9627 9555 9693 9556
rect 9630 9077 9690 9555
rect 10277 9280 10597 10304
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 12939 9620 13005 9621
rect 12939 9556 12940 9620
rect 13004 9556 13005 9620
rect 12939 9555 13005 9556
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 9627 9076 9693 9077
rect 9627 9012 9628 9076
rect 9692 9012 9693 9076
rect 9627 9011 9693 9012
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 9627 7580 9693 7581
rect 9627 7516 9628 7580
rect 9692 7516 9693 7580
rect 9627 7515 9693 7516
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 9630 5405 9690 7515
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 9627 5404 9693 5405
rect 9627 5340 9628 5404
rect 9692 5340 9693 5404
rect 9627 5339 9693 5340
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 12942 4453 13002 9555
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 12939 4452 13005 4453
rect 12939 4388 12940 4452
rect 13004 4388 13005 4452
rect 12939 4387 13005 4388
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 8070 3772 8306 3858
rect 8070 3708 8156 3772
rect 8156 3708 8220 3772
rect 8220 3708 8306 3772
rect 8070 3622 8306 3708
rect 17638 3772 17874 3858
rect 17638 3708 17724 3772
rect 17724 3708 17788 3772
rect 17788 3708 17874 3772
rect 17638 3622 17874 3708
<< metal5 >>
rect 8028 3858 17916 3900
rect 8028 3622 8070 3858
rect 8306 3622 17638 3858
rect 17874 3622 17916 3858
rect 8028 3580 17916 3622
use sky130_fd_sc_hd__fill_2  FILLER_0_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__D tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 1564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_16
timestamp 1604681595
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_12
timestamp 1604681595
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2116 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20
timestamp 1604681595
transform 1 0 2944 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2944 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_29
timestamp 1604681595
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3128 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_33
timestamp 1604681595
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4508 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4324 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51
timestamp 1604681595
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55
timestamp 1604681595
transform 1 0 6164 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6348 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59
timestamp 1604681595
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_69
timestamp 1604681595
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _057_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7176 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_73
timestamp 1604681595
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 8188 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7452 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_93
timestamp 1604681595
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_97
timestamp 1604681595
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1604681595
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1604681595
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10396 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _110_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9844 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12788 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_143
timestamp 1604681595
transform 1 0 14260 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_139
timestamp 1604681595
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_143
timestamp 1604681595
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1604681595
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_163
timestamp 1604681595
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_1_175
timestamp 1604681595
transform 1 0 17204 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_167
timestamp 1604681595
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1604681595
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604681595
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 16836 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_180
timestamp 1604681595
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_181
timestamp 1604681595
transform 1 0 17756 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_177
timestamp 1604681595
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17480 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1604681595
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_193
timestamp 1604681595
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_201 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 19596 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1604681595
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1604681595
transform 1 0 19228 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19044 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19596 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_207
timestamp 1604681595
transform 1 0 20148 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_207
timestamp 1604681595
transform 1 0 20148 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_214
timestamp 1604681595
transform 1 0 20792 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_211
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_218
timestamp 1604681595
transform 1 0 21160 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604681595
transform 1 0 21344 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 21528 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_226
timestamp 1604681595
transform 1 0 21896 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_228
timestamp 1604681595
transform 1 0 22080 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_224
timestamp 1604681595
transform 1 0 21712 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21896 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604681595
transform 1 0 22080 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_236
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604681595
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 22448 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_250
timestamp 1604681595
transform 1 0 24104 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_245
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_242
timestamp 1604681595
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_240 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604681595
transform 1 0 23920 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_230 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 22264 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 24564 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604681595
transform 1 0 25116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_259
timestamp 1604681595
transform 1 0 24932 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_254
timestamp 1604681595
transform 1 0 24472 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_259
timestamp 1604681595
transform 1 0 24932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_263
timestamp 1604681595
transform 1 0 25300 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_271
timestamp 1604681595
transform 1 0 26036 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_275
timestamp 1604681595
transform 1 0 26404 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_36
timestamp 1604681595
transform 1 0 4416 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _069_
timestamp 1604681595
transform 1 0 4140 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_40
timestamp 1604681595
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6716 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6164 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_53
timestamp 1604681595
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_57
timestamp 1604681595
transform 1 0 6348 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1604681595
transform 1 0 8556 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 8004 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_70
timestamp 1604681595
transform 1 0 7544 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_74
timestamp 1604681595
transform 1 0 7912 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_77
timestamp 1604681595
transform 1 0 8188 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9844 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1604681595
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1604681595
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1604681595
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11132 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_105
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_125
timestamp 1604681595
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13340 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_142
timestamp 1604681595
transform 1 0 14168 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15916 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14720 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_146
timestamp 1604681595
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp 1604681595
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_158
timestamp 1604681595
transform 1 0 15640 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17480 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604681595
transform 1 0 16928 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_170
timestamp 1604681595
transform 1 0 16744 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_174
timestamp 1604681595
transform 1 0 17112 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_187
timestamp 1604681595
transform 1 0 18308 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19044 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18492 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18860 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_191
timestamp 1604681595
transform 1 0 18676 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_201
timestamp 1604681595
transform 1 0 19596 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1604681595
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_219
timestamp 1604681595
transform 1 0 21252 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 23920 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_231
timestamp 1604681595
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_243
timestamp 1604681595
transform 1 0 23460 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_247
timestamp 1604681595
transform 1 0 23828 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_252
timestamp 1604681595
transform 1 0 24288 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_264
timestamp 1604681595
transform 1 0 25392 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_272
timestamp 1604681595
transform 1 0 26128 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1564 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_14
timestamp 1604681595
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_18
timestamp 1604681595
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3128 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_38
timestamp 1604681595
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_50
timestamp 1604681595
transform 1 0 5704 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_46
timestamp 1604681595
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_42
timestamp 1604681595
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_55
timestamp 1604681595
transform 1 0 6164 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8464 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_71
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_76
timestamp 1604681595
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1604681595
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_93
timestamp 1604681595
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_97
timestamp 1604681595
transform 1 0 10028 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14076 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_136
timestamp 1604681595
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_140
timestamp 1604681595
transform 1 0 13984 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15364 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_147
timestamp 1604681595
transform 1 0 14628 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_151
timestamp 1604681595
transform 1 0 14996 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_171
timestamp 1604681595
transform 1 0 16836 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_175
timestamp 1604681595
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1604681595
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19596 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1604681595
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1604681595
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_207
timestamp 1604681595
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 21988 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 20884 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604681595
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604681595
transform 1 0 20700 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604681595
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_211
timestamp 1604681595
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_219
timestamp 1604681595
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_223
timestamp 1604681595
transform 1 0 21620 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604681595
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_231
timestamp 1604681595
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_235
timestamp 1604681595
transform 1 0 22724 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_243
timestamp 1604681595
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604681595
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_269
timestamp 1604681595
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_40
timestamp 1604681595
transform 1 0 4784 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_36
timestamp 1604681595
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5520 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_46
timestamp 1604681595
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7544 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_64
timestamp 1604681595
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_72
timestamp 1604681595
transform 1 0 7728 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1604681595
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_88
timestamp 1604681595
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 11224 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_106
timestamp 1604681595
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_119
timestamp 1604681595
transform 1 0 12052 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_125
timestamp 1604681595
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12788 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1604681595
transform 1 0 13616 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_142
timestamp 1604681595
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16008 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14720 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 15456 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_146
timestamp 1604681595
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp 1604681595
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 1604681595
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18216 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_178
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_192
timestamp 1604681595
transform 1 0 18768 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_206
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_219
timestamp 1604681595
transform 1 0 21252 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_231
timestamp 1604681595
transform 1 0 22356 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_243
timestamp 1604681595
transform 1 0 23460 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_255
timestamp 1604681595
transform 1 0 24564 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_267
timestamp 1604681595
transform 1 0 25668 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1932 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_25
timestamp 1604681595
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_29
timestamp 1604681595
transform 1 0 3772 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_33
timestamp 1604681595
transform 1 0 4140 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_36
timestamp 1604681595
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_40
timestamp 1604681595
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1604681595
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604681595
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1604681595
transform 1 0 8556 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1604681595
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_75
timestamp 1604681595
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_79
timestamp 1604681595
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9568 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_84
timestamp 1604681595
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_88
timestamp 1604681595
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_108
timestamp 1604681595
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_112
timestamp 1604681595
transform 1 0 11408 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_132
timestamp 1604681595
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_136
timestamp 1604681595
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16100 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15916 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_149
timestamp 1604681595
transform 1 0 14812 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_153
timestamp 1604681595
transform 1 0 15180 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_159
timestamp 1604681595
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_172
timestamp 1604681595
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_176
timestamp 1604681595
transform 1 0 17296 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_180
timestamp 1604681595
transform 1 0 17664 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 19320 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604681595
transform 1 0 18768 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604681595
transform 1 0 19872 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_190
timestamp 1604681595
transform 1 0 18584 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_194
timestamp 1604681595
transform 1 0 18952 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_202
timestamp 1604681595
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_206
timestamp 1604681595
transform 1 0 20056 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 20516 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604681595
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_210
timestamp 1604681595
transform 1 0 20424 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_215
timestamp 1604681595
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_219
timestamp 1604681595
transform 1 0 21252 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_231
timestamp 1604681595
transform 1 0 22356 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_243
timestamp 1604681595
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604681595
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 1604681595
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1604681595
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_6
timestamp 1604681595
transform 1 0 1656 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _068_
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_11
timestamp 1604681595
transform 1 0 2116 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_10
timestamp 1604681595
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2208 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_29
timestamp 1604681595
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_25
timestamp 1604681595
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_21
timestamp 1604681595
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_40
timestamp 1604681595
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_36
timestamp 1604681595
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4232 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 4140 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_51
timestamp 1604681595
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_47
timestamp 1604681595
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_43
timestamp 1604681595
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5612 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1604681595
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_53
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 5980 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1604681595
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_69
timestamp 1604681595
transform 1 0 7452 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7728 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_79
timestamp 1604681595
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_75
timestamp 1604681595
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_74
timestamp 1604681595
transform 1 0 7912 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1604681595
transform 1 0 8188 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8740 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_88
timestamp 1604681595
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_103
timestamp 1604681595
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_99
timestamp 1604681595
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_102
timestamp 1604681595
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_112
timestamp 1604681595
transform 1 0 11408 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_107
timestamp 1604681595
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_113
timestamp 1604681595
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_106
timestamp 1604681595
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 11224 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1604681595
transform 1 0 11132 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_117
timestamp 1604681595
transform 1 0 11868 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11684 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12788 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13708 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_131
timestamp 1604681595
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_135
timestamp 1604681595
transform 1 0 13524 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_145
timestamp 1604681595
transform 1 0 14444 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_143
timestamp 1604681595
transform 1 0 14260 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14996 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_164
timestamp 1604681595
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_160
timestamp 1604681595
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_161
timestamp 1604681595
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_157
timestamp 1604681595
transform 1 0 15548 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 15732 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16284 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16560 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17296 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_181
timestamp 1604681595
transform 1 0 17756 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_174
timestamp 1604681595
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_178
timestamp 1604681595
transform 1 0 17480 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1604681595
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_187
timestamp 1604681595
transform 1 0 18308 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_191
timestamp 1604681595
transform 1 0 18676 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_193
timestamp 1604681595
transform 1 0 18860 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 18492 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_199
timestamp 1604681595
transform 1 0 19412 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_205
timestamp 1604681595
transform 1 0 19964 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 19596 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_206
timestamp 1604681595
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1604681595
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_210
timestamp 1604681595
transform 1 0 20424 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_222
timestamp 1604681595
transform 1 0 21528 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_234
timestamp 1604681595
transform 1 0 22632 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_242
timestamp 1604681595
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1604681595
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1604681595
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1604681595
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 2944 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2760 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_12
timestamp 1604681595
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_16
timestamp 1604681595
transform 1 0 2576 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4784 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_23
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_35
timestamp 1604681595
transform 1 0 4324 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_39
timestamp 1604681595
transform 1 0 4692 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5428 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_42
timestamp 1604681595
transform 1 0 4968 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7728 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_63
timestamp 1604681595
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_67
timestamp 1604681595
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_71
timestamp 1604681595
transform 1 0 7636 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_81
timestamp 1604681595
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10028 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1604681595
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1604681595
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 12052 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_113
timestamp 1604681595
transform 1 0 11500 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_117
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_121
timestamp 1604681595
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_125
timestamp 1604681595
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15640 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_149
timestamp 1604681595
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17848 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_174
timestamp 1604681595
transform 1 0 17112 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_188
timestamp 1604681595
transform 1 0 18400 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_200
timestamp 1604681595
transform 1 0 19504 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1604681595
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1604681595
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604681595
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2944 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_12
timestamp 1604681595
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_16
timestamp 1604681595
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604681595
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8004 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_65
timestamp 1604681595
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1604681595
transform 1 0 7452 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 10212 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_91
timestamp 1604681595
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_95
timestamp 1604681595
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_102
timestamp 1604681595
transform 1 0 10488 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 12512 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13708 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_127
timestamp 1604681595
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_131
timestamp 1604681595
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_135
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15916 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_153
timestamp 1604681595
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_157
timestamp 1604681595
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_170
timestamp 1604681595
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_174
timestamp 1604681595
transform 1 0 17112 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1604681595
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1604681595
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1604681595
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_19
timestamp 1604681595
transform 1 0 2852 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_36
timestamp 1604681595
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4784 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_60
timestamp 1604681595
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7176 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_64
timestamp 1604681595
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1604681595
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_86
timestamp 1604681595
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1604681595
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_97
timestamp 1604681595
transform 1 0 10028 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_101
timestamp 1604681595
transform 1 0 10396 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1604681595
transform 1 0 10120 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11132 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_107
timestamp 1604681595
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_125
timestamp 1604681595
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13340 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_129
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_142
timestamp 1604681595
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp 1604681595
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_146
timestamp 1604681595
transform 1 0 14536 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14720 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_161
timestamp 1604681595
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 1604681595
transform 1 0 15640 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1604681595
transform 1 0 16008 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1604681595
transform 1 0 16284 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1604681595
transform 1 0 17388 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_189
timestamp 1604681595
transform 1 0 18492 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1604681595
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1604681595
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604681595
transform 1 0 4140 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_25
timestamp 1604681595
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_29
timestamp 1604681595
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_36
timestamp 1604681595
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_40
timestamp 1604681595
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1604681595
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 8372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_71
timestamp 1604681595
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_75
timestamp 1604681595
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_82
timestamp 1604681595
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8832 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10396 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_93
timestamp 1604681595
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_97
timestamp 1604681595
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11868 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1604681595
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1604681595
transform 1 0 13984 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14444 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_132
timestamp 1604681595
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_136
timestamp 1604681595
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_143
timestamp 1604681595
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_147
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp 1604681595
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_175
timestamp 1604681595
transform 1 0 17204 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604681595
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1472 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_13
timestamp 1604681595
transform 1 0 2300 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_17
timestamp 1604681595
transform 1 0 2668 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_21
timestamp 1604681595
transform 1 0 3036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_25
timestamp 1604681595
transform 1 0 3404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_38
timestamp 1604681595
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 5336 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_42
timestamp 1604681595
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1604681595
transform 1 0 6808 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 7728 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_68
timestamp 1604681595
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_88
timestamp 1604681595
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_97
timestamp 1604681595
transform 1 0 10028 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1604681595
transform 1 0 9752 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_103
timestamp 1604681595
transform 1 0 10580 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_121
timestamp 1604681595
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_125
timestamp 1604681595
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12972 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1604681595
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_142
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_150
timestamp 1604681595
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1604681595
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1604681595
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604681595
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_8
timestamp 1604681595
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2024 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_19
timestamp 1604681595
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1840 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_28
timestamp 1604681595
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_24
timestamp 1604681595
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4048 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_41
timestamp 1604681595
transform 1 0 4876 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_45
timestamp 1604681595
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_45
timestamp 1604681595
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5060 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5612 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 5612 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_58
timestamp 1604681595
transform 1 0 6440 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_60
timestamp 1604681595
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_56
timestamp 1604681595
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_52
timestamp 1604681595
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6716 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7544 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7544 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_66
timestamp 1604681595
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_79
timestamp 1604681595
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_83
timestamp 1604681595
transform 1 0 8740 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_89
timestamp 1604681595
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_90
timestamp 1604681595
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_86
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_101
timestamp 1604681595
transform 1 0 10396 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_97
timestamp 1604681595
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_94
timestamp 1604681595
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10948 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604681595
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_106
timestamp 1604681595
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_123
timestamp 1604681595
transform 1 0 12420 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_133
timestamp 1604681595
transform 1 0 13340 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_129
timestamp 1604681595
transform 1 0 12972 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1604681595
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13524 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_136
timestamp 1604681595
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_137
timestamp 1604681595
transform 1 0 13708 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_140
timestamp 1604681595
transform 1 0 13984 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_152
timestamp 1604681595
transform 1 0 15088 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_164
timestamp 1604681595
transform 1 0 16192 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1604681595
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1604681595
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_176
timestamp 1604681595
transform 1 0 17296 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1604681595
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1604681595
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1604681595
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1604681595
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_220
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_232
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1604681595
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604681595
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1604681595
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4232 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_23
timestamp 1604681595
transform 1 0 3220 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_27
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1604681595
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_50
timestamp 1604681595
transform 1 0 5704 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_54
timestamp 1604681595
transform 1 0 6072 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_58
timestamp 1604681595
transform 1 0 6440 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7820 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_66
timestamp 1604681595
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_69
timestamp 1604681595
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_82
timestamp 1604681595
transform 1 0 8648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10672 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9108 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_96
timestamp 1604681595
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_100
timestamp 1604681595
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1604681595
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_117
timestamp 1604681595
transform 1 0 11868 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1604681595
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_140
timestamp 1604681595
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_144
timestamp 1604681595
transform 1 0 14352 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_156
timestamp 1604681595
transform 1 0 15456 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_168
timestamp 1604681595
transform 1 0 16560 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_180
timestamp 1604681595
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1604681595
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_232
timestamp 1604681595
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1604681595
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1604681595
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1656 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_22
timestamp 1604681595
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_26
timestamp 1604681595
transform 1 0 3496 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_41
timestamp 1604681595
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5612 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_46
timestamp 1604681595
transform 1 0 5336 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7820 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_65
timestamp 1604681595
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_69
timestamp 1604681595
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_89
timestamp 1604681595
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_102
timestamp 1604681595
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11224 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11040 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_106
timestamp 1604681595
transform 1 0 10856 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_119
timestamp 1604681595
transform 1 0 12052 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_125
timestamp 1604681595
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12788 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_136
timestamp 1604681595
transform 1 0 13616 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_148
timestamp 1604681595
transform 1 0 14720 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1604681595
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1604681595
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_190
timestamp 1604681595
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1604681595
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1604681595
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1604681595
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2668 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_9
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_13
timestamp 1604681595
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4508 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_26
timestamp 1604681595
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_30
timestamp 1604681595
transform 1 0 3864 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_34
timestamp 1604681595
transform 1 0 4232 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_53
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604681595
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_65
timestamp 1604681595
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1604681595
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_73
timestamp 1604681595
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_77
timestamp 1604681595
transform 1 0 8188 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_81
timestamp 1604681595
transform 1 0 8556 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10672 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8832 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12604 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13340 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_127
timestamp 1604681595
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_131
timestamp 1604681595
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_135
timestamp 1604681595
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1604681595
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_143
timestamp 1604681595
transform 1 0 14260 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_155
timestamp 1604681595
transform 1 0 15364 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_167
timestamp 1604681595
transform 1 0 16468 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1604681595
transform 1 0 17572 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1604681595
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1604681595
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604681595
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_226
timestamp 1604681595
transform 1 0 21896 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_238
timestamp 1604681595
transform 1 0 23000 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1472 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_13
timestamp 1604681595
transform 1 0 2300 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_19
timestamp 1604681595
transform 1 0 2852 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3036 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_40
timestamp 1604681595
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_36
timestamp 1604681595
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604681595
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5520 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_47
timestamp 1604681595
transform 1 0 5428 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_64
timestamp 1604681595
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_68
timestamp 1604681595
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_72
timestamp 1604681595
transform 1 0 7728 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_88
timestamp 1604681595
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11960 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_109
timestamp 1604681595
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_113
timestamp 1604681595
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_117
timestamp 1604681595
transform 1 0 11868 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_134
timestamp 1604681595
transform 1 0 13432 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_146
timestamp 1604681595
transform 1 0 14536 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1604681595
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1604681595
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1604681595
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1604681595
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 21712 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_223
timestamp 1604681595
transform 1 0 21620 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_228
timestamp 1604681595
transform 1 0 22080 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_240
timestamp 1604681595
transform 1 0 23184 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_252
timestamp 1604681595
transform 1 0 24288 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_264
timestamp 1604681595
transform 1 0 25392 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_272
timestamp 1604681595
transform 1 0 26128 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1472 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_17
timestamp 1604681595
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_13
timestamp 1604681595
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1748 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_40
timestamp 1604681595
transform 1 0 4784 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_36
timestamp 1604681595
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_41
timestamp 1604681595
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_37
timestamp 1604681595
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3036 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_19_49
timestamp 1604681595
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604681595
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 5244 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_62
timestamp 1604681595
transform 1 0 6808 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5336 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_20_67
timestamp 1604681595
transform 1 0 7268 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7544 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 7084 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_79
timestamp 1604681595
transform 1 0 8372 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_82
timestamp 1604681595
transform 1 0 8648 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_78
timestamp 1604681595
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_74
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 8740 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1604681595
transform 1 0 8924 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_90
timestamp 1604681595
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_86
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 9108 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10028 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10212 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9752 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1604681595
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_115
timestamp 1604681595
transform 1 0 11684 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_119
timestamp 1604681595
transform 1 0 12052 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11868 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_123
timestamp 1604681595
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1604681595
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_127
timestamp 1604681595
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_131
timestamp 1604681595
transform 1 0 13156 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_143
timestamp 1604681595
transform 1 0 14260 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_127
timestamp 1604681595
transform 1 0 12788 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_139
timestamp 1604681595
transform 1 0 13892 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_155
timestamp 1604681595
transform 1 0 15364 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1604681595
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_167
timestamp 1604681595
transform 1 0 16468 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1604681595
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1604681595
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1604681595
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_220
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_228
timestamp 1604681595
transform 1 0 22080 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 22264 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604681595
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_232
timestamp 1604681595
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_234
timestamp 1604681595
transform 1 0 22632 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_246
timestamp 1604681595
transform 1 0 23736 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1604681595
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_258
timestamp 1604681595
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_270
timestamp 1604681595
transform 1 0 25944 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_274
timestamp 1604681595
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1932 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 4140 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_25
timestamp 1604681595
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_29
timestamp 1604681595
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_36
timestamp 1604681595
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1604681595
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7820 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_65
timestamp 1604681595
transform 1 0 7084 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1604681595
transform 1 0 7452 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10028 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_89
timestamp 1604681595
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_93
timestamp 1604681595
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_106
timestamp 1604681595
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1604681595
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_126
timestamp 1604681595
transform 1 0 12696 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_130
timestamp 1604681595
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_134
timestamp 1604681595
transform 1 0 13432 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_146
timestamp 1604681595
transform 1 0 14536 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_158
timestamp 1604681595
transform 1 0 15640 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_170
timestamp 1604681595
transform 1 0 16744 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1604681595
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_232
timestamp 1604681595
transform 1 0 22448 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_249
timestamp 1604681595
transform 1 0 24012 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604681595
transform 1 0 24196 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_253
timestamp 1604681595
transform 1 0 24380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_265
timestamp 1604681595
transform 1 0 25484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_6
timestamp 1604681595
transform 1 0 1656 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_12
timestamp 1604681595
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_36
timestamp 1604681595
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_40
timestamp 1604681595
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4968 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_58
timestamp 1604681595
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_62
timestamp 1604681595
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7176 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 8740 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6992 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_75
timestamp 1604681595
transform 1 0 8004 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_79
timestamp 1604681595
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10212 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_86
timestamp 1604681595
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1604681595
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_98
timestamp 1604681595
transform 1 0 10120 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_115
timestamp 1604681595
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_119
timestamp 1604681595
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_132
timestamp 1604681595
transform 1 0 13248 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_144
timestamp 1604681595
transform 1 0 14352 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1604681595
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 23460 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_239
timestamp 1604681595
transform 1 0 23092 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_247
timestamp 1604681595
transform 1 0 23828 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_259
timestamp 1604681595
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1604681595
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2024 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1604681595
transform 1 0 1748 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_19
timestamp 1604681595
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_23
timestamp 1604681595
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_36
timestamp 1604681595
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_40
timestamp 1604681595
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7728 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_66
timestamp 1604681595
transform 1 0 7176 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_69
timestamp 1604681595
transform 1 0 7452 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9936 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_88
timestamp 1604681595
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_92
timestamp 1604681595
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_113
timestamp 1604681595
transform 1 0 11500 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_109
timestamp 1604681595
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_105
timestamp 1604681595
transform 1 0 10764 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 10948 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_132
timestamp 1604681595
transform 1 0 13248 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_144
timestamp 1604681595
transform 1 0 14352 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_156
timestamp 1604681595
transform 1 0 15456 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_168
timestamp 1604681595
transform 1 0 16560 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1604681595
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604681595
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604681595
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_269
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_6
timestamp 1604681595
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_10
timestamp 1604681595
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_35
timestamp 1604681595
transform 1 0 4324 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_39
timestamp 1604681595
transform 1 0 4692 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4508 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5060 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 6716 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_59
timestamp 1604681595
transform 1 0 6532 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7268 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_63
timestamp 1604681595
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_76
timestamp 1604681595
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_80
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10304 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 9108 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9936 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_84
timestamp 1604681595
transform 1 0 8832 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1604681595
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_98
timestamp 1604681595
transform 1 0 10120 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_116
timestamp 1604681595
transform 1 0 11776 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_120
timestamp 1604681595
transform 1 0 12144 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_125
timestamp 1604681595
transform 1 0 12604 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_137
timestamp 1604681595
transform 1 0 13708 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1604681595
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604681595
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1604681595
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1604681595
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1604681595
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2760 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_9
timestamp 1604681595
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_13
timestamp 1604681595
transform 1 0 2300 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_34
timestamp 1604681595
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_38
timestamp 1604681595
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5060 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6440 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_42
timestamp 1604681595
transform 1 0 4968 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_52
timestamp 1604681595
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_56
timestamp 1604681595
transform 1 0 6256 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_60
timestamp 1604681595
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7360 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7176 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10212 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_84
timestamp 1604681595
transform 1 0 8832 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_88
timestamp 1604681595
transform 1 0 9200 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_91
timestamp 1604681595
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_95
timestamp 1604681595
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_108
timestamp 1604681595
transform 1 0 11040 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_112
timestamp 1604681595
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_116
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_126
timestamp 1604681595
transform 1 0 12696 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_138
timestamp 1604681595
transform 1 0 13800 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_150
timestamp 1604681595
transform 1 0 14904 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_162
timestamp 1604681595
transform 1 0 16008 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_174
timestamp 1604681595
transform 1 0 17112 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1604681595
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604681595
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1604681595
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1604681595
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_9
timestamp 1604681595
transform 1 0 1932 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1656 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_16
timestamp 1604681595
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_13
timestamp 1604681595
transform 1 0 2300 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_19
timestamp 1604681595
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2760 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1604681595
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_34
timestamp 1604681595
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_41
timestamp 1604681595
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_49
timestamp 1604681595
transform 1 0 5612 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_45
timestamp 1604681595
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4968 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_55
timestamp 1604681595
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5796 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_67
timestamp 1604681595
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_71
timestamp 1604681595
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_78
timestamp 1604681595
transform 1 0 8280 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_82
timestamp 1604681595
transform 1 0 8648 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_84
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_88
timestamp 1604681595
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 9292 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_92
timestamp 1604681595
transform 1 0 9568 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_102
timestamp 1604681595
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10672 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9936 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1604681595
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_106
timestamp 1604681595
transform 1 0 10856 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1604681595
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_117
timestamp 1604681595
transform 1 0 11868 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_124
timestamp 1604681595
transform 1 0 12512 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_112
timestamp 1604681595
transform 1 0 11408 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_136
timestamp 1604681595
transform 1 0 13616 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1604681595
transform 1 0 14720 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1604681595
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1604681595
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1604681595
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1604681595
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1604681595
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1604681595
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604681595
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604681595
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1604681595
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1604681595
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_6
timestamp 1604681595
transform 1 0 1656 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_11
timestamp 1604681595
transform 1 0 2116 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5704 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6072 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_48
timestamp 1604681595
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_52
timestamp 1604681595
transform 1 0 5888 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 8556 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8280 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_72
timestamp 1604681595
transform 1 0 7728 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_76
timestamp 1604681595
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_80
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9752 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9292 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_88
timestamp 1604681595
transform 1 0 9200 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1604681595
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_110
timestamp 1604681595
transform 1 0 11224 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_122
timestamp 1604681595
transform 1 0 12328 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_134
timestamp 1604681595
transform 1 0 13432 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_146
timestamp 1604681595
transform 1 0 14536 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1604681595
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604681595
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1604681595
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1932 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_18
timestamp 1604681595
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_22
timestamp 1604681595
transform 1 0 3128 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_36
timestamp 1604681595
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_40
timestamp 1604681595
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1604681595
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7176 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_75
timestamp 1604681595
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_79
timestamp 1604681595
transform 1 0 8372 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9292 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_85
timestamp 1604681595
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10948 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11316 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_105
timestamp 1604681595
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_109
timestamp 1604681595
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1604681595
transform 1 0 11500 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1604681595
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1604681595
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1604681595
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1604681595
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1604681595
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1932 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1604681595
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_22
timestamp 1604681595
transform 1 0 3128 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_26
timestamp 1604681595
transform 1 0 3496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_36
timestamp 1604681595
transform 1 0 4416 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_40
timestamp 1604681595
transform 1 0 4784 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5244 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_43
timestamp 1604681595
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_61
timestamp 1604681595
transform 1 0 6716 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7452 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 8464 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_65
timestamp 1604681595
transform 1 0 7084 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_78
timestamp 1604681595
transform 1 0 8280 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1604681595
transform 1 0 8648 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_86
timestamp 1604681595
transform 1 0 9016 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1604681595
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_106
timestamp 1604681595
transform 1 0 10856 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_118
timestamp 1604681595
transform 1 0 11960 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_130
timestamp 1604681595
transform 1 0 13064 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_142
timestamp 1604681595
transform 1 0 14168 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_150
timestamp 1604681595
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1604681595
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1604681595
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604681595
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2852 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1604681595
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 4140 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3956 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_25
timestamp 1604681595
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_29
timestamp 1604681595
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_36
timestamp 1604681595
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_40
timestamp 1604681595
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_53
timestamp 1604681595
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604681595
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8372 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_71
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_75
timestamp 1604681595
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_95
timestamp 1604681595
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_99
timestamp 1604681595
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_112
timestamp 1604681595
transform 1 0 11408 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1604681595
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1604681595
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604681595
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604681595
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1604681595
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2668 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_9
timestamp 1604681595
transform 1 0 1932 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_13
timestamp 1604681595
transform 1 0 2300 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1604681595
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_40
timestamp 1604681595
transform 1 0 4784 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_36
timestamp 1604681595
transform 1 0 4416 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 4600 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604681595
transform 1 0 4232 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4876 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5888 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_50
timestamp 1604681595
transform 1 0 5704 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_54
timestamp 1604681595
transform 1 0 6072 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_58
timestamp 1604681595
transform 1 0 6440 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_64
timestamp 1604681595
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_88
timestamp 1604681595
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1604681595
transform 1 0 11132 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1604681595
transform 1 0 12236 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_133
timestamp 1604681595
transform 1 0 13340 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_145
timestamp 1604681595
transform 1 0 14444 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1604681595
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1604681595
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1604681595
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1604681595
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1604681595
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1604681595
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_16
timestamp 1604681595
transform 1 0 2576 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_12
timestamp 1604681595
transform 1 0 2208 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2392 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2944 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_12
timestamp 1604681595
transform 1 0 2208 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_30
timestamp 1604681595
transform 1 0 3864 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_24
timestamp 1604681595
transform 1 0 3312 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_30
timestamp 1604681595
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_26
timestamp 1604681595
transform 1 0 3496 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3680 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_40
timestamp 1604681595
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4140 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4232 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_39
timestamp 1604681595
transform 1 0 4692 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_51
timestamp 1604681595
transform 1 0 5796 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_52
timestamp 1604681595
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_44
timestamp 1604681595
transform 1 0 5152 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 5336 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 5520 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_60
timestamp 1604681595
transform 1 0 6624 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_56
timestamp 1604681595
transform 1 0 6256 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604681595
transform 1 0 6072 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6072 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 8464 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_78
timestamp 1604681595
transform 1 0 8280 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_82
timestamp 1604681595
transform 1 0 8648 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_64
timestamp 1604681595
transform 1 0 6992 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_71
timestamp 1604681595
transform 1 0 7636 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_83
timestamp 1604681595
transform 1 0 8740 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1604681595
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_90
timestamp 1604681595
transform 1 0 9384 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_99
timestamp 1604681595
transform 1 0 10212 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_95
timestamp 1604681595
transform 1 0 9844 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_102
timestamp 1604681595
transform 1 0 10488 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_103
timestamp 1604681595
transform 1 0 10580 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_115
timestamp 1604681595
transform 1 0 11684 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1604681595
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_114
timestamp 1604681595
transform 1 0 11592 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1604681595
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_126
timestamp 1604681595
transform 1 0 12696 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_138
timestamp 1604681595
transform 1 0 13800 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1604681595
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_159
timestamp 1604681595
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_150
timestamp 1604681595
transform 1 0 14904 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_171
timestamp 1604681595
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604681595
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604681595
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1604681595
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1604681595
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604681595
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 2852 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_11
timestamp 1604681595
transform 1 0 2116 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_17
timestamp 1604681595
transform 1 0 2668 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 3956 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604681595
transform 1 0 3404 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604681595
transform 1 0 4508 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604681595
transform 1 0 4876 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_23
timestamp 1604681595
transform 1 0 3220 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_35
timestamp 1604681595
transform 1 0 4324 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_39
timestamp 1604681595
transform 1 0 4692 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 5060 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604681595
transform 1 0 5612 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604681595
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_47
timestamp 1604681595
transform 1 0 5428 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_51
timestamp 1604681595
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_55
timestamp 1604681595
transform 1 0 6164 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 7912 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8648 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 7728 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_70
timestamp 1604681595
transform 1 0 7544 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_80
timestamp 1604681595
transform 1 0 8464 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 9200 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_84
timestamp 1604681595
transform 1 0 8832 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_91
timestamp 1604681595
transform 1 0 9476 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_103
timestamp 1604681595
transform 1 0 10580 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_115
timestamp 1604681595
transform 1 0 11684 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_121
timestamp 1604681595
transform 1 0 12236 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_135
timestamp 1604681595
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_147
timestamp 1604681595
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_159
timestamp 1604681595
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_171
timestamp 1604681595
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604681595
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604681595
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1604681595
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1604681595
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1604681595
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 2484 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604681595
transform 1 0 2300 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_7
timestamp 1604681595
transform 1 0 1748 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_11
timestamp 1604681595
transform 1 0 2116 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_19
timestamp 1604681595
transform 1 0 2852 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_36
timestamp 1604681595
transform 1 0 4416 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 5428 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_44
timestamp 1604681595
transform 1 0 5152 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_51
timestamp 1604681595
transform 1 0 5796 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8096 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_63
timestamp 1604681595
transform 1 0 6900 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_75
timestamp 1604681595
transform 1 0 8004 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_82
timestamp 1604681595
transform 1 0 8648 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_90
timestamp 1604681595
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1604681595
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_117
timestamp 1604681595
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1604681595
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1604681595
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_166
timestamp 1604681595
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_178
timestamp 1604681595
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_190
timestamp 1604681595
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_202
timestamp 1604681595
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604681595
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1604681595
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1604681595
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1604681595
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 2944 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2392 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2760 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_12
timestamp 1604681595
transform 1 0 2208 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_16
timestamp 1604681595
transform 1 0 2576 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 4048 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604681595
transform 1 0 3496 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604681595
transform 1 0 4600 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_24
timestamp 1604681595
transform 1 0 3312 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_28
timestamp 1604681595
transform 1 0 3680 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_36
timestamp 1604681595
transform 1 0 4416 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_40
timestamp 1604681595
transform 1 0 4784 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_52
timestamp 1604681595
transform 1 0 5888 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_60
timestamp 1604681595
transform 1 0 6624 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 7268 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8740 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604681595
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604681595
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_66
timestamp 1604681595
transform 1 0 7176 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_71
timestamp 1604681595
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_75
timestamp 1604681595
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_79
timestamp 1604681595
transform 1 0 8372 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9476 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_89
timestamp 1604681595
transform 1 0 9292 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1604681595
transform 1 0 9660 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_105
timestamp 1604681595
transform 1 0 10764 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_117
timestamp 1604681595
transform 1 0 11868 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_121
timestamp 1604681595
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_135
timestamp 1604681595
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_147
timestamp 1604681595
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_159
timestamp 1604681595
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_171
timestamp 1604681595
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1604681595
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1604681595
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_220
timestamp 1604681595
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_232
timestamp 1604681595
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1604681595
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1604681595
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_12
timestamp 1604681595
transform 1 0 2208 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_24
timestamp 1604681595
transform 1 0 3312 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_30
timestamp 1604681595
transform 1 0 3864 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604681595
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604681595
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 8096 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_68
timestamp 1604681595
transform 1 0 7360 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1604681595
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1604681595
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_117
timestamp 1604681595
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_129
timestamp 1604681595
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1604681595
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1604681595
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_178
timestamp 1604681595
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_190
timestamp 1604681595
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_202
timestamp 1604681595
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1604681595
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1604681595
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_251
timestamp 1604681595
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_263
timestamp 1604681595
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_7
timestamp 1604681595
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604681595
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_19
timestamp 1604681595
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_11
timestamp 1604681595
transform 1 0 2116 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604681595
transform 1 0 2300 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_19
timestamp 1604681595
transform 1 0 2852 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_7
timestamp 1604681595
transform 1 0 1748 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604681595
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604681595
transform 1 0 4140 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_23
timestamp 1604681595
transform 1 0 3220 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_31
timestamp 1604681595
transform 1 0 3956 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1604681595
transform 1 0 4324 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_47
timestamp 1604681595
transform 1 0 5428 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604681595
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1604681595
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1604681595
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1604681595
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_98
timestamp 1604681595
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_110
timestamp 1604681595
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1604681595
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_117
timestamp 1604681595
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_135
timestamp 1604681595
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1604681595
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1604681595
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_147
timestamp 1604681595
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_159
timestamp 1604681595
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_166
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_171
timestamp 1604681595
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1604681595
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 19780 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_196
timestamp 1604681595
transform 1 0 19136 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_202
timestamp 1604681595
transform 1 0 19688 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_207
timestamp 1604681595
transform 1 0 20148 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_190
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_202
timestamp 1604681595
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_219
timestamp 1604681595
transform 1 0 21252 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1604681595
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_231
timestamp 1604681595
transform 1 0 22356 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_243
timestamp 1604681595
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1604681595
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_257
timestamp 1604681595
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1604681595
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_251
timestamp 1604681595
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_263
timestamp 1604681595
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1604681595
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1604681595
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1604681595
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_147
timestamp 1604681595
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_159
timestamp 1604681595
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_171
timestamp 1604681595
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604681595
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604681595
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604681595
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604681595
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604681595
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604681595
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604681595
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604681595
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604681595
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604681595
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604681595
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604681595
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604681595
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604681595
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 27066 0 27122 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 7010 27520 7066 28000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 27618 0 27674 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 20994 27520 21050 28000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 4 nsew default input
rlabel metal2 s 662 0 718 480 6 bottom_left_grid_pin_43_
port 5 nsew default input
rlabel metal2 s 1214 0 1270 480 6 bottom_left_grid_pin_44_
port 6 nsew default input
rlabel metal2 s 1766 0 1822 480 6 bottom_left_grid_pin_45_
port 7 nsew default input
rlabel metal2 s 2318 0 2374 480 6 bottom_left_grid_pin_46_
port 8 nsew default input
rlabel metal2 s 2870 0 2926 480 6 bottom_left_grid_pin_47_
port 9 nsew default input
rlabel metal2 s 3422 0 3478 480 6 bottom_left_grid_pin_48_
port 10 nsew default input
rlabel metal2 s 3974 0 4030 480 6 bottom_left_grid_pin_49_
port 11 nsew default input
rlabel metal2 s 26514 0 26570 480 6 bottom_right_grid_pin_1_
port 12 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 ccff_head
port 13 nsew default input
rlabel metal3 s 27520 23264 28000 23384 6 ccff_tail
port 14 nsew default tristate
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[0]
port 15 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[10]
port 16 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[11]
port 17 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[12]
port 18 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[13]
port 19 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[14]
port 20 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[15]
port 21 nsew default input
rlabel metal3 s 0 13880 480 14000 6 chanx_left_in[16]
port 22 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[17]
port 23 nsew default input
rlabel metal3 s 0 15104 480 15224 6 chanx_left_in[18]
port 24 nsew default input
rlabel metal3 s 0 15648 480 15768 6 chanx_left_in[19]
port 25 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[1]
port 26 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[2]
port 27 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[3]
port 28 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[4]
port 29 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[5]
port 30 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[6]
port 31 nsew default input
rlabel metal3 s 0 8848 480 8968 6 chanx_left_in[7]
port 32 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[8]
port 33 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[9]
port 34 nsew default input
rlabel metal3 s 0 16192 480 16312 6 chanx_left_out[0]
port 35 nsew default tristate
rlabel metal3 s 0 21904 480 22024 6 chanx_left_out[10]
port 36 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[11]
port 37 nsew default tristate
rlabel metal3 s 0 23128 480 23248 6 chanx_left_out[12]
port 38 nsew default tristate
rlabel metal3 s 0 23672 480 23792 6 chanx_left_out[13]
port 39 nsew default tristate
rlabel metal3 s 0 24216 480 24336 6 chanx_left_out[14]
port 40 nsew default tristate
rlabel metal3 s 0 24760 480 24880 6 chanx_left_out[15]
port 41 nsew default tristate
rlabel metal3 s 0 25304 480 25424 6 chanx_left_out[16]
port 42 nsew default tristate
rlabel metal3 s 0 25984 480 26104 6 chanx_left_out[17]
port 43 nsew default tristate
rlabel metal3 s 0 26528 480 26648 6 chanx_left_out[18]
port 44 nsew default tristate
rlabel metal3 s 0 27072 480 27192 6 chanx_left_out[19]
port 45 nsew default tristate
rlabel metal3 s 0 16736 480 16856 6 chanx_left_out[1]
port 46 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 chanx_left_out[2]
port 47 nsew default tristate
rlabel metal3 s 0 17960 480 18080 6 chanx_left_out[3]
port 48 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[4]
port 49 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[5]
port 50 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chanx_left_out[6]
port 51 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[7]
port 52 nsew default tristate
rlabel metal3 s 0 20816 480 20936 6 chanx_left_out[8]
port 53 nsew default tristate
rlabel metal3 s 0 21360 480 21480 6 chanx_left_out[9]
port 54 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_in[0]
port 55 nsew default input
rlabel metal2 s 10046 0 10102 480 6 chany_bottom_in[10]
port 56 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[11]
port 57 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_in[12]
port 58 nsew default input
rlabel metal2 s 11702 0 11758 480 6 chany_bottom_in[13]
port 59 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[14]
port 60 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_in[15]
port 61 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[16]
port 62 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[17]
port 63 nsew default input
rlabel metal2 s 14370 0 14426 480 6 chany_bottom_in[18]
port 64 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[19]
port 65 nsew default input
rlabel metal2 s 5078 0 5134 480 6 chany_bottom_in[1]
port 66 nsew default input
rlabel metal2 s 5630 0 5686 480 6 chany_bottom_in[2]
port 67 nsew default input
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_in[3]
port 68 nsew default input
rlabel metal2 s 6734 0 6790 480 6 chany_bottom_in[4]
port 69 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chany_bottom_in[5]
port 70 nsew default input
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_in[6]
port 71 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[7]
port 72 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[8]
port 73 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[9]
port 74 nsew default input
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_out[0]
port 75 nsew default tristate
rlabel metal2 s 20994 0 21050 480 6 chany_bottom_out[10]
port 76 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[11]
port 77 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[12]
port 78 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[13]
port 79 nsew default tristate
rlabel metal2 s 23202 0 23258 480 6 chany_bottom_out[14]
port 80 nsew default tristate
rlabel metal2 s 23754 0 23810 480 6 chany_bottom_out[15]
port 81 nsew default tristate
rlabel metal2 s 24306 0 24362 480 6 chany_bottom_out[16]
port 82 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 chany_bottom_out[17]
port 83 nsew default tristate
rlabel metal2 s 25410 0 25466 480 6 chany_bottom_out[18]
port 84 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_bottom_out[19]
port 85 nsew default tristate
rlabel metal2 s 16026 0 16082 480 6 chany_bottom_out[1]
port 86 nsew default tristate
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_out[2]
port 87 nsew default tristate
rlabel metal2 s 17130 0 17186 480 6 chany_bottom_out[3]
port 88 nsew default tristate
rlabel metal2 s 17682 0 17738 480 6 chany_bottom_out[4]
port 89 nsew default tristate
rlabel metal2 s 18234 0 18290 480 6 chany_bottom_out[5]
port 90 nsew default tristate
rlabel metal2 s 18786 0 18842 480 6 chany_bottom_out[6]
port 91 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chany_bottom_out[7]
port 92 nsew default tristate
rlabel metal2 s 19890 0 19946 480 6 chany_bottom_out[8]
port 93 nsew default tristate
rlabel metal2 s 20442 0 20498 480 6 chany_bottom_out[9]
port 94 nsew default tristate
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_34_
port 95 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_35_
port 96 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_36_
port 97 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_37_
port 98 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_38_
port 99 nsew default input
rlabel metal3 s 0 3136 480 3256 6 left_bottom_grid_pin_39_
port 100 nsew default input
rlabel metal3 s 0 3680 480 3800 6 left_bottom_grid_pin_40_
port 101 nsew default input
rlabel metal3 s 0 4224 480 4344 6 left_bottom_grid_pin_41_
port 102 nsew default input
rlabel metal3 s 0 27616 480 27736 6 left_top_grid_pin_1_
port 103 nsew default input
rlabel metal3 s 27520 4632 28000 4752 6 prog_clk
port 104 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 105 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 106 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
