magic
tech sky130A
magscale 1 2
timestamp 1605197775
<< locali >>
rect 6929 18471 6963 18573
<< viali >>
rect 11621 20409 11655 20443
rect 13001 20341 13035 20375
rect 7849 20273 7883 20307
rect 10425 20273 10459 20307
rect 13553 20273 13587 20307
rect 16589 20273 16623 20307
rect 11437 20205 11471 20239
rect 18337 20205 18371 20239
rect 19993 20205 20027 20239
rect 7665 20137 7699 20171
rect 16405 20137 16439 20171
rect 18613 20137 18647 20171
rect 7205 20069 7239 20103
rect 7573 20069 7607 20103
rect 13369 20069 13403 20103
rect 13461 20069 13495 20103
rect 16037 20069 16071 20103
rect 16497 20069 16531 20103
rect 20177 20069 20211 20103
rect 16037 19865 16071 19899
rect 7104 19729 7138 19763
rect 9393 19729 9427 19763
rect 13625 19729 13659 19763
rect 15945 19729 15979 19763
rect 18061 19729 18095 19763
rect 19809 19729 19843 19763
rect 6837 19661 6871 19695
rect 9137 19661 9171 19695
rect 11345 19661 11379 19695
rect 13369 19661 13403 19695
rect 16129 19661 16163 19695
rect 18245 19661 18279 19695
rect 19993 19661 20027 19695
rect 15577 19593 15611 19627
rect 8217 19525 8251 19559
rect 10517 19525 10551 19559
rect 14749 19525 14783 19559
rect 8769 19321 8803 19355
rect 13277 19321 13311 19355
rect 17969 19253 18003 19287
rect 19073 19185 19107 19219
rect 6377 19117 6411 19151
rect 7389 19117 7423 19151
rect 7656 19117 7690 19151
rect 9689 19117 9723 19151
rect 9956 19117 9990 19151
rect 11897 19117 11931 19151
rect 14105 19117 14139 19151
rect 15301 19117 15335 19151
rect 15557 19117 15591 19151
rect 17785 19117 17819 19151
rect 18889 19117 18923 19151
rect 12164 19049 12198 19083
rect 11069 18981 11103 19015
rect 14289 18981 14323 19015
rect 16681 18981 16715 19015
rect 7021 18777 7055 18811
rect 7389 18777 7423 18811
rect 7481 18777 7515 18811
rect 9045 18777 9079 18811
rect 10149 18777 10183 18811
rect 10517 18777 10551 18811
rect 12449 18777 12483 18811
rect 18061 18777 18095 18811
rect 18521 18777 18555 18811
rect 20177 18709 20211 18743
rect 8953 18641 8987 18675
rect 12817 18641 12851 18675
rect 14657 18641 14691 18675
rect 16017 18641 16051 18675
rect 18429 18641 18463 18675
rect 19901 18641 19935 18675
rect 6929 18573 6963 18607
rect 7573 18573 7607 18607
rect 9229 18573 9263 18607
rect 10609 18573 10643 18607
rect 10793 18573 10827 18607
rect 12909 18573 12943 18607
rect 13001 18573 13035 18607
rect 15761 18573 15795 18607
rect 18613 18573 18647 18607
rect 8585 18505 8619 18539
rect 17141 18505 17175 18539
rect 6929 18437 6963 18471
rect 14841 18437 14875 18471
rect 6929 18233 6963 18267
rect 12081 18233 12115 18267
rect 16313 18233 16347 18267
rect 8309 18097 8343 18131
rect 9873 18097 9907 18131
rect 5549 18029 5583 18063
rect 5816 18029 5850 18063
rect 11897 18029 11931 18063
rect 13001 18029 13035 18063
rect 14105 18029 14139 18063
rect 16129 18029 16163 18063
rect 17233 18029 17267 18063
rect 19717 18029 19751 18063
rect 8125 17961 8159 17995
rect 17500 17961 17534 17995
rect 7757 17893 7791 17927
rect 8217 17893 8251 17927
rect 10885 17893 10919 17927
rect 13185 17893 13219 17927
rect 14289 17893 14323 17927
rect 18613 17893 18647 17927
rect 19901 17893 19935 17927
rect 6929 17689 6963 17723
rect 9689 17689 9723 17723
rect 11345 17689 11379 17723
rect 12909 17689 12943 17723
rect 15025 17689 15059 17723
rect 18613 17689 18647 17723
rect 7389 17621 7423 17655
rect 20177 17621 20211 17655
rect 7297 17553 7331 17587
rect 9597 17553 9631 17587
rect 12817 17553 12851 17587
rect 14933 17553 14967 17587
rect 16865 17553 16899 17587
rect 18521 17553 18555 17587
rect 19901 17553 19935 17587
rect 7481 17485 7515 17519
rect 9781 17485 9815 17519
rect 13001 17485 13035 17519
rect 15117 17485 15151 17519
rect 18705 17485 18739 17519
rect 18153 17417 18187 17451
rect 9229 17349 9263 17383
rect 12449 17349 12483 17383
rect 14565 17349 14599 17383
rect 17049 17349 17083 17383
rect 7665 17145 7699 17179
rect 14381 17145 14415 17179
rect 11897 17077 11931 17111
rect 19717 17009 19751 17043
rect 6285 16941 6319 16975
rect 6552 16941 6586 16975
rect 10517 16941 10551 16975
rect 12909 16941 12943 16975
rect 13001 16941 13035 16975
rect 15301 16941 15335 16975
rect 15557 16941 15591 16975
rect 18429 16941 18463 16975
rect 19533 16941 19567 16975
rect 10762 16873 10796 16907
rect 13268 16873 13302 16907
rect 12725 16805 12759 16839
rect 16681 16805 16715 16839
rect 18613 16805 18647 16839
rect 7389 16601 7423 16635
rect 10517 16601 10551 16635
rect 13829 16601 13863 16635
rect 14841 16601 14875 16635
rect 9404 16533 9438 16567
rect 16028 16533 16062 16567
rect 18521 16533 18555 16567
rect 20177 16533 20211 16567
rect 9045 16465 9079 16499
rect 12449 16465 12483 16499
rect 12716 16465 12750 16499
rect 14657 16465 14691 16499
rect 18429 16465 18463 16499
rect 19901 16465 19935 16499
rect 9137 16397 9171 16431
rect 11345 16397 11379 16431
rect 15761 16397 15795 16431
rect 18613 16397 18647 16431
rect 17141 16329 17175 16363
rect 8861 16261 8895 16295
rect 18061 16261 18095 16295
rect 7113 16057 7147 16091
rect 15577 16057 15611 16091
rect 10149 15989 10183 16023
rect 12817 15989 12851 16023
rect 10701 15921 10735 15955
rect 13277 15921 13311 15955
rect 13461 15921 13495 15955
rect 16129 15921 16163 15955
rect 5733 15853 5767 15887
rect 10517 15853 10551 15887
rect 13185 15853 13219 15887
rect 17325 15853 17359 15887
rect 17592 15853 17626 15887
rect 19533 15853 19567 15887
rect 6000 15785 6034 15819
rect 16037 15785 16071 15819
rect 19809 15785 19843 15819
rect 10609 15717 10643 15751
rect 15945 15717 15979 15751
rect 18705 15717 18739 15751
rect 7297 15513 7331 15547
rect 9781 15513 9815 15547
rect 11621 15513 11655 15547
rect 15853 15513 15887 15547
rect 17049 15513 17083 15547
rect 18705 15513 18739 15547
rect 7205 15445 7239 15479
rect 8668 15377 8702 15411
rect 11805 15377 11839 15411
rect 14289 15377 14323 15411
rect 16865 15377 16899 15411
rect 18613 15377 18647 15411
rect 19993 15377 20027 15411
rect 7481 15309 7515 15343
rect 8401 15309 8435 15343
rect 10609 15309 10643 15343
rect 14381 15309 14415 15343
rect 14565 15309 14599 15343
rect 18797 15309 18831 15343
rect 20177 15309 20211 15343
rect 18245 15241 18279 15275
rect 6837 15173 6871 15207
rect 13921 15173 13955 15207
rect 11253 14969 11287 15003
rect 17509 14969 17543 15003
rect 8769 14901 8803 14935
rect 9689 14901 9723 14935
rect 10241 14833 10275 14867
rect 11713 14833 11747 14867
rect 11897 14833 11931 14867
rect 12817 14833 12851 14867
rect 15853 14833 15887 14867
rect 19717 14833 19751 14867
rect 7389 14765 7423 14799
rect 10057 14765 10091 14799
rect 13084 14765 13118 14799
rect 17325 14765 17359 14799
rect 18429 14765 18463 14799
rect 19543 14765 19577 14799
rect 7656 14697 7690 14731
rect 10149 14629 10183 14663
rect 11621 14629 11655 14663
rect 14197 14629 14231 14663
rect 15301 14629 15335 14663
rect 15669 14629 15703 14663
rect 15761 14629 15795 14663
rect 18613 14629 18647 14663
rect 8217 14425 8251 14459
rect 13829 14425 13863 14459
rect 14749 14425 14783 14459
rect 17141 14425 17175 14459
rect 19441 14425 19475 14459
rect 10232 14357 10266 14391
rect 6837 14289 6871 14323
rect 7104 14289 7138 14323
rect 9965 14289 9999 14323
rect 12716 14289 12750 14323
rect 16028 14289 16062 14323
rect 18328 14289 18362 14323
rect 20545 14289 20579 14323
rect 12449 14221 12483 14255
rect 15761 14221 15795 14255
rect 18061 14221 18095 14255
rect 11345 14085 11379 14119
rect 20729 14085 20763 14119
rect 13093 13881 13127 13915
rect 17325 13881 17359 13915
rect 6929 13813 6963 13847
rect 10241 13813 10275 13847
rect 13645 13813 13679 13847
rect 7481 13745 7515 13779
rect 10701 13745 10735 13779
rect 10885 13745 10919 13779
rect 14105 13745 14139 13779
rect 14197 13745 14231 13779
rect 16129 13745 16163 13779
rect 18889 13745 18923 13779
rect 7297 13677 7331 13711
rect 11805 13677 11839 13711
rect 15853 13677 15887 13711
rect 17141 13677 17175 13711
rect 18705 13677 18739 13711
rect 14013 13609 14047 13643
rect 19809 13609 19843 13643
rect 7389 13541 7423 13575
rect 10609 13541 10643 13575
rect 18245 13541 18279 13575
rect 18613 13541 18647 13575
rect 7021 13337 7055 13371
rect 12909 13337 12943 13371
rect 16313 13337 16347 13371
rect 19073 13337 19107 13371
rect 7481 13269 7515 13303
rect 10416 13269 10450 13303
rect 14657 13269 14691 13303
rect 20453 13269 20487 13303
rect 7389 13201 7423 13235
rect 8861 13201 8895 13235
rect 12817 13201 12851 13235
rect 14381 13201 14415 13235
rect 16129 13201 16163 13235
rect 16681 13201 16715 13235
rect 18981 13201 19015 13235
rect 20177 13201 20211 13235
rect 7665 13133 7699 13167
rect 9137 13133 9171 13167
rect 10149 13133 10183 13167
rect 13093 13133 13127 13167
rect 16773 13133 16807 13167
rect 16957 13133 16991 13167
rect 19165 13133 19199 13167
rect 11529 13065 11563 13099
rect 12449 12997 12483 13031
rect 18613 12997 18647 13031
rect 7389 12793 7423 12827
rect 18889 12793 18923 12827
rect 15761 12725 15795 12759
rect 18061 12725 18095 12759
rect 14013 12657 14047 12691
rect 19349 12657 19383 12691
rect 19441 12657 19475 12691
rect 6009 12589 6043 12623
rect 6276 12589 6310 12623
rect 11253 12589 11287 12623
rect 11520 12589 11554 12623
rect 13921 12589 13955 12623
rect 15577 12589 15611 12623
rect 16681 12589 16715 12623
rect 19257 12589 19291 12623
rect 16948 12521 16982 12555
rect 12633 12453 12667 12487
rect 13461 12453 13495 12487
rect 13829 12453 13863 12487
rect 7297 12249 7331 12283
rect 10057 12249 10091 12283
rect 13093 12249 13127 12283
rect 16865 12249 16899 12283
rect 18521 12249 18555 12283
rect 19625 12249 19659 12283
rect 20729 12249 20763 12283
rect 8944 12181 8978 12215
rect 13001 12181 13035 12215
rect 8677 12113 8711 12147
rect 14381 12113 14415 12147
rect 15752 12113 15786 12147
rect 18337 12113 18371 12147
rect 19441 12113 19475 12147
rect 20545 12113 20579 12147
rect 13277 12045 13311 12079
rect 15485 12045 15519 12079
rect 12633 11909 12667 11943
rect 14565 11909 14599 11943
rect 15301 11637 15335 11671
rect 13645 11569 13679 11603
rect 15853 11569 15887 11603
rect 16865 11569 16899 11603
rect 18153 11569 18187 11603
rect 19717 11569 19751 11603
rect 12541 11501 12575 11535
rect 17877 11501 17911 11535
rect 19533 11501 19567 11535
rect 15761 11433 15795 11467
rect 12357 11365 12391 11399
rect 15669 11365 15703 11399
rect 13001 11161 13035 11195
rect 15761 11161 15795 11195
rect 17049 11161 17083 11195
rect 18061 11161 18095 11195
rect 20545 11161 20579 11195
rect 12909 11025 12943 11059
rect 14289 11025 14323 11059
rect 14637 11025 14671 11059
rect 16865 11025 16899 11059
rect 18429 11025 18463 11059
rect 20361 11025 20395 11059
rect 13185 10957 13219 10991
rect 14381 10957 14415 10991
rect 18521 10957 18555 10991
rect 18705 10957 18739 10991
rect 12541 10889 12575 10923
rect 14105 10821 14139 10855
rect 13277 10617 13311 10651
rect 15301 10617 15335 10651
rect 19901 10617 19935 10651
rect 15761 10481 15795 10515
rect 15853 10481 15887 10515
rect 10609 10413 10643 10447
rect 11897 10413 11931 10447
rect 17325 10413 17359 10447
rect 19717 10413 19751 10447
rect 12164 10345 12198 10379
rect 17592 10345 17626 10379
rect 10425 10277 10459 10311
rect 14197 10277 14231 10311
rect 15669 10277 15703 10311
rect 18705 10277 18739 10311
rect 15669 10073 15703 10107
rect 18061 10073 18095 10107
rect 20729 10073 20763 10107
rect 13246 10005 13280 10039
rect 18429 9937 18463 9971
rect 20545 9937 20579 9971
rect 13001 9869 13035 9903
rect 15761 9869 15795 9903
rect 15853 9869 15887 9903
rect 18521 9869 18555 9903
rect 18613 9869 18647 9903
rect 14381 9801 14415 9835
rect 15301 9801 15335 9835
rect 17969 9529 18003 9563
rect 11713 9461 11747 9495
rect 13277 9461 13311 9495
rect 19901 9461 19935 9495
rect 11529 9325 11563 9359
rect 13093 9325 13127 9359
rect 15301 9325 15335 9359
rect 16589 9325 16623 9359
rect 19717 9325 19751 9359
rect 15577 9257 15611 9291
rect 16834 9257 16868 9291
rect 14933 8985 14967 9019
rect 15945 8985 15979 9019
rect 18061 8985 18095 9019
rect 19625 8985 19659 9019
rect 20729 8985 20763 9019
rect 11345 8917 11379 8951
rect 13369 8917 13403 8951
rect 11069 8849 11103 8883
rect 13093 8849 13127 8883
rect 14749 8849 14783 8883
rect 16313 8849 16347 8883
rect 19441 8849 19475 8883
rect 20545 8849 20579 8883
rect 16405 8781 16439 8815
rect 16589 8781 16623 8815
rect 13553 8441 13587 8475
rect 16957 8441 16991 8475
rect 11345 8305 11379 8339
rect 14197 8305 14231 8339
rect 10333 8237 10367 8271
rect 15577 8237 15611 8271
rect 11590 8169 11624 8203
rect 14013 8169 14047 8203
rect 15822 8169 15856 8203
rect 12725 8101 12759 8135
rect 13921 8101 13955 8135
rect 11161 7897 11195 7931
rect 13277 7897 13311 7931
rect 16497 7897 16531 7931
rect 20729 7897 20763 7931
rect 14534 7829 14568 7863
rect 10048 7761 10082 7795
rect 19441 7761 19475 7795
rect 20545 7761 20579 7795
rect 9781 7693 9815 7727
rect 14289 7693 14323 7727
rect 19625 7625 19659 7659
rect 15669 7557 15703 7591
rect 10793 7353 10827 7387
rect 14197 7353 14231 7387
rect 16497 7353 16531 7387
rect 11345 7217 11379 7251
rect 12817 7217 12851 7251
rect 17049 7217 17083 7251
rect 13073 7149 13107 7183
rect 16957 7149 16991 7183
rect 11161 7081 11195 7115
rect 16865 7081 16899 7115
rect 11253 7013 11287 7047
rect 11161 6741 11195 6775
rect 14013 6741 14047 6775
rect 8197 6673 8231 6707
rect 11253 6673 11287 6707
rect 14105 6673 14139 6707
rect 19441 6673 19475 6707
rect 20545 6673 20579 6707
rect 7941 6605 7975 6639
rect 11345 6605 11379 6639
rect 14197 6605 14231 6639
rect 9321 6537 9355 6571
rect 10793 6537 10827 6571
rect 13645 6537 13679 6571
rect 19625 6537 19659 6571
rect 20729 6469 20763 6503
rect 20729 5721 20763 5755
rect 20545 5585 20579 5619
rect 13185 4633 13219 4667
rect 13001 4497 13035 4531
rect 20729 3545 20763 3579
rect 20545 3409 20579 3443
<< metal1 >>
rect 1104 20554 21896 20576
rect 1104 20502 4447 20554
rect 4499 20502 4511 20554
rect 4563 20502 4575 20554
rect 4627 20502 4639 20554
rect 4691 20502 11378 20554
rect 11430 20502 11442 20554
rect 11494 20502 11506 20554
rect 11558 20502 11570 20554
rect 11622 20502 18308 20554
rect 18360 20502 18372 20554
rect 18424 20502 18436 20554
rect 18488 20502 18500 20554
rect 18552 20502 21896 20554
rect 1104 20480 21896 20502
rect 11609 20443 11667 20449
rect 11609 20409 11621 20443
rect 11655 20440 11667 20443
rect 17862 20440 17868 20452
rect 11655 20412 17868 20440
rect 11655 20409 11667 20412
rect 11609 20403 11667 20409
rect 17862 20400 17868 20412
rect 17920 20400 17926 20452
rect 12989 20375 13047 20381
rect 12989 20341 13001 20375
rect 13035 20372 13047 20375
rect 13035 20344 18368 20372
rect 13035 20341 13047 20344
rect 12989 20335 13047 20341
rect 7837 20307 7895 20313
rect 7837 20273 7849 20307
rect 7883 20304 7895 20307
rect 8202 20304 8208 20316
rect 7883 20276 8208 20304
rect 7883 20273 7895 20276
rect 7837 20267 7895 20273
rect 8202 20264 8208 20276
rect 8260 20264 8266 20316
rect 10413 20307 10471 20313
rect 10413 20273 10425 20307
rect 10459 20304 10471 20307
rect 10459 20276 13216 20304
rect 10459 20273 10471 20276
rect 10413 20267 10471 20273
rect 5810 20196 5816 20248
rect 5868 20236 5874 20248
rect 11422 20236 11428 20248
rect 5868 20208 9168 20236
rect 11383 20208 11428 20236
rect 5868 20196 5874 20208
rect 7098 20128 7104 20180
rect 7156 20168 7162 20180
rect 7653 20171 7711 20177
rect 7653 20168 7665 20171
rect 7156 20140 7665 20168
rect 7156 20128 7162 20140
rect 7653 20137 7665 20140
rect 7699 20137 7711 20171
rect 9140 20168 9168 20208
rect 11422 20196 11428 20208
rect 11480 20196 11486 20248
rect 13078 20236 13084 20248
rect 12820 20208 13084 20236
rect 12820 20168 12848 20208
rect 13078 20196 13084 20208
rect 13136 20196 13142 20248
rect 13188 20236 13216 20276
rect 13262 20264 13268 20316
rect 13320 20304 13326 20316
rect 13541 20307 13599 20313
rect 13541 20304 13553 20307
rect 13320 20276 13553 20304
rect 13320 20264 13326 20276
rect 13541 20273 13553 20276
rect 13587 20273 13599 20307
rect 13541 20267 13599 20273
rect 16114 20264 16120 20316
rect 16172 20304 16178 20316
rect 16577 20307 16635 20313
rect 16577 20304 16589 20307
rect 16172 20276 16589 20304
rect 16172 20264 16178 20276
rect 16577 20273 16589 20276
rect 16623 20273 16635 20307
rect 16577 20267 16635 20273
rect 13188 20208 13400 20236
rect 13372 20168 13400 20208
rect 13446 20196 13452 20248
rect 13504 20236 13510 20248
rect 18340 20245 18368 20344
rect 18325 20239 18383 20245
rect 13504 20208 16528 20236
rect 13504 20196 13510 20208
rect 16393 20171 16451 20177
rect 16393 20168 16405 20171
rect 9140 20140 12848 20168
rect 12912 20140 13308 20168
rect 13372 20140 16405 20168
rect 7653 20131 7711 20137
rect 7190 20100 7196 20112
rect 7151 20072 7196 20100
rect 7190 20060 7196 20072
rect 7248 20060 7254 20112
rect 7282 20060 7288 20112
rect 7340 20100 7346 20112
rect 7561 20103 7619 20109
rect 7561 20100 7573 20103
rect 7340 20072 7573 20100
rect 7340 20060 7346 20072
rect 7561 20069 7573 20072
rect 7607 20069 7619 20103
rect 7561 20063 7619 20069
rect 11146 20060 11152 20112
rect 11204 20100 11210 20112
rect 12912 20100 12940 20140
rect 11204 20072 12940 20100
rect 13280 20100 13308 20140
rect 16393 20137 16405 20140
rect 16439 20137 16451 20171
rect 16500 20168 16528 20208
rect 18325 20205 18337 20239
rect 18371 20205 18383 20239
rect 19981 20239 20039 20245
rect 19981 20236 19993 20239
rect 18325 20199 18383 20205
rect 18432 20208 19993 20236
rect 18432 20168 18460 20208
rect 19981 20205 19993 20208
rect 20027 20205 20039 20239
rect 19981 20199 20039 20205
rect 16500 20140 18460 20168
rect 18601 20171 18659 20177
rect 16393 20131 16451 20137
rect 18601 20137 18613 20171
rect 18647 20168 18659 20171
rect 18690 20168 18696 20180
rect 18647 20140 18696 20168
rect 18647 20137 18659 20140
rect 18601 20131 18659 20137
rect 18690 20128 18696 20140
rect 18748 20128 18754 20180
rect 13357 20103 13415 20109
rect 13357 20100 13369 20103
rect 13280 20072 13369 20100
rect 11204 20060 11210 20072
rect 13357 20069 13369 20072
rect 13403 20069 13415 20103
rect 13357 20063 13415 20069
rect 13449 20103 13507 20109
rect 13449 20069 13461 20103
rect 13495 20100 13507 20103
rect 13630 20100 13636 20112
rect 13495 20072 13636 20100
rect 13495 20069 13507 20072
rect 13449 20063 13507 20069
rect 13630 20060 13636 20072
rect 13688 20060 13694 20112
rect 16025 20103 16083 20109
rect 16025 20069 16037 20103
rect 16071 20100 16083 20103
rect 16298 20100 16304 20112
rect 16071 20072 16304 20100
rect 16071 20069 16083 20072
rect 16025 20063 16083 20069
rect 16298 20060 16304 20072
rect 16356 20060 16362 20112
rect 16482 20060 16488 20112
rect 16540 20100 16546 20112
rect 16540 20072 16585 20100
rect 16540 20060 16546 20072
rect 19242 20060 19248 20112
rect 19300 20100 19306 20112
rect 20165 20103 20223 20109
rect 20165 20100 20177 20103
rect 19300 20072 20177 20100
rect 19300 20060 19306 20072
rect 20165 20069 20177 20072
rect 20211 20069 20223 20103
rect 20165 20063 20223 20069
rect 1104 20010 21896 20032
rect 1104 19958 7912 20010
rect 7964 19958 7976 20010
rect 8028 19958 8040 20010
rect 8092 19958 8104 20010
rect 8156 19958 14843 20010
rect 14895 19958 14907 20010
rect 14959 19958 14971 20010
rect 15023 19958 15035 20010
rect 15087 19958 21896 20010
rect 1104 19936 21896 19958
rect 9214 19856 9220 19908
rect 9272 19896 9278 19908
rect 15194 19896 15200 19908
rect 9272 19868 15200 19896
rect 9272 19856 9278 19868
rect 15194 19856 15200 19868
rect 15252 19856 15258 19908
rect 16022 19896 16028 19908
rect 15983 19868 16028 19896
rect 16022 19856 16028 19868
rect 16080 19856 16086 19908
rect 16390 19856 16396 19908
rect 16448 19896 16454 19908
rect 19426 19896 19432 19908
rect 16448 19868 19432 19896
rect 16448 19856 16454 19868
rect 19426 19856 19432 19868
rect 19484 19856 19490 19908
rect 7190 19788 7196 19840
rect 7248 19828 7254 19840
rect 12342 19828 12348 19840
rect 7248 19800 12348 19828
rect 7248 19788 7254 19800
rect 12342 19788 12348 19800
rect 12400 19788 12406 19840
rect 15102 19788 15108 19840
rect 15160 19828 15166 19840
rect 15160 19800 16068 19828
rect 15160 19788 15166 19800
rect 7092 19763 7150 19769
rect 7092 19729 7104 19763
rect 7138 19760 7150 19763
rect 7466 19760 7472 19772
rect 7138 19732 7472 19760
rect 7138 19729 7150 19732
rect 7092 19723 7150 19729
rect 7466 19720 7472 19732
rect 7524 19720 7530 19772
rect 8754 19720 8760 19772
rect 8812 19760 8818 19772
rect 9214 19760 9220 19772
rect 8812 19732 9220 19760
rect 8812 19720 8818 19732
rect 9214 19720 9220 19732
rect 9272 19760 9278 19772
rect 9381 19763 9439 19769
rect 9381 19760 9393 19763
rect 9272 19732 9393 19760
rect 9272 19720 9278 19732
rect 9381 19729 9393 19732
rect 9427 19729 9439 19763
rect 9381 19723 9439 19729
rect 12986 19720 12992 19772
rect 13044 19760 13050 19772
rect 13262 19760 13268 19772
rect 13044 19732 13268 19760
rect 13044 19720 13050 19732
rect 13262 19720 13268 19732
rect 13320 19760 13326 19772
rect 13613 19763 13671 19769
rect 13613 19760 13625 19763
rect 13320 19732 13625 19760
rect 13320 19720 13326 19732
rect 13613 19729 13625 19732
rect 13659 19729 13671 19763
rect 13613 19723 13671 19729
rect 15838 19720 15844 19772
rect 15896 19760 15902 19772
rect 15933 19763 15991 19769
rect 15933 19760 15945 19763
rect 15896 19732 15945 19760
rect 15896 19720 15902 19732
rect 15933 19729 15945 19732
rect 15979 19729 15991 19763
rect 16040 19760 16068 19800
rect 16224 19800 19840 19828
rect 16224 19760 16252 19800
rect 16040 19732 16252 19760
rect 15933 19723 15991 19729
rect 16298 19720 16304 19772
rect 16356 19760 16362 19772
rect 19812 19769 19840 19800
rect 18049 19763 18107 19769
rect 18049 19760 18061 19763
rect 16356 19732 18061 19760
rect 16356 19720 16362 19732
rect 18049 19729 18061 19732
rect 18095 19729 18107 19763
rect 18049 19723 18107 19729
rect 19797 19763 19855 19769
rect 19797 19729 19809 19763
rect 19843 19729 19855 19763
rect 19797 19723 19855 19729
rect 6822 19692 6828 19704
rect 6783 19664 6828 19692
rect 6822 19652 6828 19664
rect 6880 19652 6886 19704
rect 9122 19692 9128 19704
rect 9083 19664 9128 19692
rect 9122 19652 9128 19664
rect 9180 19652 9186 19704
rect 11054 19652 11060 19704
rect 11112 19692 11118 19704
rect 11333 19695 11391 19701
rect 11333 19692 11345 19695
rect 11112 19664 11345 19692
rect 11112 19652 11118 19664
rect 11333 19661 11345 19664
rect 11379 19661 11391 19695
rect 11333 19655 11391 19661
rect 12526 19652 12532 19704
rect 12584 19692 12590 19704
rect 13357 19695 13415 19701
rect 13357 19692 13369 19695
rect 12584 19664 13369 19692
rect 12584 19652 12590 19664
rect 13357 19661 13369 19664
rect 13403 19661 13415 19695
rect 13357 19655 13415 19661
rect 15654 19652 15660 19704
rect 15712 19692 15718 19704
rect 16117 19695 16175 19701
rect 16117 19692 16129 19695
rect 15712 19664 16129 19692
rect 15712 19652 15718 19664
rect 16117 19661 16129 19664
rect 16163 19661 16175 19695
rect 16117 19655 16175 19661
rect 16390 19652 16396 19704
rect 16448 19692 16454 19704
rect 18233 19695 18291 19701
rect 18233 19692 18245 19695
rect 16448 19664 18245 19692
rect 16448 19652 16454 19664
rect 18233 19661 18245 19664
rect 18279 19661 18291 19695
rect 19978 19692 19984 19704
rect 19939 19664 19984 19692
rect 18233 19655 18291 19661
rect 19978 19652 19984 19664
rect 20036 19652 20042 19704
rect 15565 19627 15623 19633
rect 15565 19593 15577 19627
rect 15611 19624 15623 19627
rect 16482 19624 16488 19636
rect 15611 19596 16488 19624
rect 15611 19593 15623 19596
rect 15565 19587 15623 19593
rect 16482 19584 16488 19596
rect 16540 19584 16546 19636
rect 8202 19556 8208 19568
rect 8163 19528 8208 19556
rect 8202 19516 8208 19528
rect 8260 19516 8266 19568
rect 10502 19556 10508 19568
rect 10463 19528 10508 19556
rect 10502 19516 10508 19528
rect 10560 19516 10566 19568
rect 14737 19559 14795 19565
rect 14737 19525 14749 19559
rect 14783 19556 14795 19559
rect 15378 19556 15384 19568
rect 14783 19528 15384 19556
rect 14783 19525 14795 19528
rect 14737 19519 14795 19525
rect 15378 19516 15384 19528
rect 15436 19516 15442 19568
rect 1104 19466 21896 19488
rect 1104 19414 4447 19466
rect 4499 19414 4511 19466
rect 4563 19414 4575 19466
rect 4627 19414 4639 19466
rect 4691 19414 11378 19466
rect 11430 19414 11442 19466
rect 11494 19414 11506 19466
rect 11558 19414 11570 19466
rect 11622 19414 18308 19466
rect 18360 19414 18372 19466
rect 18424 19414 18436 19466
rect 18488 19414 18500 19466
rect 18552 19414 21896 19466
rect 1104 19392 21896 19414
rect 8754 19352 8760 19364
rect 8715 19324 8760 19352
rect 8754 19312 8760 19324
rect 8812 19312 8818 19364
rect 12526 19352 12532 19364
rect 11900 19324 12532 19352
rect 6270 19176 6276 19228
rect 6328 19216 6334 19228
rect 6822 19216 6828 19228
rect 6328 19188 6828 19216
rect 6328 19176 6334 19188
rect 6822 19176 6828 19188
rect 6880 19216 6886 19228
rect 6880 19188 7420 19216
rect 6880 19176 6886 19188
rect 6365 19151 6423 19157
rect 6365 19117 6377 19151
rect 6411 19148 6423 19151
rect 7282 19148 7288 19160
rect 6411 19120 7288 19148
rect 6411 19117 6423 19120
rect 6365 19111 6423 19117
rect 7282 19108 7288 19120
rect 7340 19108 7346 19160
rect 7392 19157 7420 19188
rect 7377 19151 7435 19157
rect 7377 19117 7389 19151
rect 7423 19117 7435 19151
rect 7377 19111 7435 19117
rect 7644 19151 7702 19157
rect 7644 19117 7656 19151
rect 7690 19148 7702 19151
rect 8202 19148 8208 19160
rect 7690 19120 8208 19148
rect 7690 19117 7702 19120
rect 7644 19111 7702 19117
rect 8202 19108 8208 19120
rect 8260 19108 8266 19160
rect 9122 19108 9128 19160
rect 9180 19148 9186 19160
rect 9677 19151 9735 19157
rect 9677 19148 9689 19151
rect 9180 19120 9689 19148
rect 9180 19108 9186 19120
rect 9677 19117 9689 19120
rect 9723 19117 9735 19151
rect 9677 19111 9735 19117
rect 9944 19151 10002 19157
rect 9944 19117 9956 19151
rect 9990 19148 10002 19151
rect 10502 19148 10508 19160
rect 9990 19120 10508 19148
rect 9990 19117 10002 19120
rect 9944 19111 10002 19117
rect 10502 19108 10508 19120
rect 10560 19148 10566 19160
rect 10778 19148 10784 19160
rect 10560 19120 10784 19148
rect 10560 19108 10566 19120
rect 10778 19108 10784 19120
rect 10836 19108 10842 19160
rect 11900 19157 11928 19324
rect 12526 19312 12532 19324
rect 12584 19312 12590 19364
rect 13262 19352 13268 19364
rect 13223 19324 13268 19352
rect 13262 19312 13268 19324
rect 13320 19312 13326 19364
rect 13906 19312 13912 19364
rect 13964 19352 13970 19364
rect 16390 19352 16396 19364
rect 13964 19324 16396 19352
rect 13964 19312 13970 19324
rect 16390 19312 16396 19324
rect 16448 19312 16454 19364
rect 12894 19244 12900 19296
rect 12952 19284 12958 19296
rect 13630 19284 13636 19296
rect 12952 19256 13636 19284
rect 12952 19244 12958 19256
rect 13630 19244 13636 19256
rect 13688 19244 13694 19296
rect 17954 19284 17960 19296
rect 17915 19256 17960 19284
rect 17954 19244 17960 19256
rect 18012 19244 18018 19296
rect 14016 19188 14228 19216
rect 11885 19151 11943 19157
rect 11885 19117 11897 19151
rect 11931 19117 11943 19151
rect 14016 19148 14044 19188
rect 11885 19111 11943 19117
rect 11992 19120 14044 19148
rect 14093 19151 14151 19157
rect 1394 19040 1400 19092
rect 1452 19080 1458 19092
rect 1452 19052 2820 19080
rect 1452 19040 1458 19052
rect 2792 19012 2820 19052
rect 3602 19040 3608 19092
rect 3660 19080 3666 19092
rect 9490 19080 9496 19092
rect 3660 19052 9496 19080
rect 3660 19040 3666 19052
rect 9490 19040 9496 19052
rect 9548 19040 9554 19092
rect 10134 19040 10140 19092
rect 10192 19080 10198 19092
rect 11992 19080 12020 19120
rect 14093 19117 14105 19151
rect 14139 19117 14151 19151
rect 14200 19148 14228 19188
rect 15102 19176 15108 19228
rect 15160 19176 15166 19228
rect 17494 19176 17500 19228
rect 17552 19216 17558 19228
rect 17552 19188 17724 19216
rect 17552 19176 17558 19188
rect 15120 19148 15148 19176
rect 15286 19148 15292 19160
rect 14200 19120 15148 19148
rect 15247 19120 15292 19148
rect 14093 19111 14151 19117
rect 10192 19052 12020 19080
rect 12152 19083 12210 19089
rect 10192 19040 10198 19052
rect 12152 19049 12164 19083
rect 12198 19080 12210 19083
rect 12986 19080 12992 19092
rect 12198 19052 12992 19080
rect 12198 19049 12210 19052
rect 12152 19043 12210 19049
rect 8294 19012 8300 19024
rect 2792 18984 8300 19012
rect 8294 18972 8300 18984
rect 8352 18972 8358 19024
rect 8662 18972 8668 19024
rect 8720 19012 8726 19024
rect 10962 19012 10968 19024
rect 8720 18984 10968 19012
rect 8720 18972 8726 18984
rect 10962 18972 10968 18984
rect 11020 18972 11026 19024
rect 11057 19015 11115 19021
rect 11057 18981 11069 19015
rect 11103 19012 11115 19015
rect 12268 19012 12296 19052
rect 12986 19040 12992 19052
rect 13044 19040 13050 19092
rect 14108 19080 14136 19111
rect 15286 19108 15292 19120
rect 15344 19108 15350 19160
rect 15378 19108 15384 19160
rect 15436 19148 15442 19160
rect 15562 19157 15568 19160
rect 15545 19151 15568 19157
rect 15545 19148 15557 19151
rect 15436 19120 15557 19148
rect 15436 19108 15442 19120
rect 15545 19117 15557 19120
rect 15620 19148 15626 19160
rect 17696 19148 17724 19188
rect 18046 19176 18052 19228
rect 18104 19216 18110 19228
rect 19061 19219 19119 19225
rect 19061 19216 19073 19219
rect 18104 19188 19073 19216
rect 18104 19176 18110 19188
rect 19061 19185 19073 19188
rect 19107 19185 19119 19219
rect 19061 19179 19119 19185
rect 17773 19151 17831 19157
rect 17773 19148 17785 19151
rect 15620 19120 15693 19148
rect 17696 19120 17785 19148
rect 15545 19111 15568 19117
rect 15562 19108 15568 19111
rect 15620 19108 15626 19120
rect 17773 19117 17785 19120
rect 17819 19117 17831 19151
rect 17773 19111 17831 19117
rect 18138 19108 18144 19160
rect 18196 19148 18202 19160
rect 18877 19151 18935 19157
rect 18877 19148 18889 19151
rect 18196 19120 18889 19148
rect 18196 19108 18202 19120
rect 18877 19117 18889 19120
rect 18923 19117 18935 19151
rect 18877 19111 18935 19117
rect 15194 19080 15200 19092
rect 14108 19052 15200 19080
rect 15194 19040 15200 19052
rect 15252 19040 15258 19092
rect 16758 19040 16764 19092
rect 16816 19080 16822 19092
rect 19978 19080 19984 19092
rect 16816 19052 19984 19080
rect 16816 19040 16822 19052
rect 19978 19040 19984 19052
rect 20036 19040 20042 19092
rect 11103 18984 12296 19012
rect 11103 18981 11115 18984
rect 11057 18975 11115 18981
rect 12342 18972 12348 19024
rect 12400 19012 12406 19024
rect 12802 19012 12808 19024
rect 12400 18984 12808 19012
rect 12400 18972 12406 18984
rect 12802 18972 12808 18984
rect 12860 18972 12866 19024
rect 14277 19015 14335 19021
rect 14277 18981 14289 19015
rect 14323 19012 14335 19015
rect 14366 19012 14372 19024
rect 14323 18984 14372 19012
rect 14323 18981 14335 18984
rect 14277 18975 14335 18981
rect 14366 18972 14372 18984
rect 14424 18972 14430 19024
rect 16114 18972 16120 19024
rect 16172 19012 16178 19024
rect 16669 19015 16727 19021
rect 16669 19012 16681 19015
rect 16172 18984 16681 19012
rect 16172 18972 16178 18984
rect 16669 18981 16681 18984
rect 16715 18981 16727 19015
rect 16669 18975 16727 18981
rect 17034 18972 17040 19024
rect 17092 19012 17098 19024
rect 21082 19012 21088 19024
rect 17092 18984 21088 19012
rect 17092 18972 17098 18984
rect 21082 18972 21088 18984
rect 21140 18972 21146 19024
rect 1104 18922 21896 18944
rect 1104 18870 7912 18922
rect 7964 18870 7976 18922
rect 8028 18870 8040 18922
rect 8092 18870 8104 18922
rect 8156 18870 14843 18922
rect 14895 18870 14907 18922
rect 14959 18870 14971 18922
rect 15023 18870 15035 18922
rect 15087 18870 21896 18922
rect 1104 18848 21896 18870
rect 2498 18768 2504 18820
rect 2556 18808 2562 18820
rect 5534 18808 5540 18820
rect 2556 18780 5540 18808
rect 2556 18768 2562 18780
rect 5534 18768 5540 18780
rect 5592 18768 5598 18820
rect 7009 18811 7067 18817
rect 7009 18777 7021 18811
rect 7055 18808 7067 18811
rect 7098 18808 7104 18820
rect 7055 18780 7104 18808
rect 7055 18777 7067 18780
rect 7009 18771 7067 18777
rect 7098 18768 7104 18780
rect 7156 18768 7162 18820
rect 7374 18808 7380 18820
rect 7335 18780 7380 18808
rect 7374 18768 7380 18780
rect 7432 18768 7438 18820
rect 7469 18811 7527 18817
rect 7469 18777 7481 18811
rect 7515 18808 7527 18811
rect 7558 18808 7564 18820
rect 7515 18780 7564 18808
rect 7515 18777 7527 18780
rect 7469 18771 7527 18777
rect 7558 18768 7564 18780
rect 7616 18768 7622 18820
rect 7742 18768 7748 18820
rect 7800 18808 7806 18820
rect 9033 18811 9091 18817
rect 9033 18808 9045 18811
rect 7800 18780 9045 18808
rect 7800 18768 7806 18780
rect 9033 18777 9045 18780
rect 9079 18777 9091 18811
rect 10134 18808 10140 18820
rect 10095 18780 10140 18808
rect 9033 18771 9091 18777
rect 10134 18768 10140 18780
rect 10192 18768 10198 18820
rect 10505 18811 10563 18817
rect 10505 18777 10517 18811
rect 10551 18808 10563 18811
rect 11054 18808 11060 18820
rect 10551 18780 11060 18808
rect 10551 18777 10563 18780
rect 10505 18771 10563 18777
rect 11054 18768 11060 18780
rect 11112 18768 11118 18820
rect 11698 18768 11704 18820
rect 11756 18808 11762 18820
rect 12342 18808 12348 18820
rect 11756 18780 12348 18808
rect 11756 18768 11762 18780
rect 12342 18768 12348 18780
rect 12400 18768 12406 18820
rect 12437 18811 12495 18817
rect 12437 18777 12449 18811
rect 12483 18808 12495 18811
rect 12894 18808 12900 18820
rect 12483 18780 12900 18808
rect 12483 18777 12495 18780
rect 12437 18771 12495 18777
rect 12894 18768 12900 18780
rect 12952 18768 12958 18820
rect 14366 18768 14372 18820
rect 14424 18808 14430 18820
rect 17586 18808 17592 18820
rect 14424 18780 17592 18808
rect 14424 18768 14430 18780
rect 17586 18768 17592 18780
rect 17644 18768 17650 18820
rect 18046 18808 18052 18820
rect 18007 18780 18052 18808
rect 18046 18768 18052 18780
rect 18104 18768 18110 18820
rect 18506 18808 18512 18820
rect 18467 18780 18512 18808
rect 18506 18768 18512 18780
rect 18564 18768 18570 18820
rect 18598 18768 18604 18820
rect 18656 18808 18662 18820
rect 21358 18808 21364 18820
rect 18656 18780 21364 18808
rect 18656 18768 18662 18780
rect 21358 18768 21364 18780
rect 21416 18768 21422 18820
rect 4798 18700 4804 18752
rect 4856 18740 4862 18752
rect 8570 18740 8576 18752
rect 4856 18712 8576 18740
rect 4856 18700 4862 18712
rect 8570 18700 8576 18712
rect 8628 18700 8634 18752
rect 13078 18740 13084 18752
rect 8772 18712 13084 18740
rect 4154 18632 4160 18684
rect 4212 18672 4218 18684
rect 8772 18672 8800 18712
rect 13078 18700 13084 18712
rect 13136 18700 13142 18752
rect 20165 18743 20223 18749
rect 20165 18740 20177 18743
rect 14660 18712 20177 18740
rect 8938 18672 8944 18684
rect 4212 18644 8800 18672
rect 8899 18644 8944 18672
rect 4212 18632 4218 18644
rect 8938 18632 8944 18644
rect 8996 18632 9002 18684
rect 12805 18675 12863 18681
rect 12805 18641 12817 18675
rect 12851 18672 12863 18675
rect 13170 18672 13176 18684
rect 12851 18644 13176 18672
rect 12851 18641 12863 18644
rect 12805 18635 12863 18641
rect 13170 18632 13176 18644
rect 13228 18632 13234 18684
rect 14660 18681 14688 18712
rect 20165 18709 20177 18712
rect 20211 18709 20223 18743
rect 20165 18703 20223 18709
rect 16013 18681 16019 18684
rect 14645 18675 14703 18681
rect 14645 18641 14657 18675
rect 14691 18641 14703 18675
rect 14645 18635 14703 18641
rect 16005 18675 16019 18681
rect 16005 18641 16017 18675
rect 16071 18672 16077 18684
rect 16071 18644 16105 18672
rect 16005 18635 16019 18641
rect 16013 18632 16019 18635
rect 16071 18632 16077 18644
rect 17862 18632 17868 18684
rect 17920 18672 17926 18684
rect 18414 18672 18420 18684
rect 17920 18644 18276 18672
rect 18375 18644 18420 18672
rect 17920 18632 17926 18644
rect 842 18564 848 18616
rect 900 18604 906 18616
rect 6917 18607 6975 18613
rect 6917 18604 6929 18607
rect 900 18576 6929 18604
rect 900 18564 906 18576
rect 6917 18573 6929 18576
rect 6963 18573 6975 18607
rect 6917 18567 6975 18573
rect 7098 18564 7104 18616
rect 7156 18604 7162 18616
rect 7466 18604 7472 18616
rect 7156 18576 7472 18604
rect 7156 18564 7162 18576
rect 7466 18564 7472 18576
rect 7524 18604 7530 18616
rect 7561 18607 7619 18613
rect 7561 18604 7573 18607
rect 7524 18576 7573 18604
rect 7524 18564 7530 18576
rect 7561 18573 7573 18576
rect 7607 18573 7619 18607
rect 9214 18604 9220 18616
rect 9175 18576 9220 18604
rect 7561 18567 7619 18573
rect 9214 18564 9220 18576
rect 9272 18564 9278 18616
rect 10597 18607 10655 18613
rect 10597 18573 10609 18607
rect 10643 18573 10655 18607
rect 10597 18567 10655 18573
rect 290 18496 296 18548
rect 348 18536 354 18548
rect 8386 18536 8392 18548
rect 348 18508 8392 18536
rect 348 18496 354 18508
rect 8386 18496 8392 18508
rect 8444 18496 8450 18548
rect 8573 18539 8631 18545
rect 8573 18505 8585 18539
rect 8619 18536 8631 18539
rect 10612 18536 10640 18567
rect 10778 18564 10784 18616
rect 10836 18604 10842 18616
rect 10836 18576 10881 18604
rect 10836 18564 10842 18576
rect 11054 18564 11060 18616
rect 11112 18604 11118 18616
rect 12897 18607 12955 18613
rect 12897 18604 12909 18607
rect 11112 18576 12909 18604
rect 11112 18564 11118 18576
rect 12897 18573 12909 18576
rect 12943 18573 12955 18607
rect 12897 18567 12955 18573
rect 12986 18564 12992 18616
rect 13044 18604 13050 18616
rect 13044 18576 13089 18604
rect 13044 18564 13050 18576
rect 15286 18564 15292 18616
rect 15344 18604 15350 18616
rect 15749 18607 15807 18613
rect 15749 18604 15761 18607
rect 15344 18576 15761 18604
rect 15344 18564 15350 18576
rect 15749 18573 15761 18576
rect 15795 18573 15807 18607
rect 17494 18604 17500 18616
rect 15749 18567 15807 18573
rect 17144 18576 17500 18604
rect 17144 18545 17172 18576
rect 17494 18564 17500 18576
rect 17552 18604 17558 18616
rect 18248 18604 18276 18644
rect 18414 18632 18420 18644
rect 18472 18632 18478 18684
rect 18524 18644 19380 18672
rect 18524 18604 18552 18644
rect 17552 18576 18184 18604
rect 18248 18576 18552 18604
rect 18601 18607 18659 18613
rect 17552 18564 17558 18576
rect 8619 18508 10640 18536
rect 17129 18539 17187 18545
rect 8619 18505 8631 18508
rect 8573 18499 8631 18505
rect 17129 18505 17141 18539
rect 17175 18505 17187 18539
rect 18156 18536 18184 18576
rect 18601 18573 18613 18607
rect 18647 18573 18659 18607
rect 19352 18604 19380 18644
rect 19426 18632 19432 18684
rect 19484 18672 19490 18684
rect 19889 18675 19947 18681
rect 19889 18672 19901 18675
rect 19484 18644 19901 18672
rect 19484 18632 19490 18644
rect 19889 18641 19901 18644
rect 19935 18641 19947 18675
rect 19889 18635 19947 18641
rect 19794 18604 19800 18616
rect 19352 18576 19800 18604
rect 18601 18567 18659 18573
rect 18616 18536 18644 18567
rect 19794 18564 19800 18576
rect 19852 18564 19858 18616
rect 18156 18508 18644 18536
rect 17129 18499 17187 18505
rect 6917 18471 6975 18477
rect 6917 18437 6929 18471
rect 6963 18468 6975 18471
rect 11238 18468 11244 18480
rect 6963 18440 11244 18468
rect 6963 18437 6975 18440
rect 6917 18431 6975 18437
rect 11238 18428 11244 18440
rect 11296 18428 11302 18480
rect 12526 18428 12532 18480
rect 12584 18468 12590 18480
rect 14734 18468 14740 18480
rect 12584 18440 14740 18468
rect 12584 18428 12590 18440
rect 14734 18428 14740 18440
rect 14792 18428 14798 18480
rect 14829 18471 14887 18477
rect 14829 18437 14841 18471
rect 14875 18468 14887 18471
rect 17678 18468 17684 18480
rect 14875 18440 17684 18468
rect 14875 18437 14887 18440
rect 14829 18431 14887 18437
rect 17678 18428 17684 18440
rect 17736 18428 17742 18480
rect 17770 18428 17776 18480
rect 17828 18468 17834 18480
rect 20990 18468 20996 18480
rect 17828 18440 20996 18468
rect 17828 18428 17834 18440
rect 20990 18428 20996 18440
rect 21048 18428 21054 18480
rect 1104 18378 21896 18400
rect 1104 18326 4447 18378
rect 4499 18326 4511 18378
rect 4563 18326 4575 18378
rect 4627 18326 4639 18378
rect 4691 18326 11378 18378
rect 11430 18326 11442 18378
rect 11494 18326 11506 18378
rect 11558 18326 11570 18378
rect 11622 18326 18308 18378
rect 18360 18326 18372 18378
rect 18424 18326 18436 18378
rect 18488 18326 18500 18378
rect 18552 18326 21896 18378
rect 1104 18304 21896 18326
rect 1946 18224 1952 18276
rect 2004 18264 2010 18276
rect 6917 18267 6975 18273
rect 2004 18236 6500 18264
rect 2004 18224 2010 18236
rect 6472 18196 6500 18236
rect 6917 18233 6929 18267
rect 6963 18264 6975 18267
rect 7098 18264 7104 18276
rect 6963 18236 7104 18264
rect 6963 18233 6975 18236
rect 6917 18227 6975 18233
rect 7098 18224 7104 18236
rect 7156 18224 7162 18276
rect 9674 18264 9680 18276
rect 7208 18236 9680 18264
rect 7208 18196 7236 18236
rect 9674 18224 9680 18236
rect 9732 18224 9738 18276
rect 12069 18267 12127 18273
rect 12069 18233 12081 18267
rect 12115 18264 12127 18267
rect 12526 18264 12532 18276
rect 12115 18236 12532 18264
rect 12115 18233 12127 18236
rect 12069 18227 12127 18233
rect 12526 18224 12532 18236
rect 12584 18224 12590 18276
rect 12618 18224 12624 18276
rect 12676 18264 12682 18276
rect 13262 18264 13268 18276
rect 12676 18236 13268 18264
rect 12676 18224 12682 18236
rect 13262 18224 13268 18236
rect 13320 18224 13326 18276
rect 13630 18224 13636 18276
rect 13688 18264 13694 18276
rect 15378 18264 15384 18276
rect 13688 18236 15384 18264
rect 13688 18224 13694 18236
rect 15378 18224 15384 18236
rect 15436 18224 15442 18276
rect 15470 18224 15476 18276
rect 15528 18264 15534 18276
rect 16301 18267 16359 18273
rect 15528 18236 16252 18264
rect 15528 18224 15534 18236
rect 6472 18168 7236 18196
rect 7650 18156 7656 18208
rect 7708 18196 7714 18208
rect 10226 18196 10232 18208
rect 7708 18168 10232 18196
rect 7708 18156 7714 18168
rect 10226 18156 10232 18168
rect 10284 18156 10290 18208
rect 10318 18156 10324 18208
rect 10376 18196 10382 18208
rect 11698 18196 11704 18208
rect 10376 18168 11704 18196
rect 10376 18156 10382 18168
rect 11698 18156 11704 18168
rect 11756 18156 11762 18208
rect 13998 18156 14004 18208
rect 14056 18196 14062 18208
rect 16224 18196 16252 18236
rect 16301 18233 16313 18267
rect 16347 18264 16359 18267
rect 18598 18264 18604 18276
rect 16347 18236 18604 18264
rect 16347 18233 16359 18236
rect 16301 18227 16359 18233
rect 18598 18224 18604 18236
rect 18656 18224 18662 18276
rect 16482 18196 16488 18208
rect 14056 18168 16160 18196
rect 16224 18168 16488 18196
rect 14056 18156 14062 18168
rect 8297 18131 8355 18137
rect 8297 18128 8309 18131
rect 8220 18100 8309 18128
rect 5537 18063 5595 18069
rect 5537 18029 5549 18063
rect 5583 18029 5595 18063
rect 5537 18023 5595 18029
rect 5804 18063 5862 18069
rect 5804 18029 5816 18063
rect 5850 18060 5862 18063
rect 7650 18060 7656 18072
rect 5850 18032 7656 18060
rect 5850 18029 5862 18032
rect 5804 18023 5862 18029
rect 5552 17992 5580 18023
rect 7650 18020 7656 18032
rect 7708 18060 7714 18072
rect 8220 18060 8248 18100
rect 8297 18097 8309 18100
rect 8343 18097 8355 18131
rect 9858 18128 9864 18140
rect 9819 18100 9864 18128
rect 8297 18091 8355 18097
rect 9858 18088 9864 18100
rect 9916 18088 9922 18140
rect 13354 18128 13360 18140
rect 12452 18100 13360 18128
rect 7708 18032 8248 18060
rect 7708 18020 7714 18032
rect 8386 18020 8392 18072
rect 8444 18060 8450 18072
rect 10686 18060 10692 18072
rect 8444 18032 10692 18060
rect 8444 18020 8450 18032
rect 10686 18020 10692 18032
rect 10744 18020 10750 18072
rect 10870 18020 10876 18072
rect 10928 18060 10934 18072
rect 11885 18063 11943 18069
rect 11885 18060 11897 18063
rect 10928 18032 11897 18060
rect 10928 18020 10934 18032
rect 11885 18029 11897 18032
rect 11931 18029 11943 18063
rect 11885 18023 11943 18029
rect 6270 17992 6276 18004
rect 5552 17964 6276 17992
rect 6270 17952 6276 17964
rect 6328 17952 6334 18004
rect 7374 17952 7380 18004
rect 7432 17992 7438 18004
rect 8113 17995 8171 18001
rect 8113 17992 8125 17995
rect 7432 17964 8125 17992
rect 7432 17952 7438 17964
rect 8113 17961 8125 17964
rect 8159 17961 8171 17995
rect 8113 17955 8171 17961
rect 8570 17952 8576 18004
rect 8628 17992 8634 18004
rect 12452 17992 12480 18100
rect 13354 18088 13360 18100
rect 13412 18088 13418 18140
rect 16132 18128 16160 18168
rect 16482 18156 16488 18168
rect 16540 18156 16546 18208
rect 18230 18156 18236 18208
rect 18288 18196 18294 18208
rect 18874 18196 18880 18208
rect 18288 18168 18880 18196
rect 18288 18156 18294 18168
rect 18874 18156 18880 18168
rect 18932 18156 18938 18208
rect 18966 18128 18972 18140
rect 16132 18100 17356 18128
rect 12989 18063 13047 18069
rect 12989 18029 13001 18063
rect 13035 18060 13047 18063
rect 13906 18060 13912 18072
rect 13035 18032 13912 18060
rect 13035 18029 13047 18032
rect 12989 18023 13047 18029
rect 13906 18020 13912 18032
rect 13964 18020 13970 18072
rect 14093 18063 14151 18069
rect 14093 18029 14105 18063
rect 14139 18029 14151 18063
rect 14093 18023 14151 18029
rect 13630 17992 13636 18004
rect 8628 17964 12480 17992
rect 13096 17964 13636 17992
rect 8628 17952 8634 17964
rect 3050 17884 3056 17936
rect 3108 17924 3114 17936
rect 7282 17924 7288 17936
rect 3108 17896 7288 17924
rect 3108 17884 3114 17896
rect 7282 17884 7288 17896
rect 7340 17884 7346 17936
rect 7742 17924 7748 17936
rect 7703 17896 7748 17924
rect 7742 17884 7748 17896
rect 7800 17884 7806 17936
rect 8202 17924 8208 17936
rect 8163 17896 8208 17924
rect 8202 17884 8208 17896
rect 8260 17884 8266 17936
rect 8294 17884 8300 17936
rect 8352 17924 8358 17936
rect 10778 17924 10784 17936
rect 8352 17896 10784 17924
rect 8352 17884 8358 17896
rect 10778 17884 10784 17896
rect 10836 17884 10842 17936
rect 10873 17927 10931 17933
rect 10873 17893 10885 17927
rect 10919 17924 10931 17927
rect 11146 17924 11152 17936
rect 10919 17896 11152 17924
rect 10919 17893 10931 17896
rect 10873 17887 10931 17893
rect 11146 17884 11152 17896
rect 11204 17884 11210 17936
rect 11238 17884 11244 17936
rect 11296 17924 11302 17936
rect 13096 17924 13124 17964
rect 13630 17952 13636 17964
rect 13688 17952 13694 18004
rect 14108 17992 14136 18023
rect 14274 18020 14280 18072
rect 14332 18060 14338 18072
rect 14734 18060 14740 18072
rect 14332 18032 14740 18060
rect 14332 18020 14338 18032
rect 14734 18020 14740 18032
rect 14792 18020 14798 18072
rect 16117 18063 16175 18069
rect 16117 18029 16129 18063
rect 16163 18060 16175 18063
rect 17034 18060 17040 18072
rect 16163 18032 17040 18060
rect 16163 18029 16175 18032
rect 16117 18023 16175 18029
rect 17034 18020 17040 18032
rect 17092 18020 17098 18072
rect 17218 18060 17224 18072
rect 17179 18032 17224 18060
rect 17218 18020 17224 18032
rect 17276 18020 17282 18072
rect 17328 18060 17356 18100
rect 18248 18100 18972 18128
rect 18248 18060 18276 18100
rect 18966 18088 18972 18100
rect 19024 18088 19030 18140
rect 19058 18088 19064 18140
rect 19116 18088 19122 18140
rect 19886 18088 19892 18140
rect 19944 18128 19950 18140
rect 20346 18128 20352 18140
rect 19944 18100 20352 18128
rect 19944 18088 19950 18100
rect 20346 18088 20352 18100
rect 20404 18088 20410 18140
rect 17328 18032 18276 18060
rect 18874 18020 18880 18072
rect 18932 18060 18938 18072
rect 19076 18060 19104 18088
rect 19702 18060 19708 18072
rect 18932 18032 19104 18060
rect 19663 18032 19708 18060
rect 18932 18020 18938 18032
rect 19702 18020 19708 18032
rect 19760 18020 19766 18072
rect 17310 17992 17316 18004
rect 14108 17964 17316 17992
rect 17310 17952 17316 17964
rect 17368 17952 17374 18004
rect 17494 18001 17500 18004
rect 17488 17992 17500 18001
rect 17455 17964 17500 17992
rect 17488 17955 17500 17964
rect 17494 17952 17500 17955
rect 17552 17952 17558 18004
rect 17678 17952 17684 18004
rect 17736 17992 17742 18004
rect 18690 17992 18696 18004
rect 17736 17964 18696 17992
rect 17736 17952 17742 17964
rect 18690 17952 18696 17964
rect 18748 17952 18754 18004
rect 19610 17952 19616 18004
rect 19668 17992 19674 18004
rect 20438 17992 20444 18004
rect 19668 17964 20444 17992
rect 19668 17952 19674 17964
rect 20438 17952 20444 17964
rect 20496 17952 20502 18004
rect 11296 17896 13124 17924
rect 13173 17927 13231 17933
rect 11296 17884 11302 17896
rect 13173 17893 13185 17927
rect 13219 17924 13231 17927
rect 13998 17924 14004 17936
rect 13219 17896 14004 17924
rect 13219 17893 13231 17896
rect 13173 17887 13231 17893
rect 13998 17884 14004 17896
rect 14056 17884 14062 17936
rect 14277 17927 14335 17933
rect 14277 17893 14289 17927
rect 14323 17924 14335 17927
rect 18230 17924 18236 17936
rect 14323 17896 18236 17924
rect 14323 17893 14335 17896
rect 14277 17887 14335 17893
rect 18230 17884 18236 17896
rect 18288 17884 18294 17936
rect 18598 17924 18604 17936
rect 18559 17896 18604 17924
rect 18598 17884 18604 17896
rect 18656 17884 18662 17936
rect 19150 17884 19156 17936
rect 19208 17924 19214 17936
rect 19889 17927 19947 17933
rect 19889 17924 19901 17927
rect 19208 17896 19901 17924
rect 19208 17884 19214 17896
rect 19889 17893 19901 17896
rect 19935 17893 19947 17927
rect 19889 17887 19947 17893
rect 21174 17884 21180 17936
rect 21232 17924 21238 17936
rect 22646 17924 22652 17936
rect 21232 17896 22652 17924
rect 21232 17884 21238 17896
rect 22646 17884 22652 17896
rect 22704 17884 22710 17936
rect 1104 17834 21896 17856
rect 1104 17782 7912 17834
rect 7964 17782 7976 17834
rect 8028 17782 8040 17834
rect 8092 17782 8104 17834
rect 8156 17782 14843 17834
rect 14895 17782 14907 17834
rect 14959 17782 14971 17834
rect 15023 17782 15035 17834
rect 15087 17782 21896 17834
rect 1104 17760 21896 17782
rect 6917 17723 6975 17729
rect 6917 17689 6929 17723
rect 6963 17720 6975 17723
rect 8202 17720 8208 17732
rect 6963 17692 8208 17720
rect 6963 17689 6975 17692
rect 6917 17683 6975 17689
rect 8202 17680 8208 17692
rect 8260 17680 8266 17732
rect 9490 17680 9496 17732
rect 9548 17720 9554 17732
rect 9677 17723 9735 17729
rect 9677 17720 9689 17723
rect 9548 17692 9689 17720
rect 9548 17680 9554 17692
rect 9677 17689 9689 17692
rect 9723 17689 9735 17723
rect 9677 17683 9735 17689
rect 11333 17723 11391 17729
rect 11333 17689 11345 17723
rect 11379 17720 11391 17723
rect 12710 17720 12716 17732
rect 11379 17692 12716 17720
rect 11379 17689 11391 17692
rect 11333 17683 11391 17689
rect 12710 17680 12716 17692
rect 12768 17680 12774 17732
rect 12897 17723 12955 17729
rect 12897 17689 12909 17723
rect 12943 17720 12955 17723
rect 13078 17720 13084 17732
rect 12943 17692 13084 17720
rect 12943 17689 12955 17692
rect 12897 17683 12955 17689
rect 13078 17680 13084 17692
rect 13136 17680 13142 17732
rect 13354 17680 13360 17732
rect 13412 17720 13418 17732
rect 15013 17723 15071 17729
rect 15013 17720 15025 17723
rect 13412 17692 15025 17720
rect 13412 17680 13418 17692
rect 15013 17689 15025 17692
rect 15059 17689 15071 17723
rect 15013 17683 15071 17689
rect 18046 17680 18052 17732
rect 18104 17720 18110 17732
rect 18601 17723 18659 17729
rect 18601 17720 18613 17723
rect 18104 17692 18613 17720
rect 18104 17680 18110 17692
rect 18601 17689 18613 17692
rect 18647 17689 18659 17723
rect 18601 17683 18659 17689
rect 7006 17612 7012 17664
rect 7064 17652 7070 17664
rect 7377 17655 7435 17661
rect 7377 17652 7389 17655
rect 7064 17624 7389 17652
rect 7064 17612 7070 17624
rect 7377 17621 7389 17624
rect 7423 17621 7435 17655
rect 7377 17615 7435 17621
rect 7484 17624 16528 17652
rect 7190 17544 7196 17596
rect 7248 17584 7254 17596
rect 7285 17587 7343 17593
rect 7285 17584 7297 17587
rect 7248 17556 7297 17584
rect 7248 17544 7254 17556
rect 7285 17553 7297 17556
rect 7331 17553 7343 17587
rect 7484 17584 7512 17624
rect 7285 17547 7343 17553
rect 7392 17556 7512 17584
rect 4062 17476 4068 17528
rect 4120 17516 4126 17528
rect 7392 17516 7420 17556
rect 8938 17544 8944 17596
rect 8996 17584 9002 17596
rect 9582 17584 9588 17596
rect 8996 17556 9588 17584
rect 8996 17544 9002 17556
rect 9582 17544 9588 17556
rect 9640 17544 9646 17596
rect 12805 17587 12863 17593
rect 12805 17553 12817 17587
rect 12851 17584 12863 17587
rect 13170 17584 13176 17596
rect 12851 17556 13176 17584
rect 12851 17553 12863 17556
rect 12805 17547 12863 17553
rect 13170 17544 13176 17556
rect 13228 17544 13234 17596
rect 14921 17587 14979 17593
rect 14921 17553 14933 17587
rect 14967 17584 14979 17587
rect 15838 17584 15844 17596
rect 14967 17556 15844 17584
rect 14967 17553 14979 17556
rect 14921 17547 14979 17553
rect 15838 17544 15844 17556
rect 15896 17584 15902 17596
rect 16022 17584 16028 17596
rect 15896 17556 16028 17584
rect 15896 17544 15902 17556
rect 16022 17544 16028 17556
rect 16080 17544 16086 17596
rect 4120 17488 7420 17516
rect 4120 17476 4126 17488
rect 7466 17476 7472 17528
rect 7524 17516 7530 17528
rect 9766 17516 9772 17528
rect 7524 17488 7569 17516
rect 9727 17488 9772 17516
rect 7524 17476 7530 17488
rect 9766 17476 9772 17488
rect 9824 17476 9830 17528
rect 12986 17516 12992 17528
rect 12947 17488 12992 17516
rect 12986 17476 12992 17488
rect 13044 17476 13050 17528
rect 15102 17516 15108 17528
rect 15063 17488 15108 17516
rect 15102 17476 15108 17488
rect 15160 17476 15166 17528
rect 16500 17516 16528 17624
rect 17034 17612 17040 17664
rect 17092 17652 17098 17664
rect 20165 17655 20223 17661
rect 20165 17652 20177 17655
rect 17092 17624 20177 17652
rect 17092 17612 17098 17624
rect 20165 17621 20177 17624
rect 20211 17621 20223 17655
rect 20165 17615 20223 17621
rect 16850 17584 16856 17596
rect 16811 17556 16856 17584
rect 16850 17544 16856 17556
rect 16908 17544 16914 17596
rect 17862 17544 17868 17596
rect 17920 17584 17926 17596
rect 18509 17587 18567 17593
rect 18509 17584 18521 17587
rect 17920 17556 18521 17584
rect 17920 17544 17926 17556
rect 18509 17553 18521 17556
rect 18555 17553 18567 17587
rect 19886 17584 19892 17596
rect 19847 17556 19892 17584
rect 18509 17547 18567 17553
rect 19886 17544 19892 17556
rect 19944 17544 19950 17596
rect 18598 17516 18604 17528
rect 16500 17488 18604 17516
rect 18598 17476 18604 17488
rect 18656 17516 18662 17528
rect 18693 17519 18751 17525
rect 18693 17516 18705 17519
rect 18656 17488 18705 17516
rect 18656 17476 18662 17488
rect 18693 17485 18705 17488
rect 18739 17485 18751 17519
rect 18693 17479 18751 17485
rect 9858 17408 9864 17460
rect 9916 17448 9922 17460
rect 17862 17448 17868 17460
rect 9916 17420 17868 17448
rect 9916 17408 9922 17420
rect 17862 17408 17868 17420
rect 17920 17408 17926 17460
rect 18138 17448 18144 17460
rect 18099 17420 18144 17448
rect 18138 17408 18144 17420
rect 18196 17408 18202 17460
rect 9217 17383 9275 17389
rect 9217 17349 9229 17383
rect 9263 17380 9275 17383
rect 10502 17380 10508 17392
rect 9263 17352 10508 17380
rect 9263 17349 9275 17352
rect 9217 17343 9275 17349
rect 10502 17340 10508 17352
rect 10560 17340 10566 17392
rect 12434 17340 12440 17392
rect 12492 17380 12498 17392
rect 14553 17383 14611 17389
rect 12492 17352 12537 17380
rect 12492 17340 12498 17352
rect 14553 17349 14565 17383
rect 14599 17380 14611 17383
rect 15746 17380 15752 17392
rect 14599 17352 15752 17380
rect 14599 17349 14611 17352
rect 14553 17343 14611 17349
rect 15746 17340 15752 17352
rect 15804 17340 15810 17392
rect 17037 17383 17095 17389
rect 17037 17349 17049 17383
rect 17083 17380 17095 17383
rect 17954 17380 17960 17392
rect 17083 17352 17960 17380
rect 17083 17349 17095 17352
rect 17037 17343 17095 17349
rect 17954 17340 17960 17352
rect 18012 17340 18018 17392
rect 20990 17340 20996 17392
rect 21048 17380 21054 17392
rect 22094 17380 22100 17392
rect 21048 17352 22100 17380
rect 21048 17340 21054 17352
rect 22094 17340 22100 17352
rect 22152 17340 22158 17392
rect 1104 17290 21896 17312
rect 1104 17238 4447 17290
rect 4499 17238 4511 17290
rect 4563 17238 4575 17290
rect 4627 17238 4639 17290
rect 4691 17238 11378 17290
rect 11430 17238 11442 17290
rect 11494 17238 11506 17290
rect 11558 17238 11570 17290
rect 11622 17238 18308 17290
rect 18360 17238 18372 17290
rect 18424 17238 18436 17290
rect 18488 17238 18500 17290
rect 18552 17238 21896 17290
rect 1104 17216 21896 17238
rect 7650 17176 7656 17188
rect 7611 17148 7656 17176
rect 7650 17136 7656 17148
rect 7708 17136 7714 17188
rect 14369 17179 14427 17185
rect 14369 17145 14381 17179
rect 14415 17176 14427 17179
rect 15102 17176 15108 17188
rect 14415 17148 15108 17176
rect 14415 17145 14427 17148
rect 14369 17139 14427 17145
rect 15102 17136 15108 17148
rect 15160 17136 15166 17188
rect 18138 17136 18144 17188
rect 18196 17176 18202 17188
rect 18782 17176 18788 17188
rect 18196 17148 18788 17176
rect 18196 17136 18202 17148
rect 18782 17136 18788 17148
rect 18840 17136 18846 17188
rect 11885 17111 11943 17117
rect 11885 17077 11897 17111
rect 11931 17108 11943 17111
rect 12986 17108 12992 17120
rect 11931 17080 12992 17108
rect 11931 17077 11943 17080
rect 11885 17071 11943 17077
rect 12986 17068 12992 17080
rect 13044 17068 13050 17120
rect 15120 17040 15148 17136
rect 15120 17012 15424 17040
rect 6270 16972 6276 16984
rect 6231 16944 6276 16972
rect 6270 16932 6276 16944
rect 6328 16932 6334 16984
rect 6540 16975 6598 16981
rect 6540 16941 6552 16975
rect 6586 16972 6598 16975
rect 7098 16972 7104 16984
rect 6586 16944 7104 16972
rect 6586 16941 6598 16944
rect 6540 16935 6598 16941
rect 7098 16932 7104 16944
rect 7156 16972 7162 16984
rect 7466 16972 7472 16984
rect 7156 16944 7472 16972
rect 7156 16932 7162 16944
rect 7466 16932 7472 16944
rect 7524 16932 7530 16984
rect 9122 16932 9128 16984
rect 9180 16972 9186 16984
rect 10505 16975 10563 16981
rect 10505 16972 10517 16975
rect 9180 16944 10517 16972
rect 9180 16932 9186 16944
rect 10505 16941 10517 16944
rect 10551 16941 10563 16975
rect 10505 16935 10563 16941
rect 11238 16932 11244 16984
rect 11296 16972 11302 16984
rect 12897 16975 12955 16981
rect 12897 16972 12909 16975
rect 11296 16944 12909 16972
rect 11296 16932 11302 16944
rect 12897 16941 12909 16944
rect 12943 16941 12955 16975
rect 12897 16935 12955 16941
rect 12989 16975 13047 16981
rect 12989 16941 13001 16975
rect 13035 16972 13047 16975
rect 15286 16972 15292 16984
rect 13035 16944 15292 16972
rect 13035 16941 13047 16944
rect 12989 16935 13047 16941
rect 10594 16864 10600 16916
rect 10652 16904 10658 16916
rect 10750 16907 10808 16913
rect 10750 16904 10762 16907
rect 10652 16876 10762 16904
rect 10652 16864 10658 16876
rect 10750 16873 10762 16876
rect 10796 16873 10808 16907
rect 10750 16867 10808 16873
rect 12526 16796 12532 16848
rect 12584 16836 12590 16848
rect 12713 16839 12771 16845
rect 12713 16836 12725 16839
rect 12584 16808 12725 16836
rect 12584 16796 12590 16808
rect 12713 16805 12725 16808
rect 12759 16836 12771 16839
rect 13004 16836 13032 16935
rect 15286 16932 15292 16944
rect 15344 16932 15350 16984
rect 15396 16972 15424 17012
rect 16850 17000 16856 17052
rect 16908 17040 16914 17052
rect 19705 17043 19763 17049
rect 19705 17040 19717 17043
rect 16908 17012 19717 17040
rect 16908 17000 16914 17012
rect 19705 17009 19717 17012
rect 19751 17009 19763 17043
rect 19705 17003 19763 17009
rect 15545 16975 15603 16981
rect 15545 16972 15557 16975
rect 15396 16944 15557 16972
rect 15545 16941 15557 16944
rect 15591 16941 15603 16975
rect 15545 16935 15603 16941
rect 18417 16975 18475 16981
rect 18417 16941 18429 16975
rect 18463 16972 18475 16975
rect 19058 16972 19064 16984
rect 18463 16944 19064 16972
rect 18463 16941 18475 16944
rect 18417 16935 18475 16941
rect 19058 16932 19064 16944
rect 19116 16932 19122 16984
rect 19518 16972 19524 16984
rect 19479 16944 19524 16972
rect 19518 16932 19524 16944
rect 19576 16932 19582 16984
rect 13256 16907 13314 16913
rect 13256 16873 13268 16907
rect 13302 16904 13314 16907
rect 13722 16904 13728 16916
rect 13302 16876 13728 16904
rect 13302 16873 13314 16876
rect 13256 16867 13314 16873
rect 13722 16864 13728 16876
rect 13780 16864 13786 16916
rect 15194 16864 15200 16916
rect 15252 16904 15258 16916
rect 18966 16904 18972 16916
rect 15252 16876 18972 16904
rect 15252 16864 15258 16876
rect 18966 16864 18972 16876
rect 19024 16864 19030 16916
rect 12759 16808 13032 16836
rect 12759 16805 12771 16808
rect 12713 16799 12771 16805
rect 16022 16796 16028 16848
rect 16080 16836 16086 16848
rect 16669 16839 16727 16845
rect 16669 16836 16681 16839
rect 16080 16808 16681 16836
rect 16080 16796 16086 16808
rect 16669 16805 16681 16808
rect 16715 16805 16727 16839
rect 16669 16799 16727 16805
rect 18601 16839 18659 16845
rect 18601 16805 18613 16839
rect 18647 16836 18659 16839
rect 19242 16836 19248 16848
rect 18647 16808 19248 16836
rect 18647 16805 18659 16808
rect 18601 16799 18659 16805
rect 19242 16796 19248 16808
rect 19300 16796 19306 16848
rect 1104 16746 21896 16768
rect 1104 16694 7912 16746
rect 7964 16694 7976 16746
rect 8028 16694 8040 16746
rect 8092 16694 8104 16746
rect 8156 16694 14843 16746
rect 14895 16694 14907 16746
rect 14959 16694 14971 16746
rect 15023 16694 15035 16746
rect 15087 16694 21896 16746
rect 1104 16672 21896 16694
rect 7374 16632 7380 16644
rect 7335 16604 7380 16632
rect 7374 16592 7380 16604
rect 7432 16592 7438 16644
rect 10505 16635 10563 16641
rect 9140 16604 9904 16632
rect 5258 16524 5264 16576
rect 5316 16564 5322 16576
rect 9140 16564 9168 16604
rect 5316 16536 9168 16564
rect 9392 16567 9450 16573
rect 5316 16524 5322 16536
rect 9392 16533 9404 16567
rect 9438 16564 9450 16567
rect 9766 16564 9772 16576
rect 9438 16536 9772 16564
rect 9438 16533 9450 16536
rect 9392 16527 9450 16533
rect 9766 16524 9772 16536
rect 9824 16524 9830 16576
rect 9876 16564 9904 16604
rect 10505 16601 10517 16635
rect 10551 16632 10563 16635
rect 10594 16632 10600 16644
rect 10551 16604 10600 16632
rect 10551 16601 10563 16604
rect 10505 16595 10563 16601
rect 10594 16592 10600 16604
rect 10652 16592 10658 16644
rect 11698 16592 11704 16644
rect 11756 16632 11762 16644
rect 11756 16604 13584 16632
rect 11756 16592 11762 16604
rect 13556 16564 13584 16604
rect 13722 16592 13728 16644
rect 13780 16632 13786 16644
rect 13817 16635 13875 16641
rect 13817 16632 13829 16635
rect 13780 16604 13829 16632
rect 13780 16592 13786 16604
rect 13817 16601 13829 16604
rect 13863 16601 13875 16635
rect 13817 16595 13875 16601
rect 14829 16635 14887 16641
rect 14829 16601 14841 16635
rect 14875 16632 14887 16635
rect 15194 16632 15200 16644
rect 14875 16604 15200 16632
rect 14875 16601 14887 16604
rect 14829 16595 14887 16601
rect 15194 16592 15200 16604
rect 15252 16592 15258 16644
rect 16574 16592 16580 16644
rect 16632 16632 16638 16644
rect 16632 16604 18644 16632
rect 16632 16592 16638 16604
rect 16022 16573 16028 16576
rect 16016 16564 16028 16573
rect 9876 16536 13492 16564
rect 13556 16536 14688 16564
rect 15983 16536 16028 16564
rect 9033 16499 9091 16505
rect 9033 16465 9045 16499
rect 9079 16496 9091 16499
rect 11238 16496 11244 16508
rect 9079 16468 11244 16496
rect 9079 16465 9091 16468
rect 9033 16459 9091 16465
rect 11238 16456 11244 16468
rect 11296 16456 11302 16508
rect 12437 16499 12495 16505
rect 12437 16465 12449 16499
rect 12483 16496 12495 16499
rect 12526 16496 12532 16508
rect 12483 16468 12532 16496
rect 12483 16465 12495 16468
rect 12437 16459 12495 16465
rect 12526 16456 12532 16468
rect 12584 16456 12590 16508
rect 12704 16499 12762 16505
rect 12704 16465 12716 16499
rect 12750 16496 12762 16499
rect 12986 16496 12992 16508
rect 12750 16468 12992 16496
rect 12750 16465 12762 16468
rect 12704 16459 12762 16465
rect 12986 16456 12992 16468
rect 13044 16456 13050 16508
rect 13464 16496 13492 16536
rect 14660 16505 14688 16536
rect 16016 16527 16028 16536
rect 16022 16524 16028 16527
rect 16080 16524 16086 16576
rect 18509 16567 18567 16573
rect 18509 16564 18521 16567
rect 16132 16536 18521 16564
rect 14645 16499 14703 16505
rect 13464 16468 14596 16496
rect 9122 16428 9128 16440
rect 8864 16400 9128 16428
rect 8386 16252 8392 16304
rect 8444 16292 8450 16304
rect 8864 16301 8892 16400
rect 9122 16388 9128 16400
rect 9180 16388 9186 16440
rect 11054 16388 11060 16440
rect 11112 16428 11118 16440
rect 11333 16431 11391 16437
rect 11333 16428 11345 16431
rect 11112 16400 11345 16428
rect 11112 16388 11118 16400
rect 11333 16397 11345 16400
rect 11379 16397 11391 16431
rect 14568 16428 14596 16468
rect 14645 16465 14657 16499
rect 14691 16465 14703 16499
rect 16132 16496 16160 16536
rect 18509 16533 18521 16536
rect 18555 16533 18567 16567
rect 18509 16527 18567 16533
rect 14645 16459 14703 16465
rect 14752 16468 16160 16496
rect 18417 16499 18475 16505
rect 14752 16428 14780 16468
rect 18417 16465 18429 16499
rect 18463 16465 18475 16499
rect 18616 16496 18644 16604
rect 19702 16524 19708 16576
rect 19760 16564 19766 16576
rect 20165 16567 20223 16573
rect 20165 16564 20177 16567
rect 19760 16536 20177 16564
rect 19760 16524 19766 16536
rect 20165 16533 20177 16536
rect 20211 16533 20223 16567
rect 20165 16527 20223 16533
rect 19889 16499 19947 16505
rect 19889 16496 19901 16499
rect 18616 16468 19901 16496
rect 18417 16459 18475 16465
rect 19889 16465 19901 16468
rect 19935 16465 19947 16499
rect 19889 16459 19947 16465
rect 14568 16400 14780 16428
rect 11333 16391 11391 16397
rect 15286 16388 15292 16440
rect 15344 16428 15350 16440
rect 15749 16431 15807 16437
rect 15749 16428 15761 16431
rect 15344 16400 15761 16428
rect 15344 16388 15350 16400
rect 15749 16397 15761 16400
rect 15795 16397 15807 16431
rect 18432 16428 18460 16459
rect 18506 16428 18512 16440
rect 18432 16400 18512 16428
rect 15749 16391 15807 16397
rect 8849 16295 8907 16301
rect 8849 16292 8861 16295
rect 8444 16264 8861 16292
rect 8444 16252 8450 16264
rect 8849 16261 8861 16264
rect 8895 16261 8907 16295
rect 15764 16292 15792 16391
rect 18506 16388 18512 16400
rect 18564 16388 18570 16440
rect 18601 16431 18659 16437
rect 18601 16397 18613 16431
rect 18647 16397 18659 16431
rect 18601 16391 18659 16397
rect 17129 16363 17187 16369
rect 17129 16329 17141 16363
rect 17175 16360 17187 16363
rect 17586 16360 17592 16372
rect 17175 16332 17592 16360
rect 17175 16329 17187 16332
rect 17129 16323 17187 16329
rect 17586 16320 17592 16332
rect 17644 16360 17650 16372
rect 18616 16360 18644 16391
rect 17644 16332 18644 16360
rect 17644 16320 17650 16332
rect 17310 16292 17316 16304
rect 15764 16264 17316 16292
rect 8849 16255 8907 16261
rect 17310 16252 17316 16264
rect 17368 16252 17374 16304
rect 18046 16292 18052 16304
rect 18007 16264 18052 16292
rect 18046 16252 18052 16264
rect 18104 16252 18110 16304
rect 1104 16202 21896 16224
rect 1104 16150 4447 16202
rect 4499 16150 4511 16202
rect 4563 16150 4575 16202
rect 4627 16150 4639 16202
rect 4691 16150 11378 16202
rect 11430 16150 11442 16202
rect 11494 16150 11506 16202
rect 11558 16150 11570 16202
rect 11622 16150 18308 16202
rect 18360 16150 18372 16202
rect 18424 16150 18436 16202
rect 18488 16150 18500 16202
rect 18552 16150 21896 16202
rect 1104 16128 21896 16150
rect 7098 16088 7104 16100
rect 7059 16060 7104 16088
rect 7098 16048 7104 16060
rect 7156 16048 7162 16100
rect 15565 16091 15623 16097
rect 15565 16057 15577 16091
rect 15611 16088 15623 16091
rect 19518 16088 19524 16100
rect 15611 16060 19524 16088
rect 15611 16057 15623 16060
rect 15565 16051 15623 16057
rect 19518 16048 19524 16060
rect 19576 16048 19582 16100
rect 10137 16023 10195 16029
rect 10137 15989 10149 16023
rect 10183 16020 10195 16023
rect 12618 16020 12624 16032
rect 10183 15992 12624 16020
rect 10183 15989 10195 15992
rect 10137 15983 10195 15989
rect 12618 15980 12624 15992
rect 12676 15980 12682 16032
rect 12805 16023 12863 16029
rect 12805 15989 12817 16023
rect 12851 16020 12863 16023
rect 16574 16020 16580 16032
rect 12851 15992 16580 16020
rect 12851 15989 12863 15992
rect 12805 15983 12863 15989
rect 16574 15980 16580 15992
rect 16632 15980 16638 16032
rect 10594 15912 10600 15964
rect 10652 15952 10658 15964
rect 10689 15955 10747 15961
rect 10689 15952 10701 15955
rect 10652 15924 10701 15952
rect 10652 15912 10658 15924
rect 10689 15921 10701 15924
rect 10735 15921 10747 15955
rect 10689 15915 10747 15921
rect 12434 15912 12440 15964
rect 12492 15952 12498 15964
rect 13265 15955 13323 15961
rect 13265 15952 13277 15955
rect 12492 15924 13277 15952
rect 12492 15912 12498 15924
rect 13265 15921 13277 15924
rect 13311 15921 13323 15955
rect 13265 15915 13323 15921
rect 13449 15955 13507 15961
rect 13449 15921 13461 15955
rect 13495 15952 13507 15955
rect 13722 15952 13728 15964
rect 13495 15924 13728 15952
rect 13495 15921 13507 15924
rect 13449 15915 13507 15921
rect 13722 15912 13728 15924
rect 13780 15912 13786 15964
rect 16022 15912 16028 15964
rect 16080 15952 16086 15964
rect 16117 15955 16175 15961
rect 16117 15952 16129 15955
rect 16080 15924 16129 15952
rect 16080 15912 16086 15924
rect 16117 15921 16129 15924
rect 16163 15921 16175 15955
rect 16117 15915 16175 15921
rect 5721 15887 5779 15893
rect 5721 15853 5733 15887
rect 5767 15884 5779 15887
rect 6270 15884 6276 15896
rect 5767 15856 6276 15884
rect 5767 15853 5779 15856
rect 5721 15847 5779 15853
rect 6270 15844 6276 15856
rect 6328 15844 6334 15896
rect 10505 15887 10563 15893
rect 10505 15853 10517 15887
rect 10551 15884 10563 15887
rect 11054 15884 11060 15896
rect 10551 15856 11060 15884
rect 10551 15853 10563 15856
rect 10505 15847 10563 15853
rect 11054 15844 11060 15856
rect 11112 15844 11118 15896
rect 12710 15844 12716 15896
rect 12768 15884 12774 15896
rect 13173 15887 13231 15893
rect 13173 15884 13185 15887
rect 12768 15856 13185 15884
rect 12768 15844 12774 15856
rect 13173 15853 13185 15856
rect 13219 15853 13231 15887
rect 17310 15884 17316 15896
rect 13173 15847 13231 15853
rect 15672 15856 16620 15884
rect 17271 15856 17316 15884
rect 5988 15819 6046 15825
rect 5988 15785 6000 15819
rect 6034 15816 6046 15819
rect 15672 15816 15700 15856
rect 6034 15788 15700 15816
rect 6034 15785 6046 15788
rect 5988 15779 6046 15785
rect 15746 15776 15752 15828
rect 15804 15816 15810 15828
rect 16025 15819 16083 15825
rect 16025 15816 16037 15819
rect 15804 15788 16037 15816
rect 15804 15776 15810 15788
rect 16025 15785 16037 15788
rect 16071 15785 16083 15819
rect 16025 15779 16083 15785
rect 10502 15708 10508 15760
rect 10560 15748 10566 15760
rect 10597 15751 10655 15757
rect 10597 15748 10609 15751
rect 10560 15720 10609 15748
rect 10560 15708 10566 15720
rect 10597 15717 10609 15720
rect 10643 15717 10655 15751
rect 10597 15711 10655 15717
rect 15838 15708 15844 15760
rect 15896 15748 15902 15760
rect 15933 15751 15991 15757
rect 15933 15748 15945 15751
rect 15896 15720 15945 15748
rect 15896 15708 15902 15720
rect 15933 15717 15945 15720
rect 15979 15717 15991 15751
rect 16592 15748 16620 15856
rect 17310 15844 17316 15856
rect 17368 15844 17374 15896
rect 17586 15893 17592 15896
rect 17580 15884 17592 15893
rect 17547 15856 17592 15884
rect 17580 15847 17592 15856
rect 17586 15844 17592 15847
rect 17644 15844 17650 15896
rect 19518 15884 19524 15896
rect 19479 15856 19524 15884
rect 19518 15844 19524 15856
rect 19576 15844 19582 15896
rect 17678 15776 17684 15828
rect 17736 15816 17742 15828
rect 19797 15819 19855 15825
rect 19797 15816 19809 15819
rect 17736 15788 19809 15816
rect 17736 15776 17742 15788
rect 19797 15785 19809 15788
rect 19843 15785 19855 15819
rect 19797 15779 19855 15785
rect 18693 15751 18751 15757
rect 18693 15748 18705 15751
rect 16592 15720 18705 15748
rect 15933 15711 15991 15717
rect 18693 15717 18705 15720
rect 18739 15748 18751 15751
rect 18782 15748 18788 15760
rect 18739 15720 18788 15748
rect 18739 15717 18751 15720
rect 18693 15711 18751 15717
rect 18782 15708 18788 15720
rect 18840 15708 18846 15760
rect 1104 15658 21896 15680
rect 1104 15606 7912 15658
rect 7964 15606 7976 15658
rect 8028 15606 8040 15658
rect 8092 15606 8104 15658
rect 8156 15606 14843 15658
rect 14895 15606 14907 15658
rect 14959 15606 14971 15658
rect 15023 15606 15035 15658
rect 15087 15606 21896 15658
rect 1104 15584 21896 15606
rect 7282 15544 7288 15556
rect 7243 15516 7288 15544
rect 7282 15504 7288 15516
rect 7340 15504 7346 15556
rect 9766 15544 9772 15556
rect 9727 15516 9772 15544
rect 9766 15504 9772 15516
rect 9824 15504 9830 15556
rect 11238 15504 11244 15556
rect 11296 15544 11302 15556
rect 11609 15547 11667 15553
rect 11609 15544 11621 15547
rect 11296 15516 11621 15544
rect 11296 15504 11302 15516
rect 11609 15513 11621 15516
rect 11655 15513 11667 15547
rect 11609 15507 11667 15513
rect 12618 15504 12624 15556
rect 12676 15544 12682 15556
rect 15838 15544 15844 15556
rect 12676 15516 14412 15544
rect 15799 15516 15844 15544
rect 12676 15504 12682 15516
rect 7193 15479 7251 15485
rect 7193 15445 7205 15479
rect 7239 15476 7251 15479
rect 7558 15476 7564 15488
rect 7239 15448 7564 15476
rect 7239 15445 7251 15448
rect 7193 15439 7251 15445
rect 7558 15436 7564 15448
rect 7616 15476 7622 15488
rect 7616 15448 9536 15476
rect 7616 15436 7622 15448
rect 8662 15417 8668 15420
rect 8656 15408 8668 15417
rect 8623 15380 8668 15408
rect 8656 15371 8668 15380
rect 8662 15368 8668 15371
rect 8720 15368 8726 15420
rect 9508 15408 9536 15448
rect 9582 15436 9588 15488
rect 9640 15476 9646 15488
rect 14384 15476 14412 15516
rect 15838 15504 15844 15516
rect 15896 15504 15902 15556
rect 17037 15547 17095 15553
rect 17037 15513 17049 15547
rect 17083 15544 17095 15547
rect 17954 15544 17960 15556
rect 17083 15516 17960 15544
rect 17083 15513 17095 15516
rect 17037 15507 17095 15513
rect 17954 15504 17960 15516
rect 18012 15504 18018 15556
rect 18046 15504 18052 15556
rect 18104 15544 18110 15556
rect 18693 15547 18751 15553
rect 18693 15544 18705 15547
rect 18104 15516 18705 15544
rect 18104 15504 18110 15516
rect 18693 15513 18705 15516
rect 18739 15513 18751 15547
rect 18693 15507 18751 15513
rect 19426 15476 19432 15488
rect 9640 15448 14320 15476
rect 14384 15448 19432 15476
rect 9640 15436 9646 15448
rect 10502 15408 10508 15420
rect 9508 15380 10508 15408
rect 10502 15368 10508 15380
rect 10560 15368 10566 15420
rect 11793 15411 11851 15417
rect 11793 15377 11805 15411
rect 11839 15408 11851 15411
rect 13078 15408 13084 15420
rect 11839 15380 13084 15408
rect 11839 15377 11851 15380
rect 11793 15371 11851 15377
rect 13078 15368 13084 15380
rect 13136 15368 13142 15420
rect 14292 15417 14320 15448
rect 19426 15436 19432 15448
rect 19484 15436 19490 15488
rect 14277 15411 14335 15417
rect 14277 15377 14289 15411
rect 14323 15408 14335 15411
rect 15194 15408 15200 15420
rect 14323 15380 15200 15408
rect 14323 15377 14335 15380
rect 14277 15371 14335 15377
rect 15194 15368 15200 15380
rect 15252 15368 15258 15420
rect 16853 15411 16911 15417
rect 16853 15377 16865 15411
rect 16899 15408 16911 15411
rect 17678 15408 17684 15420
rect 16899 15380 17684 15408
rect 16899 15377 16911 15380
rect 16853 15371 16911 15377
rect 17678 15368 17684 15380
rect 17736 15368 17742 15420
rect 18601 15411 18659 15417
rect 18601 15377 18613 15411
rect 18647 15408 18659 15411
rect 19242 15408 19248 15420
rect 18647 15380 19248 15408
rect 18647 15377 18659 15380
rect 18601 15371 18659 15377
rect 19242 15368 19248 15380
rect 19300 15368 19306 15420
rect 19978 15408 19984 15420
rect 19939 15380 19984 15408
rect 19978 15368 19984 15380
rect 20036 15368 20042 15420
rect 7466 15340 7472 15352
rect 7427 15312 7472 15340
rect 7466 15300 7472 15312
rect 7524 15300 7530 15352
rect 8386 15340 8392 15352
rect 8347 15312 8392 15340
rect 8386 15300 8392 15312
rect 8444 15300 8450 15352
rect 10594 15340 10600 15352
rect 10555 15312 10600 15340
rect 10594 15300 10600 15312
rect 10652 15300 10658 15352
rect 13446 15300 13452 15352
rect 13504 15340 13510 15352
rect 14369 15343 14427 15349
rect 14369 15340 14381 15343
rect 13504 15312 14381 15340
rect 13504 15300 13510 15312
rect 14369 15309 14381 15312
rect 14415 15309 14427 15343
rect 14550 15340 14556 15352
rect 14511 15312 14556 15340
rect 14369 15303 14427 15309
rect 14550 15300 14556 15312
rect 14608 15300 14614 15352
rect 18782 15340 18788 15352
rect 18743 15312 18788 15340
rect 18782 15300 18788 15312
rect 18840 15300 18846 15352
rect 18874 15300 18880 15352
rect 18932 15340 18938 15352
rect 20165 15343 20223 15349
rect 20165 15340 20177 15343
rect 18932 15312 20177 15340
rect 18932 15300 18938 15312
rect 20165 15309 20177 15312
rect 20211 15309 20223 15343
rect 20165 15303 20223 15309
rect 18233 15275 18291 15281
rect 18233 15241 18245 15275
rect 18279 15272 18291 15275
rect 19518 15272 19524 15284
rect 18279 15244 19524 15272
rect 18279 15241 18291 15244
rect 18233 15235 18291 15241
rect 19518 15232 19524 15244
rect 19576 15232 19582 15284
rect 6825 15207 6883 15213
rect 6825 15173 6837 15207
rect 6871 15204 6883 15207
rect 7742 15204 7748 15216
rect 6871 15176 7748 15204
rect 6871 15173 6883 15176
rect 6825 15167 6883 15173
rect 7742 15164 7748 15176
rect 7800 15164 7806 15216
rect 13906 15204 13912 15216
rect 13867 15176 13912 15204
rect 13906 15164 13912 15176
rect 13964 15164 13970 15216
rect 19334 15164 19340 15216
rect 19392 15204 19398 15216
rect 19886 15204 19892 15216
rect 19392 15176 19892 15204
rect 19392 15164 19398 15176
rect 19886 15164 19892 15176
rect 19944 15164 19950 15216
rect 1104 15114 21896 15136
rect 1104 15062 4447 15114
rect 4499 15062 4511 15114
rect 4563 15062 4575 15114
rect 4627 15062 4639 15114
rect 4691 15062 11378 15114
rect 11430 15062 11442 15114
rect 11494 15062 11506 15114
rect 11558 15062 11570 15114
rect 11622 15062 18308 15114
rect 18360 15062 18372 15114
rect 18424 15062 18436 15114
rect 18488 15062 18500 15114
rect 18552 15062 21896 15114
rect 1104 15040 21896 15062
rect 11241 15003 11299 15009
rect 11241 14969 11253 15003
rect 11287 15000 11299 15003
rect 13446 15000 13452 15012
rect 11287 14972 13452 15000
rect 11287 14969 11299 14972
rect 11241 14963 11299 14969
rect 13446 14960 13452 14972
rect 13504 14960 13510 15012
rect 17497 15003 17555 15009
rect 17497 14969 17509 15003
rect 17543 15000 17555 15003
rect 18690 15000 18696 15012
rect 17543 14972 18696 15000
rect 17543 14969 17555 14972
rect 17497 14963 17555 14969
rect 18690 14960 18696 14972
rect 18748 14960 18754 15012
rect 19426 14960 19432 15012
rect 19484 15000 19490 15012
rect 19484 14972 19564 15000
rect 19484 14960 19490 14972
rect 8662 14892 8668 14944
rect 8720 14932 8726 14944
rect 8757 14935 8815 14941
rect 8757 14932 8769 14935
rect 8720 14904 8769 14932
rect 8720 14892 8726 14904
rect 8757 14901 8769 14904
rect 8803 14901 8815 14935
rect 8757 14895 8815 14901
rect 9677 14935 9735 14941
rect 9677 14901 9689 14935
rect 9723 14932 9735 14935
rect 9723 14904 12388 14932
rect 9723 14901 9735 14904
rect 9677 14895 9735 14901
rect 8772 14864 8800 14895
rect 10229 14867 10287 14873
rect 10229 14864 10241 14867
rect 8772 14836 10241 14864
rect 10229 14833 10241 14836
rect 10275 14833 10287 14867
rect 10229 14827 10287 14833
rect 11146 14824 11152 14876
rect 11204 14864 11210 14876
rect 11701 14867 11759 14873
rect 11701 14864 11713 14867
rect 11204 14836 11713 14864
rect 11204 14824 11210 14836
rect 11701 14833 11713 14836
rect 11747 14833 11759 14867
rect 11882 14864 11888 14876
rect 11843 14836 11888 14864
rect 11701 14827 11759 14833
rect 11882 14824 11888 14836
rect 11940 14824 11946 14876
rect 6270 14756 6276 14808
rect 6328 14796 6334 14808
rect 7377 14799 7435 14805
rect 7377 14796 7389 14799
rect 6328 14768 7389 14796
rect 6328 14756 6334 14768
rect 7377 14765 7389 14768
rect 7423 14796 7435 14799
rect 8386 14796 8392 14808
rect 7423 14768 8392 14796
rect 7423 14765 7435 14768
rect 7377 14759 7435 14765
rect 8386 14756 8392 14768
rect 8444 14756 8450 14808
rect 10045 14799 10103 14805
rect 10045 14765 10057 14799
rect 10091 14796 10103 14799
rect 10594 14796 10600 14808
rect 10091 14768 10600 14796
rect 10091 14765 10103 14768
rect 10045 14759 10103 14765
rect 10594 14756 10600 14768
rect 10652 14756 10658 14808
rect 12360 14796 12388 14904
rect 12526 14824 12532 14876
rect 12584 14864 12590 14876
rect 12805 14867 12863 14873
rect 12805 14864 12817 14867
rect 12584 14836 12817 14864
rect 12584 14824 12590 14836
rect 12805 14833 12817 14836
rect 12851 14833 12863 14867
rect 12805 14827 12863 14833
rect 14550 14824 14556 14876
rect 14608 14864 14614 14876
rect 15841 14867 15899 14873
rect 15841 14864 15853 14867
rect 14608 14836 15853 14864
rect 14608 14824 14614 14836
rect 15841 14833 15853 14836
rect 15887 14833 15899 14867
rect 18874 14864 18880 14876
rect 15841 14827 15899 14833
rect 17328 14836 18880 14864
rect 13072 14799 13130 14805
rect 12360 14768 13032 14796
rect 7466 14688 7472 14740
rect 7524 14728 7530 14740
rect 7644 14731 7702 14737
rect 7644 14728 7656 14731
rect 7524 14700 7656 14728
rect 7524 14688 7530 14700
rect 7644 14697 7656 14700
rect 7690 14728 7702 14731
rect 8202 14728 8208 14740
rect 7690 14700 8208 14728
rect 7690 14697 7702 14700
rect 7644 14691 7702 14697
rect 8202 14688 8208 14700
rect 8260 14688 8266 14740
rect 13004 14728 13032 14768
rect 13072 14765 13084 14799
rect 13118 14796 13130 14799
rect 14568 14796 14596 14824
rect 17328 14805 17356 14836
rect 18874 14824 18880 14836
rect 18932 14824 18938 14876
rect 19058 14824 19064 14876
rect 19116 14864 19122 14876
rect 19426 14864 19432 14876
rect 19116 14836 19432 14864
rect 19116 14824 19122 14836
rect 19426 14824 19432 14836
rect 19484 14824 19490 14876
rect 13118 14768 14596 14796
rect 17313 14799 17371 14805
rect 13118 14765 13130 14768
rect 13072 14759 13130 14765
rect 17313 14765 17325 14799
rect 17359 14765 17371 14799
rect 17313 14759 17371 14765
rect 17402 14756 17408 14808
rect 17460 14796 17466 14808
rect 19536 14805 19564 14972
rect 19702 14864 19708 14876
rect 19663 14836 19708 14864
rect 19702 14824 19708 14836
rect 19760 14824 19766 14876
rect 18417 14799 18475 14805
rect 18417 14796 18429 14799
rect 17460 14768 18429 14796
rect 17460 14756 17466 14768
rect 18417 14765 18429 14768
rect 18463 14765 18475 14799
rect 18417 14759 18475 14765
rect 19531 14799 19589 14805
rect 19531 14765 19543 14799
rect 19577 14765 19589 14799
rect 19531 14759 19589 14765
rect 19334 14728 19340 14740
rect 13004 14700 19340 14728
rect 19334 14688 19340 14700
rect 19392 14688 19398 14740
rect 7742 14620 7748 14672
rect 7800 14660 7806 14672
rect 10137 14663 10195 14669
rect 10137 14660 10149 14663
rect 7800 14632 10149 14660
rect 7800 14620 7806 14632
rect 10137 14629 10149 14632
rect 10183 14629 10195 14663
rect 10137 14623 10195 14629
rect 11238 14620 11244 14672
rect 11296 14660 11302 14672
rect 11609 14663 11667 14669
rect 11609 14660 11621 14663
rect 11296 14632 11621 14660
rect 11296 14620 11302 14632
rect 11609 14629 11621 14632
rect 11655 14629 11667 14663
rect 14182 14660 14188 14672
rect 14143 14632 14188 14660
rect 11609 14623 11667 14629
rect 14182 14620 14188 14632
rect 14240 14620 14246 14672
rect 15286 14660 15292 14672
rect 15247 14632 15292 14660
rect 15286 14620 15292 14632
rect 15344 14620 15350 14672
rect 15654 14660 15660 14672
rect 15615 14632 15660 14660
rect 15654 14620 15660 14632
rect 15712 14620 15718 14672
rect 15749 14663 15807 14669
rect 15749 14629 15761 14663
rect 15795 14660 15807 14663
rect 15838 14660 15844 14672
rect 15795 14632 15844 14660
rect 15795 14629 15807 14632
rect 15749 14623 15807 14629
rect 15838 14620 15844 14632
rect 15896 14620 15902 14672
rect 18598 14660 18604 14672
rect 18559 14632 18604 14660
rect 18598 14620 18604 14632
rect 18656 14620 18662 14672
rect 1104 14570 21896 14592
rect 1104 14518 7912 14570
rect 7964 14518 7976 14570
rect 8028 14518 8040 14570
rect 8092 14518 8104 14570
rect 8156 14518 14843 14570
rect 14895 14518 14907 14570
rect 14959 14518 14971 14570
rect 15023 14518 15035 14570
rect 15087 14518 21896 14570
rect 1104 14496 21896 14518
rect 8202 14456 8208 14468
rect 8163 14428 8208 14456
rect 8202 14416 8208 14428
rect 8260 14416 8266 14468
rect 13817 14459 13875 14465
rect 13817 14425 13829 14459
rect 13863 14456 13875 14459
rect 14550 14456 14556 14468
rect 13863 14428 14556 14456
rect 13863 14425 13875 14428
rect 13817 14419 13875 14425
rect 14550 14416 14556 14428
rect 14608 14416 14614 14468
rect 14737 14459 14795 14465
rect 14737 14425 14749 14459
rect 14783 14456 14795 14459
rect 15654 14456 15660 14468
rect 14783 14428 15660 14456
rect 14783 14425 14795 14428
rect 14737 14419 14795 14425
rect 15654 14416 15660 14428
rect 15712 14416 15718 14468
rect 17129 14459 17187 14465
rect 17129 14425 17141 14459
rect 17175 14425 17187 14459
rect 19058 14456 19064 14468
rect 17129 14419 17187 14425
rect 18248 14428 19064 14456
rect 10220 14391 10278 14397
rect 6840 14360 8432 14388
rect 6840 14329 6868 14360
rect 8404 14332 8432 14360
rect 10220 14357 10232 14391
rect 10266 14388 10278 14391
rect 14182 14388 14188 14400
rect 10266 14360 14188 14388
rect 10266 14357 10278 14360
rect 10220 14351 10278 14357
rect 14182 14348 14188 14360
rect 14240 14348 14246 14400
rect 17144 14388 17172 14419
rect 14292 14360 17172 14388
rect 6825 14323 6883 14329
rect 6825 14289 6837 14323
rect 6871 14289 6883 14323
rect 6825 14283 6883 14289
rect 7092 14323 7150 14329
rect 7092 14289 7104 14323
rect 7138 14320 7150 14323
rect 7466 14320 7472 14332
rect 7138 14292 7472 14320
rect 7138 14289 7150 14292
rect 7092 14283 7150 14289
rect 7466 14280 7472 14292
rect 7524 14280 7530 14332
rect 8386 14280 8392 14332
rect 8444 14320 8450 14332
rect 9953 14323 10011 14329
rect 9953 14320 9965 14323
rect 8444 14292 9965 14320
rect 8444 14280 8450 14292
rect 9953 14289 9965 14292
rect 9999 14289 10011 14323
rect 9953 14283 10011 14289
rect 11882 14280 11888 14332
rect 11940 14320 11946 14332
rect 12704 14323 12762 14329
rect 12704 14320 12716 14323
rect 11940 14292 12716 14320
rect 11940 14280 11946 14292
rect 12704 14289 12716 14292
rect 12750 14320 12762 14323
rect 14292 14320 14320 14360
rect 12750 14292 14320 14320
rect 16016 14323 16074 14329
rect 12750 14289 12762 14292
rect 12704 14283 12762 14289
rect 16016 14289 16028 14323
rect 16062 14320 16074 14323
rect 18248 14320 18276 14428
rect 19058 14416 19064 14428
rect 19116 14456 19122 14468
rect 19429 14459 19487 14465
rect 19429 14456 19441 14459
rect 19116 14428 19441 14456
rect 19116 14416 19122 14428
rect 19429 14425 19441 14428
rect 19475 14425 19487 14459
rect 19429 14419 19487 14425
rect 16062 14292 18276 14320
rect 18316 14323 18374 14329
rect 16062 14289 16074 14292
rect 16016 14283 16074 14289
rect 18316 14289 18328 14323
rect 18362 14320 18374 14323
rect 19150 14320 19156 14332
rect 18362 14292 19156 14320
rect 18362 14289 18374 14292
rect 18316 14283 18374 14289
rect 19150 14280 19156 14292
rect 19208 14280 19214 14332
rect 20438 14280 20444 14332
rect 20496 14320 20502 14332
rect 20533 14323 20591 14329
rect 20533 14320 20545 14323
rect 20496 14292 20545 14320
rect 20496 14280 20502 14292
rect 20533 14289 20545 14292
rect 20579 14289 20591 14323
rect 20533 14283 20591 14289
rect 12437 14255 12495 14261
rect 12437 14221 12449 14255
rect 12483 14221 12495 14255
rect 12437 14215 12495 14221
rect 15749 14255 15807 14261
rect 15749 14221 15761 14255
rect 15795 14221 15807 14255
rect 15749 14215 15807 14221
rect 18049 14255 18107 14261
rect 18049 14221 18061 14255
rect 18095 14221 18107 14255
rect 18049 14215 18107 14221
rect 10870 14076 10876 14128
rect 10928 14116 10934 14128
rect 11333 14119 11391 14125
rect 11333 14116 11345 14119
rect 10928 14088 11345 14116
rect 10928 14076 10934 14088
rect 11333 14085 11345 14088
rect 11379 14085 11391 14119
rect 12452 14116 12480 14215
rect 13722 14116 13728 14128
rect 12452 14088 13728 14116
rect 11333 14079 11391 14085
rect 13722 14076 13728 14088
rect 13780 14076 13786 14128
rect 15764 14116 15792 14215
rect 17310 14116 17316 14128
rect 15764 14088 17316 14116
rect 17310 14076 17316 14088
rect 17368 14116 17374 14128
rect 18064 14116 18092 14215
rect 17368 14088 18092 14116
rect 17368 14076 17374 14088
rect 20622 14076 20628 14128
rect 20680 14116 20686 14128
rect 20717 14119 20775 14125
rect 20717 14116 20729 14119
rect 20680 14088 20729 14116
rect 20680 14076 20686 14088
rect 20717 14085 20729 14088
rect 20763 14085 20775 14119
rect 20717 14079 20775 14085
rect 1104 14026 21896 14048
rect 1104 13974 4447 14026
rect 4499 13974 4511 14026
rect 4563 13974 4575 14026
rect 4627 13974 4639 14026
rect 4691 13974 11378 14026
rect 11430 13974 11442 14026
rect 11494 13974 11506 14026
rect 11558 13974 11570 14026
rect 11622 13974 18308 14026
rect 18360 13974 18372 14026
rect 18424 13974 18436 14026
rect 18488 13974 18500 14026
rect 18552 13974 21896 14026
rect 1104 13952 21896 13974
rect 13078 13912 13084 13924
rect 13039 13884 13084 13912
rect 13078 13872 13084 13884
rect 13136 13872 13142 13924
rect 17313 13915 17371 13921
rect 13556 13884 13768 13912
rect 6917 13847 6975 13853
rect 6917 13813 6929 13847
rect 6963 13844 6975 13847
rect 8846 13844 8852 13856
rect 6963 13816 8852 13844
rect 6963 13813 6975 13816
rect 6917 13807 6975 13813
rect 8846 13804 8852 13816
rect 8904 13804 8910 13856
rect 10229 13847 10287 13853
rect 10229 13813 10241 13847
rect 10275 13844 10287 13847
rect 11330 13844 11336 13856
rect 10275 13816 11336 13844
rect 10275 13813 10287 13816
rect 10229 13807 10287 13813
rect 11330 13804 11336 13816
rect 11388 13804 11394 13856
rect 7466 13776 7472 13788
rect 7427 13748 7472 13776
rect 7466 13736 7472 13748
rect 7524 13736 7530 13788
rect 9674 13736 9680 13788
rect 9732 13776 9738 13788
rect 10689 13779 10747 13785
rect 10689 13776 10701 13779
rect 9732 13748 10701 13776
rect 9732 13736 9738 13748
rect 10689 13745 10701 13748
rect 10735 13745 10747 13779
rect 10870 13776 10876 13788
rect 10831 13748 10876 13776
rect 10689 13739 10747 13745
rect 10870 13736 10876 13748
rect 10928 13736 10934 13788
rect 7282 13708 7288 13720
rect 7243 13680 7288 13708
rect 7282 13668 7288 13680
rect 7340 13668 7346 13720
rect 11793 13711 11851 13717
rect 11793 13677 11805 13711
rect 11839 13708 11851 13711
rect 13556 13708 13584 13884
rect 13633 13847 13691 13853
rect 13633 13813 13645 13847
rect 13679 13813 13691 13847
rect 13740 13844 13768 13884
rect 17313 13881 17325 13915
rect 17359 13912 17371 13915
rect 17954 13912 17960 13924
rect 17359 13884 17960 13912
rect 17359 13881 17371 13884
rect 17313 13875 17371 13881
rect 17954 13872 17960 13884
rect 18012 13872 18018 13924
rect 18966 13844 18972 13856
rect 13740 13816 18972 13844
rect 13633 13807 13691 13813
rect 11839 13680 13584 13708
rect 13648 13708 13676 13807
rect 18966 13804 18972 13816
rect 19024 13804 19030 13856
rect 13906 13736 13912 13788
rect 13964 13776 13970 13788
rect 14093 13779 14151 13785
rect 14093 13776 14105 13779
rect 13964 13748 14105 13776
rect 13964 13736 13970 13748
rect 14093 13745 14105 13748
rect 14139 13745 14151 13779
rect 14093 13739 14151 13745
rect 14182 13736 14188 13788
rect 14240 13776 14246 13788
rect 16117 13779 16175 13785
rect 14240 13748 14285 13776
rect 14240 13736 14246 13748
rect 16117 13745 16129 13779
rect 16163 13776 16175 13779
rect 18877 13779 18935 13785
rect 16163 13748 18828 13776
rect 16163 13745 16175 13748
rect 16117 13739 16175 13745
rect 15841 13711 15899 13717
rect 15841 13708 15853 13711
rect 13648 13680 15853 13708
rect 11839 13677 11851 13680
rect 11793 13671 11851 13677
rect 15841 13677 15853 13680
rect 15887 13677 15899 13711
rect 15841 13671 15899 13677
rect 15930 13668 15936 13720
rect 15988 13708 15994 13720
rect 17129 13711 17187 13717
rect 17129 13708 17141 13711
rect 15988 13680 17141 13708
rect 15988 13668 15994 13680
rect 17129 13677 17141 13680
rect 17175 13677 17187 13711
rect 17129 13671 17187 13677
rect 17218 13668 17224 13720
rect 17276 13708 17282 13720
rect 18693 13711 18751 13717
rect 18693 13708 18705 13711
rect 17276 13680 18705 13708
rect 17276 13668 17282 13680
rect 18693 13677 18705 13680
rect 18739 13677 18751 13711
rect 18800 13708 18828 13748
rect 18877 13745 18889 13779
rect 18923 13776 18935 13779
rect 19150 13776 19156 13788
rect 18923 13748 19156 13776
rect 18923 13745 18935 13748
rect 18877 13739 18935 13745
rect 19150 13736 19156 13748
rect 19208 13736 19214 13788
rect 20530 13708 20536 13720
rect 18800 13680 20536 13708
rect 18693 13671 18751 13677
rect 20530 13668 20536 13680
rect 20588 13668 20594 13720
rect 7190 13600 7196 13652
rect 7248 13640 7254 13652
rect 11238 13640 11244 13652
rect 7248 13612 11244 13640
rect 7248 13600 7254 13612
rect 11238 13600 11244 13612
rect 11296 13640 11302 13652
rect 12342 13640 12348 13652
rect 11296 13612 12348 13640
rect 11296 13600 11302 13612
rect 12342 13600 12348 13612
rect 12400 13600 12406 13652
rect 14001 13643 14059 13649
rect 14001 13609 14013 13643
rect 14047 13640 14059 13643
rect 15286 13640 15292 13652
rect 14047 13612 15292 13640
rect 14047 13609 14059 13612
rect 14001 13603 14059 13609
rect 15286 13600 15292 13612
rect 15344 13600 15350 13652
rect 19242 13600 19248 13652
rect 19300 13640 19306 13652
rect 19797 13643 19855 13649
rect 19797 13640 19809 13643
rect 19300 13612 19809 13640
rect 19300 13600 19306 13612
rect 19797 13609 19809 13612
rect 19843 13609 19855 13643
rect 19797 13603 19855 13609
rect 7374 13572 7380 13584
rect 7335 13544 7380 13572
rect 7374 13532 7380 13544
rect 7432 13532 7438 13584
rect 10502 13532 10508 13584
rect 10560 13572 10566 13584
rect 10597 13575 10655 13581
rect 10597 13572 10609 13575
rect 10560 13544 10609 13572
rect 10560 13532 10566 13544
rect 10597 13541 10609 13544
rect 10643 13572 10655 13575
rect 16666 13572 16672 13584
rect 10643 13544 16672 13572
rect 10643 13541 10655 13544
rect 10597 13535 10655 13541
rect 16666 13532 16672 13544
rect 16724 13532 16730 13584
rect 18138 13532 18144 13584
rect 18196 13572 18202 13584
rect 18233 13575 18291 13581
rect 18233 13572 18245 13575
rect 18196 13544 18245 13572
rect 18196 13532 18202 13544
rect 18233 13541 18245 13544
rect 18279 13541 18291 13575
rect 18598 13572 18604 13584
rect 18559 13544 18604 13572
rect 18233 13535 18291 13541
rect 18598 13532 18604 13544
rect 18656 13532 18662 13584
rect 1104 13482 21896 13504
rect 1104 13430 7912 13482
rect 7964 13430 7976 13482
rect 8028 13430 8040 13482
rect 8092 13430 8104 13482
rect 8156 13430 14843 13482
rect 14895 13430 14907 13482
rect 14959 13430 14971 13482
rect 15023 13430 15035 13482
rect 15087 13430 21896 13482
rect 1104 13408 21896 13430
rect 7009 13371 7067 13377
rect 7009 13337 7021 13371
rect 7055 13368 7067 13371
rect 7374 13368 7380 13380
rect 7055 13340 7380 13368
rect 7055 13337 7067 13340
rect 7009 13331 7067 13337
rect 7374 13328 7380 13340
rect 7432 13328 7438 13380
rect 11330 13328 11336 13380
rect 11388 13368 11394 13380
rect 12897 13371 12955 13377
rect 12897 13368 12909 13371
rect 11388 13340 12909 13368
rect 11388 13328 11394 13340
rect 12897 13337 12909 13340
rect 12943 13337 12955 13371
rect 16301 13371 16359 13377
rect 12897 13331 12955 13337
rect 13004 13340 16059 13368
rect 5534 13260 5540 13312
rect 5592 13300 5598 13312
rect 7469 13303 7527 13309
rect 7469 13300 7481 13303
rect 5592 13272 7481 13300
rect 5592 13260 5598 13272
rect 7469 13269 7481 13272
rect 7515 13269 7527 13303
rect 7469 13263 7527 13269
rect 10404 13303 10462 13309
rect 10404 13269 10416 13303
rect 10450 13300 10462 13303
rect 10870 13300 10876 13312
rect 10450 13272 10876 13300
rect 10450 13269 10462 13272
rect 10404 13263 10462 13269
rect 10870 13260 10876 13272
rect 10928 13260 10934 13312
rect 13004 13300 13032 13340
rect 12728 13272 13032 13300
rect 14645 13303 14703 13309
rect 7190 13192 7196 13244
rect 7248 13232 7254 13244
rect 7377 13235 7435 13241
rect 7377 13232 7389 13235
rect 7248 13204 7389 13232
rect 7248 13192 7254 13204
rect 7377 13201 7389 13204
rect 7423 13201 7435 13235
rect 8846 13232 8852 13244
rect 8807 13204 8852 13232
rect 7377 13195 7435 13201
rect 8846 13192 8852 13204
rect 8904 13192 8910 13244
rect 9398 13192 9404 13244
rect 9456 13192 9462 13244
rect 9582 13192 9588 13244
rect 9640 13232 9646 13244
rect 12728 13232 12756 13272
rect 14645 13269 14657 13303
rect 14691 13300 14703 13303
rect 15930 13300 15936 13312
rect 14691 13272 15936 13300
rect 14691 13269 14703 13272
rect 14645 13263 14703 13269
rect 15930 13260 15936 13272
rect 15988 13260 15994 13312
rect 16031 13300 16059 13340
rect 16301 13337 16313 13371
rect 16347 13368 16359 13371
rect 17218 13368 17224 13380
rect 16347 13340 17224 13368
rect 16347 13337 16359 13340
rect 16301 13331 16359 13337
rect 17218 13328 17224 13340
rect 17276 13328 17282 13380
rect 18690 13328 18696 13380
rect 18748 13368 18754 13380
rect 18966 13368 18972 13380
rect 18748 13340 18972 13368
rect 18748 13328 18754 13340
rect 18966 13328 18972 13340
rect 19024 13368 19030 13380
rect 19061 13371 19119 13377
rect 19061 13368 19073 13371
rect 19024 13340 19073 13368
rect 19024 13328 19030 13340
rect 19061 13337 19073 13340
rect 19107 13337 19119 13371
rect 19061 13331 19119 13337
rect 17402 13300 17408 13312
rect 16031 13272 17408 13300
rect 17402 13260 17408 13272
rect 17460 13260 17466 13312
rect 20438 13300 20444 13312
rect 20399 13272 20444 13300
rect 20438 13260 20444 13272
rect 20496 13260 20502 13312
rect 9640 13204 12756 13232
rect 12805 13235 12863 13241
rect 9640 13192 9646 13204
rect 12805 13201 12817 13235
rect 12851 13232 12863 13235
rect 13170 13232 13176 13244
rect 12851 13204 13176 13232
rect 12851 13201 12863 13204
rect 12805 13195 12863 13201
rect 13170 13192 13176 13204
rect 13228 13192 13234 13244
rect 13906 13192 13912 13244
rect 13964 13232 13970 13244
rect 14369 13235 14427 13241
rect 14369 13232 14381 13235
rect 13964 13204 14381 13232
rect 13964 13192 13970 13204
rect 14369 13201 14381 13204
rect 14415 13201 14427 13235
rect 14369 13195 14427 13201
rect 15378 13192 15384 13244
rect 15436 13232 15442 13244
rect 16117 13235 16175 13241
rect 16117 13232 16129 13235
rect 15436 13204 16129 13232
rect 15436 13192 15442 13204
rect 16117 13201 16129 13204
rect 16163 13201 16175 13235
rect 16666 13232 16672 13244
rect 16579 13204 16672 13232
rect 16117 13195 16175 13201
rect 7650 13164 7656 13176
rect 7611 13136 7656 13164
rect 7650 13124 7656 13136
rect 7708 13124 7714 13176
rect 9125 13167 9183 13173
rect 9125 13133 9137 13167
rect 9171 13164 9183 13167
rect 9416 13164 9444 13192
rect 10137 13167 10195 13173
rect 10137 13164 10149 13167
rect 9171 13136 9444 13164
rect 9600 13136 10149 13164
rect 9171 13133 9183 13136
rect 9125 13127 9183 13133
rect 9600 13108 9628 13136
rect 10137 13133 10149 13136
rect 10183 13133 10195 13167
rect 11790 13164 11796 13176
rect 10137 13127 10195 13133
rect 11532 13136 11796 13164
rect 9582 13056 9588 13108
rect 9640 13056 9646 13108
rect 11532 13105 11560 13136
rect 11790 13124 11796 13136
rect 11848 13164 11854 13176
rect 13078 13164 13084 13176
rect 11848 13136 13084 13164
rect 11848 13124 11854 13136
rect 13078 13124 13084 13136
rect 13136 13124 13142 13176
rect 16132 13164 16160 13195
rect 16666 13192 16672 13204
rect 16724 13232 16730 13244
rect 16724 13204 17080 13232
rect 16724 13192 16730 13204
rect 16761 13167 16819 13173
rect 16761 13164 16773 13167
rect 16132 13136 16773 13164
rect 16761 13133 16773 13136
rect 16807 13133 16819 13167
rect 16942 13164 16948 13176
rect 16903 13136 16948 13164
rect 16761 13127 16819 13133
rect 16942 13124 16948 13136
rect 17000 13124 17006 13176
rect 17052 13164 17080 13204
rect 17954 13192 17960 13244
rect 18012 13232 18018 13244
rect 18969 13235 19027 13241
rect 18969 13232 18981 13235
rect 18012 13204 18981 13232
rect 18012 13192 18018 13204
rect 18969 13201 18981 13204
rect 19015 13201 19027 13235
rect 20162 13232 20168 13244
rect 20123 13204 20168 13232
rect 18969 13195 19027 13201
rect 20162 13192 20168 13204
rect 20220 13192 20226 13244
rect 18874 13164 18880 13176
rect 17052 13136 18880 13164
rect 18874 13124 18880 13136
rect 18932 13124 18938 13176
rect 19150 13164 19156 13176
rect 19111 13136 19156 13164
rect 19150 13124 19156 13136
rect 19208 13124 19214 13176
rect 11517 13099 11575 13105
rect 11517 13065 11529 13099
rect 11563 13065 11575 13099
rect 11517 13059 11575 13065
rect 15746 13056 15752 13108
rect 15804 13096 15810 13108
rect 21542 13096 21548 13108
rect 15804 13068 21548 13096
rect 15804 13056 15810 13068
rect 21542 13056 21548 13068
rect 21600 13056 21606 13108
rect 12437 13031 12495 13037
rect 12437 12997 12449 13031
rect 12483 13028 12495 13031
rect 12986 13028 12992 13040
rect 12483 13000 12992 13028
rect 12483 12997 12495 13000
rect 12437 12991 12495 12997
rect 12986 12988 12992 13000
rect 13044 12988 13050 13040
rect 18601 13031 18659 13037
rect 18601 12997 18613 13031
rect 18647 13028 18659 13031
rect 19242 13028 19248 13040
rect 18647 13000 19248 13028
rect 18647 12997 18659 13000
rect 18601 12991 18659 12997
rect 19242 12988 19248 13000
rect 19300 12988 19306 13040
rect 1104 12938 21896 12960
rect 1104 12886 4447 12938
rect 4499 12886 4511 12938
rect 4563 12886 4575 12938
rect 4627 12886 4639 12938
rect 4691 12886 11378 12938
rect 11430 12886 11442 12938
rect 11494 12886 11506 12938
rect 11558 12886 11570 12938
rect 11622 12886 18308 12938
rect 18360 12886 18372 12938
rect 18424 12886 18436 12938
rect 18488 12886 18500 12938
rect 18552 12886 21896 12938
rect 1104 12864 21896 12886
rect 7377 12827 7435 12833
rect 7377 12793 7389 12827
rect 7423 12824 7435 12827
rect 7466 12824 7472 12836
rect 7423 12796 7472 12824
rect 7423 12793 7435 12796
rect 7377 12787 7435 12793
rect 7466 12784 7472 12796
rect 7524 12784 7530 12836
rect 18877 12827 18935 12833
rect 18877 12793 18889 12827
rect 18923 12824 18935 12827
rect 20162 12824 20168 12836
rect 18923 12796 20168 12824
rect 18923 12793 18935 12796
rect 18877 12787 18935 12793
rect 20162 12784 20168 12796
rect 20220 12784 20226 12836
rect 15746 12756 15752 12768
rect 15707 12728 15752 12756
rect 15746 12716 15752 12728
rect 15804 12716 15810 12768
rect 18049 12759 18107 12765
rect 18049 12725 18061 12759
rect 18095 12756 18107 12759
rect 19150 12756 19156 12768
rect 18095 12728 19156 12756
rect 18095 12725 18107 12728
rect 18049 12719 18107 12725
rect 19150 12716 19156 12728
rect 19208 12716 19214 12768
rect 13078 12648 13084 12700
rect 13136 12688 13142 12700
rect 14001 12691 14059 12697
rect 14001 12688 14013 12691
rect 13136 12660 14013 12688
rect 13136 12648 13142 12660
rect 14001 12657 14013 12660
rect 14047 12657 14059 12691
rect 14001 12651 14059 12657
rect 15212 12660 16804 12688
rect 5994 12620 6000 12632
rect 5955 12592 6000 12620
rect 5994 12580 6000 12592
rect 6052 12580 6058 12632
rect 6264 12623 6322 12629
rect 6264 12589 6276 12623
rect 6310 12620 6322 12623
rect 7650 12620 7656 12632
rect 6310 12592 7656 12620
rect 6310 12589 6322 12592
rect 6264 12583 6322 12589
rect 7650 12580 7656 12592
rect 7708 12580 7714 12632
rect 11241 12623 11299 12629
rect 11241 12589 11253 12623
rect 11287 12589 11299 12623
rect 11241 12583 11299 12589
rect 11508 12623 11566 12629
rect 11508 12589 11520 12623
rect 11554 12620 11566 12623
rect 11790 12620 11796 12632
rect 11554 12592 11796 12620
rect 11554 12589 11566 12592
rect 11508 12583 11566 12589
rect 8662 12512 8668 12564
rect 8720 12552 8726 12564
rect 9398 12552 9404 12564
rect 8720 12524 9404 12552
rect 8720 12512 8726 12524
rect 9398 12512 9404 12524
rect 9456 12552 9462 12564
rect 11256 12552 11284 12583
rect 11790 12580 11796 12592
rect 11848 12580 11854 12632
rect 13909 12623 13967 12629
rect 13909 12589 13921 12623
rect 13955 12620 13967 12623
rect 15212 12620 15240 12660
rect 13955 12592 15240 12620
rect 15565 12623 15623 12629
rect 13955 12589 13967 12592
rect 13909 12583 13967 12589
rect 15565 12589 15577 12623
rect 15611 12589 15623 12623
rect 16666 12620 16672 12632
rect 16627 12592 16672 12620
rect 15565 12583 15623 12589
rect 9456 12524 11284 12552
rect 9456 12512 9462 12524
rect 13170 12512 13176 12564
rect 13228 12552 13234 12564
rect 15580 12552 15608 12583
rect 16666 12580 16672 12592
rect 16724 12580 16730 12632
rect 16776 12620 16804 12660
rect 18138 12648 18144 12700
rect 18196 12688 18202 12700
rect 19337 12691 19395 12697
rect 19337 12688 19349 12691
rect 18196 12660 19349 12688
rect 18196 12648 18202 12660
rect 19337 12657 19349 12660
rect 19383 12657 19395 12691
rect 19337 12651 19395 12657
rect 19429 12691 19487 12697
rect 19429 12657 19441 12691
rect 19475 12657 19487 12691
rect 19429 12651 19487 12657
rect 18966 12620 18972 12632
rect 16776 12592 18972 12620
rect 18966 12580 18972 12592
rect 19024 12580 19030 12632
rect 19242 12620 19248 12632
rect 19203 12592 19248 12620
rect 19242 12580 19248 12592
rect 19300 12580 19306 12632
rect 19444 12620 19472 12651
rect 19352 12592 19472 12620
rect 16574 12552 16580 12564
rect 13228 12524 14044 12552
rect 15580 12524 16580 12552
rect 13228 12512 13234 12524
rect 12618 12484 12624 12496
rect 12579 12456 12624 12484
rect 12618 12444 12624 12456
rect 12676 12444 12682 12496
rect 13446 12484 13452 12496
rect 13407 12456 13452 12484
rect 13446 12444 13452 12456
rect 13504 12444 13510 12496
rect 13814 12484 13820 12496
rect 13775 12456 13820 12484
rect 13814 12444 13820 12456
rect 13872 12444 13878 12496
rect 14016 12484 14044 12524
rect 16574 12512 16580 12524
rect 16632 12512 16638 12564
rect 16942 12561 16948 12564
rect 16936 12552 16948 12561
rect 16903 12524 16948 12552
rect 16936 12515 16948 12524
rect 16942 12512 16948 12515
rect 17000 12512 17006 12564
rect 19058 12512 19064 12564
rect 19116 12552 19122 12564
rect 19352 12552 19380 12592
rect 19116 12524 19380 12552
rect 19116 12512 19122 12524
rect 18598 12484 18604 12496
rect 14016 12456 18604 12484
rect 18598 12444 18604 12456
rect 18656 12444 18662 12496
rect 1104 12394 21896 12416
rect 1104 12342 7912 12394
rect 7964 12342 7976 12394
rect 8028 12342 8040 12394
rect 8092 12342 8104 12394
rect 8156 12342 14843 12394
rect 14895 12342 14907 12394
rect 14959 12342 14971 12394
rect 15023 12342 15035 12394
rect 15087 12342 21896 12394
rect 1104 12320 21896 12342
rect 7282 12280 7288 12292
rect 7243 12252 7288 12280
rect 7282 12240 7288 12252
rect 7340 12240 7346 12292
rect 7650 12240 7656 12292
rect 7708 12280 7714 12292
rect 10045 12283 10103 12289
rect 10045 12280 10057 12283
rect 7708 12252 10057 12280
rect 7708 12240 7714 12252
rect 10045 12249 10057 12252
rect 10091 12249 10103 12283
rect 13078 12280 13084 12292
rect 13039 12252 13084 12280
rect 10045 12243 10103 12249
rect 13078 12240 13084 12252
rect 13136 12240 13142 12292
rect 16853 12283 16911 12289
rect 16853 12249 16865 12283
rect 16899 12280 16911 12283
rect 16942 12280 16948 12292
rect 16899 12252 16948 12280
rect 16899 12249 16911 12252
rect 16853 12243 16911 12249
rect 16942 12240 16948 12252
rect 17000 12240 17006 12292
rect 18046 12240 18052 12292
rect 18104 12280 18110 12292
rect 18509 12283 18567 12289
rect 18509 12280 18521 12283
rect 18104 12252 18521 12280
rect 18104 12240 18110 12252
rect 18509 12249 18521 12252
rect 18555 12249 18567 12283
rect 19610 12280 19616 12292
rect 19571 12252 19616 12280
rect 18509 12243 18567 12249
rect 19610 12240 19616 12252
rect 19668 12240 19674 12292
rect 20714 12280 20720 12292
rect 20675 12252 20720 12280
rect 20714 12240 20720 12252
rect 20772 12240 20778 12292
rect 8932 12215 8990 12221
rect 8932 12181 8944 12215
rect 8978 12212 8990 12215
rect 12618 12212 12624 12224
rect 8978 12184 12624 12212
rect 8978 12181 8990 12184
rect 8932 12175 8990 12181
rect 5994 12104 6000 12156
rect 6052 12144 6058 12156
rect 8662 12144 8668 12156
rect 6052 12116 8668 12144
rect 6052 12104 6058 12116
rect 8662 12104 8668 12116
rect 8720 12104 8726 12156
rect 12452 12144 12480 12184
rect 12618 12172 12624 12184
rect 12676 12172 12682 12224
rect 12989 12215 13047 12221
rect 12989 12181 13001 12215
rect 13035 12212 13047 12215
rect 13446 12212 13452 12224
rect 13035 12184 13452 12212
rect 13035 12181 13047 12184
rect 12989 12175 13047 12181
rect 13446 12172 13452 12184
rect 13504 12172 13510 12224
rect 18414 12212 18420 12224
rect 14384 12184 18420 12212
rect 14384 12153 14412 12184
rect 18414 12172 18420 12184
rect 18472 12172 18478 12224
rect 15746 12153 15752 12156
rect 14369 12147 14427 12153
rect 12452 12116 13308 12144
rect 13280 12085 13308 12116
rect 14369 12113 14381 12147
rect 14415 12113 14427 12147
rect 14369 12107 14427 12113
rect 15740 12107 15752 12153
rect 15804 12144 15810 12156
rect 15804 12116 15840 12144
rect 15746 12104 15752 12107
rect 15804 12104 15810 12116
rect 18138 12104 18144 12156
rect 18196 12144 18202 12156
rect 18325 12147 18383 12153
rect 18325 12144 18337 12147
rect 18196 12116 18337 12144
rect 18196 12104 18202 12116
rect 18325 12113 18337 12116
rect 18371 12113 18383 12147
rect 18325 12107 18383 12113
rect 19429 12147 19487 12153
rect 19429 12113 19441 12147
rect 19475 12144 19487 12147
rect 19702 12144 19708 12156
rect 19475 12116 19708 12144
rect 19475 12113 19487 12116
rect 19429 12107 19487 12113
rect 19702 12104 19708 12116
rect 19760 12104 19766 12156
rect 20530 12144 20536 12156
rect 20491 12116 20536 12144
rect 20530 12104 20536 12116
rect 20588 12104 20594 12156
rect 13265 12079 13323 12085
rect 13265 12045 13277 12079
rect 13311 12045 13323 12079
rect 13265 12039 13323 12045
rect 13722 12036 13728 12088
rect 13780 12076 13786 12088
rect 15473 12079 15531 12085
rect 15473 12076 15485 12079
rect 13780 12048 15485 12076
rect 13780 12036 13786 12048
rect 15473 12045 15485 12048
rect 15519 12045 15531 12079
rect 15473 12039 15531 12045
rect 16574 11968 16580 12020
rect 16632 12008 16638 12020
rect 18690 12008 18696 12020
rect 16632 11980 18696 12008
rect 16632 11968 16638 11980
rect 18690 11968 18696 11980
rect 18748 11968 18754 12020
rect 12621 11943 12679 11949
rect 12621 11909 12633 11943
rect 12667 11940 12679 11943
rect 13906 11940 13912 11952
rect 12667 11912 13912 11940
rect 12667 11909 12679 11912
rect 12621 11903 12679 11909
rect 13906 11900 13912 11912
rect 13964 11900 13970 11952
rect 14553 11943 14611 11949
rect 14553 11909 14565 11943
rect 14599 11940 14611 11943
rect 20990 11940 20996 11952
rect 14599 11912 20996 11940
rect 14599 11909 14611 11912
rect 14553 11903 14611 11909
rect 20990 11900 20996 11912
rect 21048 11900 21054 11952
rect 1104 11850 21896 11872
rect 1104 11798 4447 11850
rect 4499 11798 4511 11850
rect 4563 11798 4575 11850
rect 4627 11798 4639 11850
rect 4691 11798 11378 11850
rect 11430 11798 11442 11850
rect 11494 11798 11506 11850
rect 11558 11798 11570 11850
rect 11622 11798 18308 11850
rect 18360 11798 18372 11850
rect 18424 11798 18436 11850
rect 18488 11798 18500 11850
rect 18552 11798 21896 11850
rect 1104 11776 21896 11798
rect 15289 11671 15347 11677
rect 15289 11637 15301 11671
rect 15335 11668 15347 11671
rect 15335 11640 19564 11668
rect 15335 11637 15347 11640
rect 15289 11631 15347 11637
rect 13633 11603 13691 11609
rect 13633 11569 13645 11603
rect 13679 11600 13691 11603
rect 13814 11600 13820 11612
rect 13679 11572 13820 11600
rect 13679 11569 13691 11572
rect 13633 11563 13691 11569
rect 13814 11560 13820 11572
rect 13872 11560 13878 11612
rect 15746 11560 15752 11612
rect 15804 11600 15810 11612
rect 15841 11603 15899 11609
rect 15841 11600 15853 11603
rect 15804 11572 15853 11600
rect 15804 11560 15810 11572
rect 15841 11569 15853 11572
rect 15887 11569 15899 11603
rect 15841 11563 15899 11569
rect 16853 11603 16911 11609
rect 16853 11569 16865 11603
rect 16899 11600 16911 11603
rect 17954 11600 17960 11612
rect 16899 11572 17960 11600
rect 16899 11569 16911 11572
rect 16853 11563 16911 11569
rect 17954 11560 17960 11572
rect 18012 11560 18018 11612
rect 18138 11600 18144 11612
rect 18099 11572 18144 11600
rect 18138 11560 18144 11572
rect 18196 11560 18202 11612
rect 12529 11535 12587 11541
rect 12529 11501 12541 11535
rect 12575 11532 12587 11535
rect 12894 11532 12900 11544
rect 12575 11504 12900 11532
rect 12575 11501 12587 11504
rect 12529 11495 12587 11501
rect 12894 11492 12900 11504
rect 12952 11492 12958 11544
rect 17865 11535 17923 11541
rect 17865 11501 17877 11535
rect 17911 11532 17923 11535
rect 18046 11532 18052 11544
rect 17911 11504 18052 11532
rect 17911 11501 17923 11504
rect 17865 11495 17923 11501
rect 18046 11492 18052 11504
rect 18104 11492 18110 11544
rect 19536 11541 19564 11640
rect 19702 11600 19708 11612
rect 19663 11572 19708 11600
rect 19702 11560 19708 11572
rect 19760 11560 19766 11612
rect 19521 11535 19579 11541
rect 19521 11501 19533 11535
rect 19567 11501 19579 11535
rect 19521 11495 19579 11501
rect 15378 11424 15384 11476
rect 15436 11464 15442 11476
rect 15749 11467 15807 11473
rect 15749 11464 15761 11467
rect 15436 11436 15761 11464
rect 15436 11424 15442 11436
rect 15749 11433 15761 11436
rect 15795 11433 15807 11467
rect 15749 11427 15807 11433
rect 11790 11356 11796 11408
rect 11848 11396 11854 11408
rect 12345 11399 12403 11405
rect 12345 11396 12357 11399
rect 11848 11368 12357 11396
rect 11848 11356 11854 11368
rect 12345 11365 12357 11368
rect 12391 11365 12403 11399
rect 15654 11396 15660 11408
rect 15615 11368 15660 11396
rect 12345 11359 12403 11365
rect 15654 11356 15660 11368
rect 15712 11356 15718 11408
rect 1104 11306 21896 11328
rect 1104 11254 7912 11306
rect 7964 11254 7976 11306
rect 8028 11254 8040 11306
rect 8092 11254 8104 11306
rect 8156 11254 14843 11306
rect 14895 11254 14907 11306
rect 14959 11254 14971 11306
rect 15023 11254 15035 11306
rect 15087 11254 21896 11306
rect 1104 11232 21896 11254
rect 12802 11152 12808 11204
rect 12860 11192 12866 11204
rect 12989 11195 13047 11201
rect 12989 11192 13001 11195
rect 12860 11164 13001 11192
rect 12860 11152 12866 11164
rect 12989 11161 13001 11164
rect 13035 11161 13047 11195
rect 12989 11155 13047 11161
rect 13078 11152 13084 11204
rect 13136 11192 13142 11204
rect 15746 11192 15752 11204
rect 13136 11164 14504 11192
rect 15707 11164 15752 11192
rect 13136 11152 13142 11164
rect 11790 11084 11796 11136
rect 11848 11124 11854 11136
rect 14476 11124 14504 11164
rect 15746 11152 15752 11164
rect 15804 11152 15810 11204
rect 17037 11195 17095 11201
rect 17037 11161 17049 11195
rect 17083 11192 17095 11195
rect 17770 11192 17776 11204
rect 17083 11164 17776 11192
rect 17083 11161 17095 11164
rect 17037 11155 17095 11161
rect 17770 11152 17776 11164
rect 17828 11152 17834 11204
rect 18046 11192 18052 11204
rect 18007 11164 18052 11192
rect 18046 11152 18052 11164
rect 18104 11152 18110 11204
rect 20346 11152 20352 11204
rect 20404 11192 20410 11204
rect 20533 11195 20591 11201
rect 20533 11192 20545 11195
rect 20404 11164 20545 11192
rect 20404 11152 20410 11164
rect 20533 11161 20545 11164
rect 20579 11161 20591 11195
rect 20533 11155 20591 11161
rect 18966 11124 18972 11136
rect 11848 11096 14320 11124
rect 14476 11096 18972 11124
rect 11848 11084 11854 11096
rect 12434 11016 12440 11068
rect 12492 11056 12498 11068
rect 12897 11059 12955 11065
rect 12897 11056 12909 11059
rect 12492 11028 12909 11056
rect 12492 11016 12498 11028
rect 12897 11025 12909 11028
rect 12943 11056 12955 11059
rect 13078 11056 13084 11068
rect 12943 11028 13084 11056
rect 12943 11025 12955 11028
rect 12897 11019 12955 11025
rect 13078 11016 13084 11028
rect 13136 11016 13142 11068
rect 14292 11065 14320 11096
rect 18966 11084 18972 11096
rect 19024 11084 19030 11136
rect 14277 11059 14335 11065
rect 14277 11025 14289 11059
rect 14323 11025 14335 11059
rect 14277 11019 14335 11025
rect 14458 11016 14464 11068
rect 14516 11056 14522 11068
rect 14625 11059 14683 11065
rect 14625 11056 14637 11059
rect 14516 11028 14637 11056
rect 14516 11016 14522 11028
rect 14625 11025 14637 11028
rect 14671 11025 14683 11059
rect 14625 11019 14683 11025
rect 16853 11059 16911 11065
rect 16853 11025 16865 11059
rect 16899 11056 16911 11059
rect 17954 11056 17960 11068
rect 16899 11028 17960 11056
rect 16899 11025 16911 11028
rect 16853 11019 16911 11025
rect 17954 11016 17960 11028
rect 18012 11016 18018 11068
rect 18138 11016 18144 11068
rect 18196 11056 18202 11068
rect 18417 11059 18475 11065
rect 18417 11056 18429 11059
rect 18196 11028 18429 11056
rect 18196 11016 18202 11028
rect 18417 11025 18429 11028
rect 18463 11025 18475 11059
rect 20346 11056 20352 11068
rect 20307 11028 20352 11056
rect 18417 11019 18475 11025
rect 20346 11016 20352 11028
rect 20404 11016 20410 11068
rect 13170 10988 13176 11000
rect 13131 10960 13176 10988
rect 13170 10948 13176 10960
rect 13228 10948 13234 11000
rect 14369 10991 14427 10997
rect 14369 10988 14381 10991
rect 14292 10960 14381 10988
rect 12529 10923 12587 10929
rect 12529 10889 12541 10923
rect 12575 10920 12587 10923
rect 14182 10920 14188 10932
rect 12575 10892 14188 10920
rect 12575 10889 12587 10892
rect 12529 10883 12587 10889
rect 14182 10880 14188 10892
rect 14240 10880 14246 10932
rect 12802 10812 12808 10864
rect 12860 10852 12866 10864
rect 13722 10852 13728 10864
rect 12860 10824 13728 10852
rect 12860 10812 12866 10824
rect 13722 10812 13728 10824
rect 13780 10852 13786 10864
rect 14093 10855 14151 10861
rect 14093 10852 14105 10855
rect 13780 10824 14105 10852
rect 13780 10812 13786 10824
rect 14093 10821 14105 10824
rect 14139 10852 14151 10855
rect 14292 10852 14320 10960
rect 14369 10957 14381 10960
rect 14415 10957 14427 10991
rect 14369 10951 14427 10957
rect 18046 10948 18052 11000
rect 18104 10988 18110 11000
rect 18509 10991 18567 10997
rect 18509 10988 18521 10991
rect 18104 10960 18521 10988
rect 18104 10948 18110 10960
rect 18509 10957 18521 10960
rect 18555 10957 18567 10991
rect 18690 10988 18696 11000
rect 18651 10960 18696 10988
rect 18509 10951 18567 10957
rect 18690 10948 18696 10960
rect 18748 10948 18754 11000
rect 14139 10824 14320 10852
rect 14139 10821 14151 10824
rect 14093 10815 14151 10821
rect 1104 10762 21896 10784
rect 1104 10710 4447 10762
rect 4499 10710 4511 10762
rect 4563 10710 4575 10762
rect 4627 10710 4639 10762
rect 4691 10710 11378 10762
rect 11430 10710 11442 10762
rect 11494 10710 11506 10762
rect 11558 10710 11570 10762
rect 11622 10710 18308 10762
rect 18360 10710 18372 10762
rect 18424 10710 18436 10762
rect 18488 10710 18500 10762
rect 18552 10710 21896 10762
rect 1104 10688 21896 10710
rect 13170 10608 13176 10660
rect 13228 10648 13234 10660
rect 13265 10651 13323 10657
rect 13265 10648 13277 10651
rect 13228 10620 13277 10648
rect 13228 10608 13234 10620
rect 13265 10617 13277 10620
rect 13311 10617 13323 10651
rect 13265 10611 13323 10617
rect 15289 10651 15347 10657
rect 15289 10617 15301 10651
rect 15335 10648 15347 10651
rect 15378 10648 15384 10660
rect 15335 10620 15384 10648
rect 15335 10617 15347 10620
rect 15289 10611 15347 10617
rect 15378 10608 15384 10620
rect 15436 10608 15442 10660
rect 19886 10648 19892 10660
rect 19847 10620 19892 10648
rect 19886 10608 19892 10620
rect 19944 10608 19950 10660
rect 14458 10540 14464 10592
rect 14516 10580 14522 10592
rect 14516 10552 15884 10580
rect 14516 10540 14522 10552
rect 14182 10472 14188 10524
rect 14240 10512 14246 10524
rect 15856 10521 15884 10552
rect 15749 10515 15807 10521
rect 15749 10512 15761 10515
rect 14240 10484 15761 10512
rect 14240 10472 14246 10484
rect 15749 10481 15761 10484
rect 15795 10481 15807 10515
rect 15749 10475 15807 10481
rect 15841 10515 15899 10521
rect 15841 10481 15853 10515
rect 15887 10481 15899 10515
rect 15841 10475 15899 10481
rect 10597 10447 10655 10453
rect 10597 10413 10609 10447
rect 10643 10444 10655 10447
rect 11790 10444 11796 10456
rect 10643 10416 11796 10444
rect 10643 10413 10655 10416
rect 10597 10407 10655 10413
rect 11790 10404 11796 10416
rect 11848 10404 11854 10456
rect 11885 10447 11943 10453
rect 11885 10413 11897 10447
rect 11931 10413 11943 10447
rect 11885 10407 11943 10413
rect 9398 10336 9404 10388
rect 9456 10376 9462 10388
rect 11900 10376 11928 10407
rect 16666 10404 16672 10456
rect 16724 10444 16730 10456
rect 17313 10447 17371 10453
rect 17313 10444 17325 10447
rect 16724 10416 17325 10444
rect 16724 10404 16730 10416
rect 17313 10413 17325 10416
rect 17359 10413 17371 10447
rect 17313 10407 17371 10413
rect 19242 10404 19248 10456
rect 19300 10444 19306 10456
rect 19705 10447 19763 10453
rect 19705 10444 19717 10447
rect 19300 10416 19717 10444
rect 19300 10404 19306 10416
rect 19705 10413 19717 10416
rect 19751 10413 19763 10447
rect 19705 10407 19763 10413
rect 9456 10348 11928 10376
rect 12152 10379 12210 10385
rect 9456 10336 9462 10348
rect 10428 10320 10456 10348
rect 12152 10345 12164 10379
rect 12198 10376 12210 10379
rect 17580 10379 17638 10385
rect 12198 10348 16620 10376
rect 12198 10345 12210 10348
rect 12152 10339 12210 10345
rect 10410 10308 10416 10320
rect 10371 10280 10416 10308
rect 10410 10268 10416 10280
rect 10468 10268 10474 10320
rect 14182 10308 14188 10320
rect 14143 10280 14188 10308
rect 14182 10268 14188 10280
rect 14240 10268 14246 10320
rect 15194 10268 15200 10320
rect 15252 10308 15258 10320
rect 15657 10311 15715 10317
rect 15657 10308 15669 10311
rect 15252 10280 15669 10308
rect 15252 10268 15258 10280
rect 15657 10277 15669 10280
rect 15703 10308 15715 10311
rect 15930 10308 15936 10320
rect 15703 10280 15936 10308
rect 15703 10277 15715 10280
rect 15657 10271 15715 10277
rect 15930 10268 15936 10280
rect 15988 10268 15994 10320
rect 16592 10308 16620 10348
rect 17580 10345 17592 10379
rect 17626 10376 17638 10379
rect 17954 10376 17960 10388
rect 17626 10348 17960 10376
rect 17626 10345 17638 10348
rect 17580 10339 17638 10345
rect 17954 10336 17960 10348
rect 18012 10336 18018 10388
rect 18690 10308 18696 10320
rect 16592 10280 18696 10308
rect 18690 10268 18696 10280
rect 18748 10268 18754 10320
rect 1104 10218 21896 10240
rect 1104 10166 7912 10218
rect 7964 10166 7976 10218
rect 8028 10166 8040 10218
rect 8092 10166 8104 10218
rect 8156 10166 14843 10218
rect 14895 10166 14907 10218
rect 14959 10166 14971 10218
rect 15023 10166 15035 10218
rect 15087 10166 21896 10218
rect 1104 10144 21896 10166
rect 14182 10064 14188 10116
rect 14240 10104 14246 10116
rect 15657 10107 15715 10113
rect 15657 10104 15669 10107
rect 14240 10076 15669 10104
rect 14240 10064 14246 10076
rect 15657 10073 15669 10076
rect 15703 10073 15715 10107
rect 18046 10104 18052 10116
rect 18007 10076 18052 10104
rect 15657 10067 15715 10073
rect 18046 10064 18052 10076
rect 18104 10064 18110 10116
rect 20717 10107 20775 10113
rect 20717 10073 20729 10107
rect 20763 10104 20775 10107
rect 21358 10104 21364 10116
rect 20763 10076 21364 10104
rect 20763 10073 20775 10076
rect 20717 10067 20775 10073
rect 21358 10064 21364 10076
rect 21416 10064 21422 10116
rect 13170 9996 13176 10048
rect 13228 10045 13234 10048
rect 13228 10039 13292 10045
rect 13228 10005 13246 10039
rect 13280 10005 13292 10039
rect 13228 9999 13292 10005
rect 13228 9996 13234 9999
rect 14458 9928 14464 9980
rect 14516 9968 14522 9980
rect 18417 9971 18475 9977
rect 14516 9940 15884 9968
rect 14516 9928 14522 9940
rect 12802 9860 12808 9912
rect 12860 9900 12866 9912
rect 12989 9903 13047 9909
rect 12989 9900 13001 9903
rect 12860 9872 13001 9900
rect 12860 9860 12866 9872
rect 12989 9869 13001 9872
rect 13035 9869 13047 9903
rect 15746 9900 15752 9912
rect 15707 9872 15752 9900
rect 12989 9863 13047 9869
rect 15746 9860 15752 9872
rect 15804 9860 15810 9912
rect 15856 9909 15884 9940
rect 18417 9937 18429 9971
rect 18463 9968 18475 9971
rect 18874 9968 18880 9980
rect 18463 9940 18880 9968
rect 18463 9937 18475 9940
rect 18417 9931 18475 9937
rect 18874 9928 18880 9940
rect 18932 9928 18938 9980
rect 20530 9968 20536 9980
rect 20491 9940 20536 9968
rect 20530 9928 20536 9940
rect 20588 9928 20594 9980
rect 15841 9903 15899 9909
rect 15841 9869 15853 9903
rect 15887 9869 15899 9903
rect 15841 9863 15899 9869
rect 18046 9860 18052 9912
rect 18104 9900 18110 9912
rect 18509 9903 18567 9909
rect 18509 9900 18521 9903
rect 18104 9872 18521 9900
rect 18104 9860 18110 9872
rect 18509 9869 18521 9872
rect 18555 9869 18567 9903
rect 18509 9863 18567 9869
rect 18601 9903 18659 9909
rect 18601 9869 18613 9903
rect 18647 9869 18659 9903
rect 18601 9863 18659 9869
rect 14369 9835 14427 9841
rect 14369 9801 14381 9835
rect 14415 9832 14427 9835
rect 14458 9832 14464 9844
rect 14415 9804 14464 9832
rect 14415 9801 14427 9804
rect 14369 9795 14427 9801
rect 14458 9792 14464 9804
rect 14516 9792 14522 9844
rect 15289 9835 15347 9841
rect 15289 9801 15301 9835
rect 15335 9832 15347 9835
rect 15654 9832 15660 9844
rect 15335 9804 15660 9832
rect 15335 9801 15347 9804
rect 15289 9795 15347 9801
rect 15654 9792 15660 9804
rect 15712 9792 15718 9844
rect 17954 9792 17960 9844
rect 18012 9832 18018 9844
rect 18616 9832 18644 9863
rect 18012 9804 18644 9832
rect 18012 9792 18018 9804
rect 11146 9724 11152 9776
rect 11204 9764 11210 9776
rect 12434 9764 12440 9776
rect 11204 9736 12440 9764
rect 11204 9724 11210 9736
rect 12434 9724 12440 9736
rect 12492 9724 12498 9776
rect 1104 9674 21896 9696
rect 1104 9622 4447 9674
rect 4499 9622 4511 9674
rect 4563 9622 4575 9674
rect 4627 9622 4639 9674
rect 4691 9622 11378 9674
rect 11430 9622 11442 9674
rect 11494 9622 11506 9674
rect 11558 9622 11570 9674
rect 11622 9622 18308 9674
rect 18360 9622 18372 9674
rect 18424 9622 18436 9674
rect 18488 9622 18500 9674
rect 18552 9622 21896 9674
rect 1104 9600 21896 9622
rect 17954 9560 17960 9572
rect 17915 9532 17960 9560
rect 17954 9520 17960 9532
rect 18012 9520 18018 9572
rect 11701 9495 11759 9501
rect 11701 9461 11713 9495
rect 11747 9492 11759 9495
rect 12066 9492 12072 9504
rect 11747 9464 12072 9492
rect 11747 9461 11759 9464
rect 11701 9455 11759 9461
rect 12066 9452 12072 9464
rect 12124 9452 12130 9504
rect 13265 9495 13323 9501
rect 13265 9461 13277 9495
rect 13311 9492 13323 9495
rect 13538 9492 13544 9504
rect 13311 9464 13544 9492
rect 13311 9461 13323 9464
rect 13265 9455 13323 9461
rect 13538 9452 13544 9464
rect 13596 9452 13602 9504
rect 19518 9452 19524 9504
rect 19576 9492 19582 9504
rect 19889 9495 19947 9501
rect 19889 9492 19901 9495
rect 19576 9464 19901 9492
rect 19576 9452 19582 9464
rect 19889 9461 19901 9464
rect 19935 9461 19947 9495
rect 19889 9455 19947 9461
rect 19058 9384 19064 9436
rect 19116 9384 19122 9436
rect 11330 9316 11336 9368
rect 11388 9356 11394 9368
rect 11517 9359 11575 9365
rect 11517 9356 11529 9359
rect 11388 9328 11529 9356
rect 11388 9316 11394 9328
rect 11517 9325 11529 9328
rect 11563 9325 11575 9359
rect 11517 9319 11575 9325
rect 13081 9359 13139 9365
rect 13081 9325 13093 9359
rect 13127 9356 13139 9359
rect 13354 9356 13360 9368
rect 13127 9328 13360 9356
rect 13127 9325 13139 9328
rect 13081 9319 13139 9325
rect 13354 9316 13360 9328
rect 13412 9316 13418 9368
rect 15289 9359 15347 9365
rect 15289 9325 15301 9359
rect 15335 9356 15347 9359
rect 15930 9356 15936 9368
rect 15335 9328 15936 9356
rect 15335 9325 15347 9328
rect 15289 9319 15347 9325
rect 15930 9316 15936 9328
rect 15988 9316 15994 9368
rect 16577 9359 16635 9365
rect 16577 9325 16589 9359
rect 16623 9356 16635 9359
rect 16666 9356 16672 9368
rect 16623 9328 16672 9356
rect 16623 9325 16635 9328
rect 16577 9319 16635 9325
rect 16666 9316 16672 9328
rect 16724 9316 16730 9368
rect 14734 9248 14740 9300
rect 14792 9288 14798 9300
rect 15565 9291 15623 9297
rect 15565 9288 15577 9291
rect 14792 9260 15577 9288
rect 14792 9248 14798 9260
rect 15565 9257 15577 9260
rect 15611 9257 15623 9291
rect 16822 9291 16880 9297
rect 16822 9288 16834 9291
rect 15565 9251 15623 9257
rect 16592 9260 16834 9288
rect 16592 9232 16620 9260
rect 16822 9257 16834 9260
rect 16868 9257 16880 9291
rect 16822 9251 16880 9257
rect 16574 9180 16580 9232
rect 16632 9180 16638 9232
rect 18874 9180 18880 9232
rect 18932 9220 18938 9232
rect 19076 9220 19104 9384
rect 19702 9356 19708 9368
rect 19663 9328 19708 9356
rect 19702 9316 19708 9328
rect 19760 9316 19766 9368
rect 18932 9192 19104 9220
rect 18932 9180 18938 9192
rect 1104 9130 21896 9152
rect 1104 9078 7912 9130
rect 7964 9078 7976 9130
rect 8028 9078 8040 9130
rect 8092 9078 8104 9130
rect 8156 9078 14843 9130
rect 14895 9078 14907 9130
rect 14959 9078 14971 9130
rect 15023 9078 15035 9130
rect 15087 9078 21896 9130
rect 1104 9056 21896 9078
rect 14642 8976 14648 9028
rect 14700 9016 14706 9028
rect 14921 9019 14979 9025
rect 14921 9016 14933 9019
rect 14700 8988 14933 9016
rect 14700 8976 14706 8988
rect 14921 8985 14933 8988
rect 14967 8985 14979 9019
rect 15930 9016 15936 9028
rect 15891 8988 15936 9016
rect 14921 8979 14979 8985
rect 15930 8976 15936 8988
rect 15988 8976 15994 9028
rect 18049 9019 18107 9025
rect 18049 8985 18061 9019
rect 18095 9016 18107 9019
rect 18138 9016 18144 9028
rect 18095 8988 18144 9016
rect 18095 8985 18107 8988
rect 18049 8979 18107 8985
rect 18138 8976 18144 8988
rect 18196 8976 18202 9028
rect 19613 9019 19671 9025
rect 19613 8985 19625 9019
rect 19659 9016 19671 9019
rect 19794 9016 19800 9028
rect 19659 8988 19800 9016
rect 19659 8985 19671 8988
rect 19613 8979 19671 8985
rect 19794 8976 19800 8988
rect 19852 8976 19858 9028
rect 20717 9019 20775 9025
rect 20717 8985 20729 9019
rect 20763 9016 20775 9019
rect 21082 9016 21088 9028
rect 20763 8988 21088 9016
rect 20763 8985 20775 8988
rect 20717 8979 20775 8985
rect 21082 8976 21088 8988
rect 21140 8976 21146 9028
rect 11330 8948 11336 8960
rect 11291 8920 11336 8948
rect 11330 8908 11336 8920
rect 11388 8908 11394 8960
rect 13354 8948 13360 8960
rect 13315 8920 13360 8948
rect 13354 8908 13360 8920
rect 13412 8908 13418 8960
rect 11054 8880 11060 8892
rect 11015 8852 11060 8880
rect 11054 8840 11060 8852
rect 11112 8840 11118 8892
rect 13081 8883 13139 8889
rect 13081 8849 13093 8883
rect 13127 8880 13139 8883
rect 13538 8880 13544 8892
rect 13127 8852 13544 8880
rect 13127 8849 13139 8852
rect 13081 8843 13139 8849
rect 13538 8840 13544 8852
rect 13596 8840 13602 8892
rect 14734 8880 14740 8892
rect 14695 8852 14740 8880
rect 14734 8840 14740 8852
rect 14792 8840 14798 8892
rect 16298 8880 16304 8892
rect 16259 8852 16304 8880
rect 16298 8840 16304 8852
rect 16356 8840 16362 8892
rect 19242 8840 19248 8892
rect 19300 8880 19306 8892
rect 19429 8883 19487 8889
rect 19429 8880 19441 8883
rect 19300 8852 19441 8880
rect 19300 8840 19306 8852
rect 19429 8849 19441 8852
rect 19475 8849 19487 8883
rect 19429 8843 19487 8849
rect 20533 8883 20591 8889
rect 20533 8849 20545 8883
rect 20579 8880 20591 8883
rect 20622 8880 20628 8892
rect 20579 8852 20628 8880
rect 20579 8849 20591 8852
rect 20533 8843 20591 8849
rect 20622 8840 20628 8852
rect 20680 8840 20686 8892
rect 16390 8812 16396 8824
rect 16351 8784 16396 8812
rect 16390 8772 16396 8784
rect 16448 8772 16454 8824
rect 16574 8812 16580 8824
rect 16535 8784 16580 8812
rect 16574 8772 16580 8784
rect 16632 8772 16638 8824
rect 1104 8586 21896 8608
rect 1104 8534 4447 8586
rect 4499 8534 4511 8586
rect 4563 8534 4575 8586
rect 4627 8534 4639 8586
rect 4691 8534 11378 8586
rect 11430 8534 11442 8586
rect 11494 8534 11506 8586
rect 11558 8534 11570 8586
rect 11622 8534 18308 8586
rect 18360 8534 18372 8586
rect 18424 8534 18436 8586
rect 18488 8534 18500 8586
rect 18552 8534 21896 8586
rect 1104 8512 21896 8534
rect 13538 8472 13544 8484
rect 13499 8444 13544 8472
rect 13538 8432 13544 8444
rect 13596 8432 13602 8484
rect 16574 8432 16580 8484
rect 16632 8472 16638 8484
rect 16945 8475 17003 8481
rect 16945 8472 16957 8475
rect 16632 8444 16957 8472
rect 16632 8432 16638 8444
rect 16945 8441 16957 8444
rect 16991 8441 17003 8475
rect 16945 8435 17003 8441
rect 9766 8296 9772 8348
rect 9824 8336 9830 8348
rect 10410 8336 10416 8348
rect 9824 8308 10416 8336
rect 9824 8296 9830 8308
rect 10410 8296 10416 8308
rect 10468 8336 10474 8348
rect 11333 8339 11391 8345
rect 11333 8336 11345 8339
rect 10468 8308 11345 8336
rect 10468 8296 10474 8308
rect 11333 8305 11345 8308
rect 11379 8305 11391 8339
rect 14182 8336 14188 8348
rect 14143 8308 14188 8336
rect 11333 8299 11391 8305
rect 14182 8296 14188 8308
rect 14240 8296 14246 8348
rect 10321 8271 10379 8277
rect 10321 8237 10333 8271
rect 10367 8268 10379 8271
rect 11238 8268 11244 8280
rect 10367 8240 11244 8268
rect 10367 8237 10379 8240
rect 10321 8231 10379 8237
rect 11238 8228 11244 8240
rect 11296 8228 11302 8280
rect 15565 8271 15623 8277
rect 15565 8237 15577 8271
rect 15611 8268 15623 8271
rect 16666 8268 16672 8280
rect 15611 8240 16672 8268
rect 15611 8237 15623 8240
rect 15565 8231 15623 8237
rect 11146 8160 11152 8212
rect 11204 8200 11210 8212
rect 11578 8203 11636 8209
rect 11578 8200 11590 8203
rect 11204 8172 11590 8200
rect 11204 8160 11210 8172
rect 11578 8169 11590 8172
rect 11624 8169 11636 8203
rect 11578 8163 11636 8169
rect 13630 8160 13636 8212
rect 13688 8200 13694 8212
rect 14001 8203 14059 8209
rect 14001 8200 14013 8203
rect 13688 8172 14013 8200
rect 13688 8160 13694 8172
rect 14001 8169 14013 8172
rect 14047 8169 14059 8203
rect 15580 8200 15608 8231
rect 16666 8228 16672 8240
rect 16724 8228 16730 8280
rect 14001 8163 14059 8169
rect 15120 8172 15608 8200
rect 12713 8135 12771 8141
rect 12713 8101 12725 8135
rect 12759 8132 12771 8135
rect 12894 8132 12900 8144
rect 12759 8104 12900 8132
rect 12759 8101 12771 8104
rect 12713 8095 12771 8101
rect 12894 8092 12900 8104
rect 12952 8092 12958 8144
rect 13906 8132 13912 8144
rect 13867 8104 13912 8132
rect 13906 8092 13912 8104
rect 13964 8092 13970 8144
rect 14274 8092 14280 8144
rect 14332 8132 14338 8144
rect 15120 8132 15148 8172
rect 15654 8160 15660 8212
rect 15712 8200 15718 8212
rect 15810 8203 15868 8209
rect 15810 8200 15822 8203
rect 15712 8172 15822 8200
rect 15712 8160 15718 8172
rect 15810 8169 15822 8172
rect 15856 8169 15868 8203
rect 15810 8163 15868 8169
rect 14332 8104 15148 8132
rect 14332 8092 14338 8104
rect 1104 8042 21896 8064
rect 1104 7990 7912 8042
rect 7964 7990 7976 8042
rect 8028 7990 8040 8042
rect 8092 7990 8104 8042
rect 8156 7990 14843 8042
rect 14895 7990 14907 8042
rect 14959 7990 14971 8042
rect 15023 7990 15035 8042
rect 15087 7990 21896 8042
rect 1104 7968 21896 7990
rect 11146 7928 11152 7940
rect 11107 7900 11152 7928
rect 11146 7888 11152 7900
rect 11204 7888 11210 7940
rect 13265 7931 13323 7937
rect 13265 7897 13277 7931
rect 13311 7928 13323 7931
rect 13906 7928 13912 7940
rect 13311 7900 13912 7928
rect 13311 7897 13323 7900
rect 13265 7891 13323 7897
rect 13906 7888 13912 7900
rect 13964 7888 13970 7940
rect 16298 7888 16304 7940
rect 16356 7928 16362 7940
rect 16485 7931 16543 7937
rect 16485 7928 16497 7931
rect 16356 7900 16497 7928
rect 16356 7888 16362 7900
rect 16485 7897 16497 7900
rect 16531 7897 16543 7931
rect 16485 7891 16543 7897
rect 20717 7931 20775 7937
rect 20717 7897 20729 7931
rect 20763 7897 20775 7931
rect 20717 7891 20775 7897
rect 14182 7820 14188 7872
rect 14240 7860 14246 7872
rect 14522 7863 14580 7869
rect 14522 7860 14534 7863
rect 14240 7832 14534 7860
rect 14240 7820 14246 7832
rect 14522 7829 14534 7832
rect 14568 7829 14580 7863
rect 14522 7823 14580 7829
rect 15470 7820 15476 7872
rect 15528 7860 15534 7872
rect 20732 7860 20760 7891
rect 15528 7832 20760 7860
rect 15528 7820 15534 7832
rect 10042 7801 10048 7804
rect 10036 7792 10048 7801
rect 10003 7764 10048 7792
rect 10036 7755 10048 7764
rect 10042 7752 10048 7755
rect 10100 7752 10106 7804
rect 19242 7752 19248 7804
rect 19300 7792 19306 7804
rect 19429 7795 19487 7801
rect 19429 7792 19441 7795
rect 19300 7764 19441 7792
rect 19300 7752 19306 7764
rect 19429 7761 19441 7764
rect 19475 7761 19487 7795
rect 20530 7792 20536 7804
rect 20491 7764 20536 7792
rect 19429 7755 19487 7761
rect 20530 7752 20536 7764
rect 20588 7752 20594 7804
rect 9766 7724 9772 7736
rect 9727 7696 9772 7724
rect 9766 7684 9772 7696
rect 9824 7684 9830 7736
rect 12802 7684 12808 7736
rect 12860 7724 12866 7736
rect 14274 7724 14280 7736
rect 12860 7696 14280 7724
rect 12860 7684 12866 7696
rect 14274 7684 14280 7696
rect 14332 7684 14338 7736
rect 16206 7616 16212 7668
rect 16264 7656 16270 7668
rect 19613 7659 19671 7665
rect 19613 7656 19625 7659
rect 16264 7628 19625 7656
rect 16264 7616 16270 7628
rect 19613 7625 19625 7628
rect 19659 7625 19671 7659
rect 19613 7619 19671 7625
rect 15654 7588 15660 7600
rect 15615 7560 15660 7588
rect 15654 7548 15660 7560
rect 15712 7548 15718 7600
rect 1104 7498 21896 7520
rect 1104 7446 4447 7498
rect 4499 7446 4511 7498
rect 4563 7446 4575 7498
rect 4627 7446 4639 7498
rect 4691 7446 11378 7498
rect 11430 7446 11442 7498
rect 11494 7446 11506 7498
rect 11558 7446 11570 7498
rect 11622 7446 18308 7498
rect 18360 7446 18372 7498
rect 18424 7446 18436 7498
rect 18488 7446 18500 7498
rect 18552 7446 21896 7498
rect 1104 7424 21896 7446
rect 10781 7387 10839 7393
rect 10781 7353 10793 7387
rect 10827 7384 10839 7387
rect 11054 7384 11060 7396
rect 10827 7356 11060 7384
rect 10827 7353 10839 7356
rect 10781 7347 10839 7353
rect 11054 7344 11060 7356
rect 11112 7344 11118 7396
rect 14182 7384 14188 7396
rect 14143 7356 14188 7384
rect 14182 7344 14188 7356
rect 14240 7344 14246 7396
rect 16390 7344 16396 7396
rect 16448 7384 16454 7396
rect 16485 7387 16543 7393
rect 16485 7384 16497 7387
rect 16448 7356 16497 7384
rect 16448 7344 16454 7356
rect 16485 7353 16497 7356
rect 16531 7353 16543 7387
rect 16485 7347 16543 7353
rect 11146 7208 11152 7260
rect 11204 7248 11210 7260
rect 11333 7251 11391 7257
rect 11333 7248 11345 7251
rect 11204 7220 11345 7248
rect 11204 7208 11210 7220
rect 11333 7217 11345 7220
rect 11379 7217 11391 7251
rect 12802 7248 12808 7260
rect 12763 7220 12808 7248
rect 11333 7211 11391 7217
rect 12802 7208 12808 7220
rect 12860 7208 12866 7260
rect 15654 7208 15660 7260
rect 15712 7248 15718 7260
rect 17037 7251 17095 7257
rect 17037 7248 17049 7251
rect 15712 7220 17049 7248
rect 15712 7208 15718 7220
rect 17037 7217 17049 7220
rect 17083 7217 17095 7251
rect 17037 7211 17095 7217
rect 11238 7180 11244 7192
rect 11164 7152 11244 7180
rect 11164 7121 11192 7152
rect 11238 7140 11244 7152
rect 11296 7140 11302 7192
rect 12894 7140 12900 7192
rect 12952 7180 12958 7192
rect 13061 7183 13119 7189
rect 13061 7180 13073 7183
rect 12952 7152 13073 7180
rect 12952 7140 12958 7152
rect 13061 7149 13073 7152
rect 13107 7149 13119 7183
rect 16942 7180 16948 7192
rect 16855 7152 16948 7180
rect 13061 7143 13119 7149
rect 16942 7140 16948 7152
rect 17000 7180 17006 7192
rect 18046 7180 18052 7192
rect 17000 7152 18052 7180
rect 17000 7140 17006 7152
rect 18046 7140 18052 7152
rect 18104 7140 18110 7192
rect 11149 7115 11207 7121
rect 11149 7081 11161 7115
rect 11195 7081 11207 7115
rect 11149 7075 11207 7081
rect 16853 7115 16911 7121
rect 16853 7081 16865 7115
rect 16899 7112 16911 7115
rect 18690 7112 18696 7124
rect 16899 7084 18696 7112
rect 16899 7081 16911 7084
rect 16853 7075 16911 7081
rect 18690 7072 18696 7084
rect 18748 7072 18754 7124
rect 11238 7044 11244 7056
rect 11199 7016 11244 7044
rect 11238 7004 11244 7016
rect 11296 7004 11302 7056
rect 1104 6954 21896 6976
rect 1104 6902 7912 6954
rect 7964 6902 7976 6954
rect 8028 6902 8040 6954
rect 8092 6902 8104 6954
rect 8156 6902 14843 6954
rect 14895 6902 14907 6954
rect 14959 6902 14971 6954
rect 15023 6902 15035 6954
rect 15087 6902 21896 6954
rect 1104 6880 21896 6902
rect 11149 6775 11207 6781
rect 11149 6741 11161 6775
rect 11195 6772 11207 6775
rect 13722 6772 13728 6784
rect 11195 6744 13728 6772
rect 11195 6741 11207 6744
rect 11149 6735 11207 6741
rect 13722 6732 13728 6744
rect 13780 6732 13786 6784
rect 14001 6775 14059 6781
rect 14001 6741 14013 6775
rect 14047 6772 14059 6775
rect 17954 6772 17960 6784
rect 14047 6744 17960 6772
rect 14047 6741 14059 6744
rect 14001 6735 14059 6741
rect 17954 6732 17960 6744
rect 18012 6732 18018 6784
rect 3694 6664 3700 6716
rect 3752 6704 3758 6716
rect 8185 6707 8243 6713
rect 8185 6704 8197 6707
rect 3752 6676 8197 6704
rect 3752 6664 3758 6676
rect 8185 6673 8197 6676
rect 8231 6673 8243 6707
rect 8185 6667 8243 6673
rect 11241 6707 11299 6713
rect 11241 6673 11253 6707
rect 11287 6704 11299 6707
rect 12434 6704 12440 6716
rect 11287 6676 12440 6704
rect 11287 6673 11299 6676
rect 11241 6667 11299 6673
rect 12434 6664 12440 6676
rect 12492 6704 12498 6716
rect 14093 6707 14151 6713
rect 14093 6704 14105 6707
rect 12492 6676 14105 6704
rect 12492 6664 12498 6676
rect 14093 6673 14105 6676
rect 14139 6704 14151 6707
rect 16942 6704 16948 6716
rect 14139 6676 16948 6704
rect 14139 6673 14151 6676
rect 14093 6667 14151 6673
rect 16942 6664 16948 6676
rect 17000 6664 17006 6716
rect 19242 6664 19248 6716
rect 19300 6704 19306 6716
rect 19429 6707 19487 6713
rect 19429 6704 19441 6707
rect 19300 6676 19441 6704
rect 19300 6664 19306 6676
rect 19429 6673 19441 6676
rect 19475 6673 19487 6707
rect 20530 6704 20536 6716
rect 20491 6676 20536 6704
rect 19429 6667 19487 6673
rect 20530 6664 20536 6676
rect 20588 6664 20594 6716
rect 7929 6639 7987 6645
rect 7929 6605 7941 6639
rect 7975 6605 7987 6639
rect 10042 6636 10048 6648
rect 7929 6599 7987 6605
rect 9324 6608 10048 6636
rect 7944 6500 7972 6599
rect 9324 6577 9352 6608
rect 10042 6596 10048 6608
rect 10100 6636 10106 6648
rect 11333 6639 11391 6645
rect 11333 6636 11345 6639
rect 10100 6608 11345 6636
rect 10100 6596 10106 6608
rect 11333 6605 11345 6608
rect 11379 6605 11391 6639
rect 11333 6599 11391 6605
rect 12894 6596 12900 6648
rect 12952 6636 12958 6648
rect 14185 6639 14243 6645
rect 12952 6608 14044 6636
rect 12952 6596 12958 6608
rect 9309 6571 9367 6577
rect 9309 6537 9321 6571
rect 9355 6537 9367 6571
rect 9309 6531 9367 6537
rect 10781 6571 10839 6577
rect 10781 6537 10793 6571
rect 10827 6568 10839 6571
rect 11238 6568 11244 6580
rect 10827 6540 11244 6568
rect 10827 6537 10839 6540
rect 10781 6531 10839 6537
rect 11238 6528 11244 6540
rect 11296 6528 11302 6580
rect 13630 6568 13636 6580
rect 13591 6540 13636 6568
rect 13630 6528 13636 6540
rect 13688 6528 13694 6580
rect 14016 6568 14044 6608
rect 14185 6605 14197 6639
rect 14231 6605 14243 6639
rect 14185 6599 14243 6605
rect 14200 6568 14228 6599
rect 14016 6540 14228 6568
rect 16482 6528 16488 6580
rect 16540 6568 16546 6580
rect 19613 6571 19671 6577
rect 19613 6568 19625 6571
rect 16540 6540 19625 6568
rect 16540 6528 16546 6540
rect 19613 6537 19625 6540
rect 19659 6537 19671 6571
rect 19613 6531 19671 6537
rect 9766 6500 9772 6512
rect 7944 6472 9772 6500
rect 9766 6460 9772 6472
rect 9824 6460 9830 6512
rect 14550 6460 14556 6512
rect 14608 6500 14614 6512
rect 20717 6503 20775 6509
rect 20717 6500 20729 6503
rect 14608 6472 20729 6500
rect 14608 6460 14614 6472
rect 20717 6469 20729 6472
rect 20763 6469 20775 6503
rect 20717 6463 20775 6469
rect 1104 6410 21896 6432
rect 1104 6358 4447 6410
rect 4499 6358 4511 6410
rect 4563 6358 4575 6410
rect 4627 6358 4639 6410
rect 4691 6358 11378 6410
rect 11430 6358 11442 6410
rect 11494 6358 11506 6410
rect 11558 6358 11570 6410
rect 11622 6358 18308 6410
rect 18360 6358 18372 6410
rect 18424 6358 18436 6410
rect 18488 6358 18500 6410
rect 18552 6358 21896 6410
rect 1104 6336 21896 6358
rect 1104 5866 21896 5888
rect 1104 5814 7912 5866
rect 7964 5814 7976 5866
rect 8028 5814 8040 5866
rect 8092 5814 8104 5866
rect 8156 5814 14843 5866
rect 14895 5814 14907 5866
rect 14959 5814 14971 5866
rect 15023 5814 15035 5866
rect 15087 5814 21896 5866
rect 1104 5792 21896 5814
rect 13538 5712 13544 5764
rect 13596 5752 13602 5764
rect 20717 5755 20775 5761
rect 20717 5752 20729 5755
rect 13596 5724 20729 5752
rect 13596 5712 13602 5724
rect 20717 5721 20729 5724
rect 20763 5721 20775 5755
rect 20717 5715 20775 5721
rect 20530 5616 20536 5628
rect 20491 5588 20536 5616
rect 20530 5576 20536 5588
rect 20588 5576 20594 5628
rect 1104 5322 21896 5344
rect 1104 5270 4447 5322
rect 4499 5270 4511 5322
rect 4563 5270 4575 5322
rect 4627 5270 4639 5322
rect 4691 5270 11378 5322
rect 11430 5270 11442 5322
rect 11494 5270 11506 5322
rect 11558 5270 11570 5322
rect 11622 5270 18308 5322
rect 18360 5270 18372 5322
rect 18424 5270 18436 5322
rect 18488 5270 18500 5322
rect 18552 5270 21896 5322
rect 1104 5248 21896 5270
rect 1104 4778 21896 4800
rect 1104 4726 7912 4778
rect 7964 4726 7976 4778
rect 8028 4726 8040 4778
rect 8092 4726 8104 4778
rect 8156 4726 14843 4778
rect 14895 4726 14907 4778
rect 14959 4726 14971 4778
rect 15023 4726 15035 4778
rect 15087 4726 21896 4778
rect 1104 4704 21896 4726
rect 13173 4667 13231 4673
rect 13173 4633 13185 4667
rect 13219 4664 13231 4667
rect 13262 4664 13268 4676
rect 13219 4636 13268 4664
rect 13219 4633 13231 4636
rect 13173 4627 13231 4633
rect 13262 4624 13268 4636
rect 13320 4624 13326 4676
rect 12989 4531 13047 4537
rect 12989 4497 13001 4531
rect 13035 4528 13047 4531
rect 13814 4528 13820 4540
rect 13035 4500 13820 4528
rect 13035 4497 13047 4500
rect 12989 4491 13047 4497
rect 13814 4488 13820 4500
rect 13872 4488 13878 4540
rect 1104 4234 21896 4256
rect 1104 4182 4447 4234
rect 4499 4182 4511 4234
rect 4563 4182 4575 4234
rect 4627 4182 4639 4234
rect 4691 4182 11378 4234
rect 11430 4182 11442 4234
rect 11494 4182 11506 4234
rect 11558 4182 11570 4234
rect 11622 4182 18308 4234
rect 18360 4182 18372 4234
rect 18424 4182 18436 4234
rect 18488 4182 18500 4234
rect 18552 4182 21896 4234
rect 1104 4160 21896 4182
rect 13814 3944 13820 3996
rect 13872 3984 13878 3996
rect 17954 3984 17960 3996
rect 13872 3956 17960 3984
rect 13872 3944 13878 3956
rect 17954 3944 17960 3956
rect 18012 3944 18018 3996
rect 13722 3876 13728 3928
rect 13780 3916 13786 3928
rect 18046 3916 18052 3928
rect 13780 3888 18052 3916
rect 13780 3876 13786 3888
rect 18046 3876 18052 3888
rect 18104 3876 18110 3928
rect 1104 3690 21896 3712
rect 1104 3638 7912 3690
rect 7964 3638 7976 3690
rect 8028 3638 8040 3690
rect 8092 3638 8104 3690
rect 8156 3638 14843 3690
rect 14895 3638 14907 3690
rect 14959 3638 14971 3690
rect 15023 3638 15035 3690
rect 15087 3638 21896 3690
rect 1104 3616 21896 3638
rect 20717 3579 20775 3585
rect 20717 3545 20729 3579
rect 20763 3576 20775 3579
rect 21174 3576 21180 3588
rect 20763 3548 21180 3576
rect 20763 3545 20775 3548
rect 20717 3539 20775 3545
rect 21174 3536 21180 3548
rect 21232 3536 21238 3588
rect 20530 3440 20536 3452
rect 20491 3412 20536 3440
rect 20530 3400 20536 3412
rect 20588 3400 20594 3452
rect 1104 3146 21896 3168
rect 1104 3094 4447 3146
rect 4499 3094 4511 3146
rect 4563 3094 4575 3146
rect 4627 3094 4639 3146
rect 4691 3094 11378 3146
rect 11430 3094 11442 3146
rect 11494 3094 11506 3146
rect 11558 3094 11570 3146
rect 11622 3094 18308 3146
rect 18360 3094 18372 3146
rect 18424 3094 18436 3146
rect 18488 3094 18500 3146
rect 18552 3094 21896 3146
rect 1104 3072 21896 3094
rect 1104 2602 21896 2624
rect 1104 2550 7912 2602
rect 7964 2550 7976 2602
rect 8028 2550 8040 2602
rect 8092 2550 8104 2602
rect 8156 2550 14843 2602
rect 14895 2550 14907 2602
rect 14959 2550 14971 2602
rect 15023 2550 15035 2602
rect 15087 2550 21896 2602
rect 1104 2528 21896 2550
rect 15746 2448 15752 2500
rect 15804 2488 15810 2500
rect 19242 2488 19248 2500
rect 15804 2460 19248 2488
rect 15804 2448 15810 2460
rect 19242 2448 19248 2460
rect 19300 2448 19306 2500
rect 1104 2058 21896 2080
rect 1104 2006 4447 2058
rect 4499 2006 4511 2058
rect 4563 2006 4575 2058
rect 4627 2006 4639 2058
rect 4691 2006 11378 2058
rect 11430 2006 11442 2058
rect 11494 2006 11506 2058
rect 11558 2006 11570 2058
rect 11622 2006 18308 2058
rect 18360 2006 18372 2058
rect 18424 2006 18436 2058
rect 18488 2006 18500 2058
rect 18552 2006 21896 2058
rect 1104 1984 21896 2006
rect 15838 1156 15844 1208
rect 15896 1196 15902 1208
rect 19242 1196 19248 1208
rect 15896 1168 19248 1196
rect 15896 1156 15902 1168
rect 19242 1156 19248 1168
rect 19300 1156 19306 1208
<< via1 >>
rect 4447 20502 4499 20554
rect 4511 20502 4563 20554
rect 4575 20502 4627 20554
rect 4639 20502 4691 20554
rect 11378 20502 11430 20554
rect 11442 20502 11494 20554
rect 11506 20502 11558 20554
rect 11570 20502 11622 20554
rect 18308 20502 18360 20554
rect 18372 20502 18424 20554
rect 18436 20502 18488 20554
rect 18500 20502 18552 20554
rect 17868 20400 17920 20452
rect 8208 20264 8260 20316
rect 5816 20196 5868 20248
rect 11428 20239 11480 20248
rect 7104 20128 7156 20180
rect 11428 20205 11437 20239
rect 11437 20205 11471 20239
rect 11471 20205 11480 20239
rect 11428 20196 11480 20205
rect 13084 20196 13136 20248
rect 13268 20264 13320 20316
rect 16120 20264 16172 20316
rect 13452 20196 13504 20248
rect 7196 20103 7248 20112
rect 7196 20069 7205 20103
rect 7205 20069 7239 20103
rect 7239 20069 7248 20103
rect 7196 20060 7248 20069
rect 7288 20060 7340 20112
rect 11152 20060 11204 20112
rect 18696 20128 18748 20180
rect 13636 20060 13688 20112
rect 16304 20060 16356 20112
rect 16488 20103 16540 20112
rect 16488 20069 16497 20103
rect 16497 20069 16531 20103
rect 16531 20069 16540 20103
rect 16488 20060 16540 20069
rect 19248 20060 19300 20112
rect 7912 19958 7964 20010
rect 7976 19958 8028 20010
rect 8040 19958 8092 20010
rect 8104 19958 8156 20010
rect 14843 19958 14895 20010
rect 14907 19958 14959 20010
rect 14971 19958 15023 20010
rect 15035 19958 15087 20010
rect 9220 19856 9272 19908
rect 15200 19856 15252 19908
rect 16028 19899 16080 19908
rect 16028 19865 16037 19899
rect 16037 19865 16071 19899
rect 16071 19865 16080 19899
rect 16028 19856 16080 19865
rect 16396 19856 16448 19908
rect 19432 19856 19484 19908
rect 7196 19788 7248 19840
rect 12348 19788 12400 19840
rect 15108 19788 15160 19840
rect 7472 19720 7524 19772
rect 8760 19720 8812 19772
rect 9220 19720 9272 19772
rect 12992 19720 13044 19772
rect 13268 19720 13320 19772
rect 15844 19720 15896 19772
rect 16304 19720 16356 19772
rect 6828 19695 6880 19704
rect 6828 19661 6837 19695
rect 6837 19661 6871 19695
rect 6871 19661 6880 19695
rect 6828 19652 6880 19661
rect 9128 19695 9180 19704
rect 9128 19661 9137 19695
rect 9137 19661 9171 19695
rect 9171 19661 9180 19695
rect 9128 19652 9180 19661
rect 11060 19652 11112 19704
rect 12532 19652 12584 19704
rect 15660 19652 15712 19704
rect 16396 19652 16448 19704
rect 19984 19695 20036 19704
rect 19984 19661 19993 19695
rect 19993 19661 20027 19695
rect 20027 19661 20036 19695
rect 19984 19652 20036 19661
rect 16488 19584 16540 19636
rect 8208 19559 8260 19568
rect 8208 19525 8217 19559
rect 8217 19525 8251 19559
rect 8251 19525 8260 19559
rect 8208 19516 8260 19525
rect 10508 19559 10560 19568
rect 10508 19525 10517 19559
rect 10517 19525 10551 19559
rect 10551 19525 10560 19559
rect 10508 19516 10560 19525
rect 15384 19516 15436 19568
rect 4447 19414 4499 19466
rect 4511 19414 4563 19466
rect 4575 19414 4627 19466
rect 4639 19414 4691 19466
rect 11378 19414 11430 19466
rect 11442 19414 11494 19466
rect 11506 19414 11558 19466
rect 11570 19414 11622 19466
rect 18308 19414 18360 19466
rect 18372 19414 18424 19466
rect 18436 19414 18488 19466
rect 18500 19414 18552 19466
rect 8760 19355 8812 19364
rect 8760 19321 8769 19355
rect 8769 19321 8803 19355
rect 8803 19321 8812 19355
rect 8760 19312 8812 19321
rect 6276 19176 6328 19228
rect 6828 19176 6880 19228
rect 7288 19108 7340 19160
rect 8208 19108 8260 19160
rect 9128 19108 9180 19160
rect 10508 19108 10560 19160
rect 10784 19108 10836 19160
rect 12532 19312 12584 19364
rect 13268 19355 13320 19364
rect 13268 19321 13277 19355
rect 13277 19321 13311 19355
rect 13311 19321 13320 19355
rect 13268 19312 13320 19321
rect 13912 19312 13964 19364
rect 16396 19312 16448 19364
rect 12900 19244 12952 19296
rect 13636 19244 13688 19296
rect 17960 19287 18012 19296
rect 17960 19253 17969 19287
rect 17969 19253 18003 19287
rect 18003 19253 18012 19287
rect 17960 19244 18012 19253
rect 1400 19040 1452 19092
rect 3608 19040 3660 19092
rect 9496 19040 9548 19092
rect 10140 19040 10192 19092
rect 15108 19176 15160 19228
rect 17500 19176 17552 19228
rect 15292 19151 15344 19160
rect 8300 18972 8352 19024
rect 8668 18972 8720 19024
rect 10968 18972 11020 19024
rect 12992 19040 13044 19092
rect 15292 19117 15301 19151
rect 15301 19117 15335 19151
rect 15335 19117 15344 19151
rect 15292 19108 15344 19117
rect 15384 19108 15436 19160
rect 15568 19151 15620 19160
rect 15568 19117 15591 19151
rect 15591 19117 15620 19151
rect 18052 19176 18104 19228
rect 15568 19108 15620 19117
rect 18144 19108 18196 19160
rect 15200 19040 15252 19092
rect 16764 19040 16816 19092
rect 19984 19040 20036 19092
rect 12348 18972 12400 19024
rect 12808 18972 12860 19024
rect 14372 18972 14424 19024
rect 16120 18972 16172 19024
rect 17040 18972 17092 19024
rect 21088 18972 21140 19024
rect 7912 18870 7964 18922
rect 7976 18870 8028 18922
rect 8040 18870 8092 18922
rect 8104 18870 8156 18922
rect 14843 18870 14895 18922
rect 14907 18870 14959 18922
rect 14971 18870 15023 18922
rect 15035 18870 15087 18922
rect 2504 18768 2556 18820
rect 5540 18768 5592 18820
rect 7104 18768 7156 18820
rect 7380 18811 7432 18820
rect 7380 18777 7389 18811
rect 7389 18777 7423 18811
rect 7423 18777 7432 18811
rect 7380 18768 7432 18777
rect 7564 18768 7616 18820
rect 7748 18768 7800 18820
rect 10140 18811 10192 18820
rect 10140 18777 10149 18811
rect 10149 18777 10183 18811
rect 10183 18777 10192 18811
rect 10140 18768 10192 18777
rect 11060 18768 11112 18820
rect 11704 18768 11756 18820
rect 12348 18768 12400 18820
rect 12900 18768 12952 18820
rect 14372 18768 14424 18820
rect 17592 18768 17644 18820
rect 18052 18811 18104 18820
rect 18052 18777 18061 18811
rect 18061 18777 18095 18811
rect 18095 18777 18104 18811
rect 18052 18768 18104 18777
rect 18512 18811 18564 18820
rect 18512 18777 18521 18811
rect 18521 18777 18555 18811
rect 18555 18777 18564 18811
rect 18512 18768 18564 18777
rect 18604 18768 18656 18820
rect 21364 18768 21416 18820
rect 4804 18700 4856 18752
rect 8576 18700 8628 18752
rect 4160 18632 4212 18684
rect 13084 18700 13136 18752
rect 8944 18675 8996 18684
rect 8944 18641 8953 18675
rect 8953 18641 8987 18675
rect 8987 18641 8996 18675
rect 8944 18632 8996 18641
rect 13176 18632 13228 18684
rect 16019 18675 16071 18684
rect 16019 18641 16051 18675
rect 16051 18641 16071 18675
rect 16019 18632 16071 18641
rect 17868 18632 17920 18684
rect 18420 18675 18472 18684
rect 848 18564 900 18616
rect 7104 18564 7156 18616
rect 7472 18564 7524 18616
rect 9220 18607 9272 18616
rect 9220 18573 9229 18607
rect 9229 18573 9263 18607
rect 9263 18573 9272 18607
rect 9220 18564 9272 18573
rect 296 18496 348 18548
rect 8392 18496 8444 18548
rect 10784 18607 10836 18616
rect 10784 18573 10793 18607
rect 10793 18573 10827 18607
rect 10827 18573 10836 18607
rect 10784 18564 10836 18573
rect 11060 18564 11112 18616
rect 12992 18607 13044 18616
rect 12992 18573 13001 18607
rect 13001 18573 13035 18607
rect 13035 18573 13044 18607
rect 12992 18564 13044 18573
rect 15292 18564 15344 18616
rect 17500 18564 17552 18616
rect 18420 18641 18429 18675
rect 18429 18641 18463 18675
rect 18463 18641 18472 18675
rect 18420 18632 18472 18641
rect 19432 18632 19484 18684
rect 19800 18564 19852 18616
rect 11244 18428 11296 18480
rect 12532 18428 12584 18480
rect 14740 18428 14792 18480
rect 17684 18428 17736 18480
rect 17776 18428 17828 18480
rect 20996 18428 21048 18480
rect 4447 18326 4499 18378
rect 4511 18326 4563 18378
rect 4575 18326 4627 18378
rect 4639 18326 4691 18378
rect 11378 18326 11430 18378
rect 11442 18326 11494 18378
rect 11506 18326 11558 18378
rect 11570 18326 11622 18378
rect 18308 18326 18360 18378
rect 18372 18326 18424 18378
rect 18436 18326 18488 18378
rect 18500 18326 18552 18378
rect 1952 18224 2004 18276
rect 7104 18224 7156 18276
rect 9680 18224 9732 18276
rect 12532 18224 12584 18276
rect 12624 18224 12676 18276
rect 13268 18224 13320 18276
rect 13636 18224 13688 18276
rect 15384 18224 15436 18276
rect 15476 18224 15528 18276
rect 7656 18156 7708 18208
rect 10232 18156 10284 18208
rect 10324 18156 10376 18208
rect 11704 18156 11756 18208
rect 14004 18156 14056 18208
rect 18604 18224 18656 18276
rect 7656 18020 7708 18072
rect 9864 18131 9916 18140
rect 9864 18097 9873 18131
rect 9873 18097 9907 18131
rect 9907 18097 9916 18131
rect 9864 18088 9916 18097
rect 8392 18020 8444 18072
rect 10692 18020 10744 18072
rect 10876 18020 10928 18072
rect 6276 17952 6328 18004
rect 7380 17952 7432 18004
rect 8576 17952 8628 18004
rect 13360 18088 13412 18140
rect 16488 18156 16540 18208
rect 18236 18156 18288 18208
rect 18880 18156 18932 18208
rect 13912 18020 13964 18072
rect 3056 17884 3108 17936
rect 7288 17884 7340 17936
rect 7748 17927 7800 17936
rect 7748 17893 7757 17927
rect 7757 17893 7791 17927
rect 7791 17893 7800 17927
rect 7748 17884 7800 17893
rect 8208 17927 8260 17936
rect 8208 17893 8217 17927
rect 8217 17893 8251 17927
rect 8251 17893 8260 17927
rect 8208 17884 8260 17893
rect 8300 17884 8352 17936
rect 10784 17884 10836 17936
rect 11152 17884 11204 17936
rect 11244 17884 11296 17936
rect 13636 17952 13688 18004
rect 14280 18020 14332 18072
rect 14740 18020 14792 18072
rect 17040 18020 17092 18072
rect 17224 18063 17276 18072
rect 17224 18029 17233 18063
rect 17233 18029 17267 18063
rect 17267 18029 17276 18063
rect 17224 18020 17276 18029
rect 18972 18088 19024 18140
rect 19064 18088 19116 18140
rect 19892 18088 19944 18140
rect 20352 18088 20404 18140
rect 18880 18020 18932 18072
rect 19708 18063 19760 18072
rect 19708 18029 19717 18063
rect 19717 18029 19751 18063
rect 19751 18029 19760 18063
rect 19708 18020 19760 18029
rect 17316 17952 17368 18004
rect 17500 17995 17552 18004
rect 17500 17961 17534 17995
rect 17534 17961 17552 17995
rect 17500 17952 17552 17961
rect 17684 17952 17736 18004
rect 18696 17952 18748 18004
rect 19616 17952 19668 18004
rect 20444 17952 20496 18004
rect 14004 17884 14056 17936
rect 18236 17884 18288 17936
rect 18604 17927 18656 17936
rect 18604 17893 18613 17927
rect 18613 17893 18647 17927
rect 18647 17893 18656 17927
rect 18604 17884 18656 17893
rect 19156 17884 19208 17936
rect 21180 17884 21232 17936
rect 22652 17884 22704 17936
rect 7912 17782 7964 17834
rect 7976 17782 8028 17834
rect 8040 17782 8092 17834
rect 8104 17782 8156 17834
rect 14843 17782 14895 17834
rect 14907 17782 14959 17834
rect 14971 17782 15023 17834
rect 15035 17782 15087 17834
rect 8208 17680 8260 17732
rect 9496 17680 9548 17732
rect 12716 17680 12768 17732
rect 13084 17680 13136 17732
rect 13360 17680 13412 17732
rect 18052 17680 18104 17732
rect 7012 17612 7064 17664
rect 7196 17544 7248 17596
rect 4068 17476 4120 17528
rect 8944 17544 8996 17596
rect 9588 17587 9640 17596
rect 9588 17553 9597 17587
rect 9597 17553 9631 17587
rect 9631 17553 9640 17587
rect 9588 17544 9640 17553
rect 13176 17544 13228 17596
rect 15844 17544 15896 17596
rect 16028 17544 16080 17596
rect 7472 17519 7524 17528
rect 7472 17485 7481 17519
rect 7481 17485 7515 17519
rect 7515 17485 7524 17519
rect 9772 17519 9824 17528
rect 7472 17476 7524 17485
rect 9772 17485 9781 17519
rect 9781 17485 9815 17519
rect 9815 17485 9824 17519
rect 9772 17476 9824 17485
rect 12992 17519 13044 17528
rect 12992 17485 13001 17519
rect 13001 17485 13035 17519
rect 13035 17485 13044 17519
rect 12992 17476 13044 17485
rect 15108 17519 15160 17528
rect 15108 17485 15117 17519
rect 15117 17485 15151 17519
rect 15151 17485 15160 17519
rect 15108 17476 15160 17485
rect 17040 17612 17092 17664
rect 16856 17587 16908 17596
rect 16856 17553 16865 17587
rect 16865 17553 16899 17587
rect 16899 17553 16908 17587
rect 16856 17544 16908 17553
rect 17868 17544 17920 17596
rect 19892 17587 19944 17596
rect 19892 17553 19901 17587
rect 19901 17553 19935 17587
rect 19935 17553 19944 17587
rect 19892 17544 19944 17553
rect 18604 17476 18656 17528
rect 9864 17408 9916 17460
rect 17868 17408 17920 17460
rect 18144 17451 18196 17460
rect 18144 17417 18153 17451
rect 18153 17417 18187 17451
rect 18187 17417 18196 17451
rect 18144 17408 18196 17417
rect 10508 17340 10560 17392
rect 12440 17383 12492 17392
rect 12440 17349 12449 17383
rect 12449 17349 12483 17383
rect 12483 17349 12492 17383
rect 12440 17340 12492 17349
rect 15752 17340 15804 17392
rect 17960 17340 18012 17392
rect 20996 17340 21048 17392
rect 22100 17340 22152 17392
rect 4447 17238 4499 17290
rect 4511 17238 4563 17290
rect 4575 17238 4627 17290
rect 4639 17238 4691 17290
rect 11378 17238 11430 17290
rect 11442 17238 11494 17290
rect 11506 17238 11558 17290
rect 11570 17238 11622 17290
rect 18308 17238 18360 17290
rect 18372 17238 18424 17290
rect 18436 17238 18488 17290
rect 18500 17238 18552 17290
rect 7656 17179 7708 17188
rect 7656 17145 7665 17179
rect 7665 17145 7699 17179
rect 7699 17145 7708 17179
rect 7656 17136 7708 17145
rect 15108 17136 15160 17188
rect 18144 17136 18196 17188
rect 18788 17136 18840 17188
rect 12992 17068 13044 17120
rect 6276 16975 6328 16984
rect 6276 16941 6285 16975
rect 6285 16941 6319 16975
rect 6319 16941 6328 16975
rect 6276 16932 6328 16941
rect 7104 16932 7156 16984
rect 7472 16932 7524 16984
rect 9128 16932 9180 16984
rect 11244 16932 11296 16984
rect 15292 16975 15344 16984
rect 10600 16864 10652 16916
rect 12532 16796 12584 16848
rect 15292 16941 15301 16975
rect 15301 16941 15335 16975
rect 15335 16941 15344 16975
rect 15292 16932 15344 16941
rect 16856 17000 16908 17052
rect 19064 16932 19116 16984
rect 19524 16975 19576 16984
rect 19524 16941 19533 16975
rect 19533 16941 19567 16975
rect 19567 16941 19576 16975
rect 19524 16932 19576 16941
rect 13728 16864 13780 16916
rect 15200 16864 15252 16916
rect 18972 16864 19024 16916
rect 16028 16796 16080 16848
rect 19248 16796 19300 16848
rect 7912 16694 7964 16746
rect 7976 16694 8028 16746
rect 8040 16694 8092 16746
rect 8104 16694 8156 16746
rect 14843 16694 14895 16746
rect 14907 16694 14959 16746
rect 14971 16694 15023 16746
rect 15035 16694 15087 16746
rect 7380 16635 7432 16644
rect 7380 16601 7389 16635
rect 7389 16601 7423 16635
rect 7423 16601 7432 16635
rect 7380 16592 7432 16601
rect 5264 16524 5316 16576
rect 9772 16524 9824 16576
rect 10600 16592 10652 16644
rect 11704 16592 11756 16644
rect 13728 16592 13780 16644
rect 15200 16592 15252 16644
rect 16580 16592 16632 16644
rect 16028 16567 16080 16576
rect 11244 16456 11296 16508
rect 12532 16456 12584 16508
rect 12992 16456 13044 16508
rect 16028 16533 16062 16567
rect 16062 16533 16080 16567
rect 16028 16524 16080 16533
rect 9128 16431 9180 16440
rect 8392 16252 8444 16304
rect 9128 16397 9137 16431
rect 9137 16397 9171 16431
rect 9171 16397 9180 16431
rect 9128 16388 9180 16397
rect 11060 16388 11112 16440
rect 19708 16524 19760 16576
rect 15292 16388 15344 16440
rect 18512 16388 18564 16440
rect 17592 16320 17644 16372
rect 17316 16252 17368 16304
rect 18052 16295 18104 16304
rect 18052 16261 18061 16295
rect 18061 16261 18095 16295
rect 18095 16261 18104 16295
rect 18052 16252 18104 16261
rect 4447 16150 4499 16202
rect 4511 16150 4563 16202
rect 4575 16150 4627 16202
rect 4639 16150 4691 16202
rect 11378 16150 11430 16202
rect 11442 16150 11494 16202
rect 11506 16150 11558 16202
rect 11570 16150 11622 16202
rect 18308 16150 18360 16202
rect 18372 16150 18424 16202
rect 18436 16150 18488 16202
rect 18500 16150 18552 16202
rect 7104 16091 7156 16100
rect 7104 16057 7113 16091
rect 7113 16057 7147 16091
rect 7147 16057 7156 16091
rect 7104 16048 7156 16057
rect 19524 16048 19576 16100
rect 12624 15980 12676 16032
rect 16580 15980 16632 16032
rect 10600 15912 10652 15964
rect 12440 15912 12492 15964
rect 13728 15912 13780 15964
rect 16028 15912 16080 15964
rect 6276 15844 6328 15896
rect 11060 15844 11112 15896
rect 12716 15844 12768 15896
rect 17316 15887 17368 15896
rect 15752 15776 15804 15828
rect 10508 15708 10560 15760
rect 15844 15708 15896 15760
rect 17316 15853 17325 15887
rect 17325 15853 17359 15887
rect 17359 15853 17368 15887
rect 17316 15844 17368 15853
rect 17592 15887 17644 15896
rect 17592 15853 17626 15887
rect 17626 15853 17644 15887
rect 17592 15844 17644 15853
rect 19524 15887 19576 15896
rect 19524 15853 19533 15887
rect 19533 15853 19567 15887
rect 19567 15853 19576 15887
rect 19524 15844 19576 15853
rect 17684 15776 17736 15828
rect 18788 15708 18840 15760
rect 7912 15606 7964 15658
rect 7976 15606 8028 15658
rect 8040 15606 8092 15658
rect 8104 15606 8156 15658
rect 14843 15606 14895 15658
rect 14907 15606 14959 15658
rect 14971 15606 15023 15658
rect 15035 15606 15087 15658
rect 7288 15547 7340 15556
rect 7288 15513 7297 15547
rect 7297 15513 7331 15547
rect 7331 15513 7340 15547
rect 7288 15504 7340 15513
rect 9772 15547 9824 15556
rect 9772 15513 9781 15547
rect 9781 15513 9815 15547
rect 9815 15513 9824 15547
rect 9772 15504 9824 15513
rect 11244 15504 11296 15556
rect 12624 15504 12676 15556
rect 15844 15547 15896 15556
rect 7564 15436 7616 15488
rect 8668 15411 8720 15420
rect 8668 15377 8702 15411
rect 8702 15377 8720 15411
rect 8668 15368 8720 15377
rect 9588 15436 9640 15488
rect 15844 15513 15853 15547
rect 15853 15513 15887 15547
rect 15887 15513 15896 15547
rect 15844 15504 15896 15513
rect 17960 15504 18012 15556
rect 18052 15504 18104 15556
rect 10508 15368 10560 15420
rect 13084 15368 13136 15420
rect 19432 15436 19484 15488
rect 15200 15368 15252 15420
rect 17684 15368 17736 15420
rect 19248 15368 19300 15420
rect 19984 15411 20036 15420
rect 19984 15377 19993 15411
rect 19993 15377 20027 15411
rect 20027 15377 20036 15411
rect 19984 15368 20036 15377
rect 7472 15343 7524 15352
rect 7472 15309 7481 15343
rect 7481 15309 7515 15343
rect 7515 15309 7524 15343
rect 7472 15300 7524 15309
rect 8392 15343 8444 15352
rect 8392 15309 8401 15343
rect 8401 15309 8435 15343
rect 8435 15309 8444 15343
rect 8392 15300 8444 15309
rect 10600 15343 10652 15352
rect 10600 15309 10609 15343
rect 10609 15309 10643 15343
rect 10643 15309 10652 15343
rect 10600 15300 10652 15309
rect 13452 15300 13504 15352
rect 14556 15343 14608 15352
rect 14556 15309 14565 15343
rect 14565 15309 14599 15343
rect 14599 15309 14608 15343
rect 14556 15300 14608 15309
rect 18788 15343 18840 15352
rect 18788 15309 18797 15343
rect 18797 15309 18831 15343
rect 18831 15309 18840 15343
rect 18788 15300 18840 15309
rect 18880 15300 18932 15352
rect 19524 15232 19576 15284
rect 7748 15164 7800 15216
rect 13912 15207 13964 15216
rect 13912 15173 13921 15207
rect 13921 15173 13955 15207
rect 13955 15173 13964 15207
rect 13912 15164 13964 15173
rect 19340 15164 19392 15216
rect 19892 15164 19944 15216
rect 4447 15062 4499 15114
rect 4511 15062 4563 15114
rect 4575 15062 4627 15114
rect 4639 15062 4691 15114
rect 11378 15062 11430 15114
rect 11442 15062 11494 15114
rect 11506 15062 11558 15114
rect 11570 15062 11622 15114
rect 18308 15062 18360 15114
rect 18372 15062 18424 15114
rect 18436 15062 18488 15114
rect 18500 15062 18552 15114
rect 13452 14960 13504 15012
rect 18696 14960 18748 15012
rect 19432 14960 19484 15012
rect 8668 14892 8720 14944
rect 11152 14824 11204 14876
rect 11888 14867 11940 14876
rect 11888 14833 11897 14867
rect 11897 14833 11931 14867
rect 11931 14833 11940 14867
rect 11888 14824 11940 14833
rect 6276 14756 6328 14808
rect 8392 14756 8444 14808
rect 10600 14756 10652 14808
rect 12532 14824 12584 14876
rect 14556 14824 14608 14876
rect 7472 14688 7524 14740
rect 8208 14688 8260 14740
rect 18880 14824 18932 14876
rect 19064 14824 19116 14876
rect 19432 14824 19484 14876
rect 17408 14756 17460 14808
rect 19708 14867 19760 14876
rect 19708 14833 19717 14867
rect 19717 14833 19751 14867
rect 19751 14833 19760 14867
rect 19708 14824 19760 14833
rect 19340 14688 19392 14740
rect 7748 14620 7800 14672
rect 11244 14620 11296 14672
rect 14188 14663 14240 14672
rect 14188 14629 14197 14663
rect 14197 14629 14231 14663
rect 14231 14629 14240 14663
rect 14188 14620 14240 14629
rect 15292 14663 15344 14672
rect 15292 14629 15301 14663
rect 15301 14629 15335 14663
rect 15335 14629 15344 14663
rect 15292 14620 15344 14629
rect 15660 14663 15712 14672
rect 15660 14629 15669 14663
rect 15669 14629 15703 14663
rect 15703 14629 15712 14663
rect 15660 14620 15712 14629
rect 15844 14620 15896 14672
rect 18604 14663 18656 14672
rect 18604 14629 18613 14663
rect 18613 14629 18647 14663
rect 18647 14629 18656 14663
rect 18604 14620 18656 14629
rect 7912 14518 7964 14570
rect 7976 14518 8028 14570
rect 8040 14518 8092 14570
rect 8104 14518 8156 14570
rect 14843 14518 14895 14570
rect 14907 14518 14959 14570
rect 14971 14518 15023 14570
rect 15035 14518 15087 14570
rect 8208 14459 8260 14468
rect 8208 14425 8217 14459
rect 8217 14425 8251 14459
rect 8251 14425 8260 14459
rect 8208 14416 8260 14425
rect 14556 14416 14608 14468
rect 15660 14416 15712 14468
rect 14188 14348 14240 14400
rect 7472 14280 7524 14332
rect 8392 14280 8444 14332
rect 11888 14280 11940 14332
rect 19064 14416 19116 14468
rect 19156 14280 19208 14332
rect 20444 14280 20496 14332
rect 10876 14076 10928 14128
rect 13728 14076 13780 14128
rect 17316 14076 17368 14128
rect 20628 14076 20680 14128
rect 4447 13974 4499 14026
rect 4511 13974 4563 14026
rect 4575 13974 4627 14026
rect 4639 13974 4691 14026
rect 11378 13974 11430 14026
rect 11442 13974 11494 14026
rect 11506 13974 11558 14026
rect 11570 13974 11622 14026
rect 18308 13974 18360 14026
rect 18372 13974 18424 14026
rect 18436 13974 18488 14026
rect 18500 13974 18552 14026
rect 13084 13915 13136 13924
rect 13084 13881 13093 13915
rect 13093 13881 13127 13915
rect 13127 13881 13136 13915
rect 13084 13872 13136 13881
rect 8852 13804 8904 13856
rect 11336 13804 11388 13856
rect 7472 13779 7524 13788
rect 7472 13745 7481 13779
rect 7481 13745 7515 13779
rect 7515 13745 7524 13779
rect 7472 13736 7524 13745
rect 9680 13736 9732 13788
rect 10876 13779 10928 13788
rect 10876 13745 10885 13779
rect 10885 13745 10919 13779
rect 10919 13745 10928 13779
rect 10876 13736 10928 13745
rect 7288 13711 7340 13720
rect 7288 13677 7297 13711
rect 7297 13677 7331 13711
rect 7331 13677 7340 13711
rect 7288 13668 7340 13677
rect 17960 13872 18012 13924
rect 18972 13804 19024 13856
rect 13912 13736 13964 13788
rect 14188 13779 14240 13788
rect 14188 13745 14197 13779
rect 14197 13745 14231 13779
rect 14231 13745 14240 13779
rect 14188 13736 14240 13745
rect 15936 13668 15988 13720
rect 17224 13668 17276 13720
rect 19156 13736 19208 13788
rect 20536 13668 20588 13720
rect 7196 13600 7248 13652
rect 11244 13600 11296 13652
rect 12348 13600 12400 13652
rect 15292 13600 15344 13652
rect 19248 13600 19300 13652
rect 7380 13575 7432 13584
rect 7380 13541 7389 13575
rect 7389 13541 7423 13575
rect 7423 13541 7432 13575
rect 7380 13532 7432 13541
rect 10508 13532 10560 13584
rect 16672 13532 16724 13584
rect 18144 13532 18196 13584
rect 18604 13575 18656 13584
rect 18604 13541 18613 13575
rect 18613 13541 18647 13575
rect 18647 13541 18656 13575
rect 18604 13532 18656 13541
rect 7912 13430 7964 13482
rect 7976 13430 8028 13482
rect 8040 13430 8092 13482
rect 8104 13430 8156 13482
rect 14843 13430 14895 13482
rect 14907 13430 14959 13482
rect 14971 13430 15023 13482
rect 15035 13430 15087 13482
rect 7380 13328 7432 13380
rect 11336 13328 11388 13380
rect 5540 13260 5592 13312
rect 10876 13260 10928 13312
rect 7196 13192 7248 13244
rect 8852 13235 8904 13244
rect 8852 13201 8861 13235
rect 8861 13201 8895 13235
rect 8895 13201 8904 13235
rect 8852 13192 8904 13201
rect 9404 13192 9456 13244
rect 9588 13192 9640 13244
rect 15936 13260 15988 13312
rect 17224 13328 17276 13380
rect 18696 13328 18748 13380
rect 18972 13328 19024 13380
rect 17408 13260 17460 13312
rect 20444 13303 20496 13312
rect 20444 13269 20453 13303
rect 20453 13269 20487 13303
rect 20487 13269 20496 13303
rect 20444 13260 20496 13269
rect 13176 13192 13228 13244
rect 13912 13192 13964 13244
rect 15384 13192 15436 13244
rect 16672 13235 16724 13244
rect 7656 13167 7708 13176
rect 7656 13133 7665 13167
rect 7665 13133 7699 13167
rect 7699 13133 7708 13167
rect 7656 13124 7708 13133
rect 9588 13056 9640 13108
rect 11796 13124 11848 13176
rect 13084 13167 13136 13176
rect 13084 13133 13093 13167
rect 13093 13133 13127 13167
rect 13127 13133 13136 13167
rect 13084 13124 13136 13133
rect 16672 13201 16681 13235
rect 16681 13201 16715 13235
rect 16715 13201 16724 13235
rect 16672 13192 16724 13201
rect 16948 13167 17000 13176
rect 16948 13133 16957 13167
rect 16957 13133 16991 13167
rect 16991 13133 17000 13167
rect 16948 13124 17000 13133
rect 17960 13192 18012 13244
rect 20168 13235 20220 13244
rect 20168 13201 20177 13235
rect 20177 13201 20211 13235
rect 20211 13201 20220 13235
rect 20168 13192 20220 13201
rect 18880 13124 18932 13176
rect 19156 13167 19208 13176
rect 19156 13133 19165 13167
rect 19165 13133 19199 13167
rect 19199 13133 19208 13167
rect 19156 13124 19208 13133
rect 15752 13056 15804 13108
rect 21548 13056 21600 13108
rect 12992 12988 13044 13040
rect 19248 12988 19300 13040
rect 4447 12886 4499 12938
rect 4511 12886 4563 12938
rect 4575 12886 4627 12938
rect 4639 12886 4691 12938
rect 11378 12886 11430 12938
rect 11442 12886 11494 12938
rect 11506 12886 11558 12938
rect 11570 12886 11622 12938
rect 18308 12886 18360 12938
rect 18372 12886 18424 12938
rect 18436 12886 18488 12938
rect 18500 12886 18552 12938
rect 7472 12784 7524 12836
rect 20168 12784 20220 12836
rect 15752 12759 15804 12768
rect 15752 12725 15761 12759
rect 15761 12725 15795 12759
rect 15795 12725 15804 12759
rect 15752 12716 15804 12725
rect 19156 12716 19208 12768
rect 13084 12648 13136 12700
rect 6000 12623 6052 12632
rect 6000 12589 6009 12623
rect 6009 12589 6043 12623
rect 6043 12589 6052 12623
rect 6000 12580 6052 12589
rect 7656 12580 7708 12632
rect 8668 12512 8720 12564
rect 9404 12512 9456 12564
rect 11796 12580 11848 12632
rect 16672 12623 16724 12632
rect 13176 12512 13228 12564
rect 16672 12589 16681 12623
rect 16681 12589 16715 12623
rect 16715 12589 16724 12623
rect 16672 12580 16724 12589
rect 18144 12648 18196 12700
rect 18972 12580 19024 12632
rect 19248 12623 19300 12632
rect 19248 12589 19257 12623
rect 19257 12589 19291 12623
rect 19291 12589 19300 12623
rect 19248 12580 19300 12589
rect 12624 12487 12676 12496
rect 12624 12453 12633 12487
rect 12633 12453 12667 12487
rect 12667 12453 12676 12487
rect 12624 12444 12676 12453
rect 13452 12487 13504 12496
rect 13452 12453 13461 12487
rect 13461 12453 13495 12487
rect 13495 12453 13504 12487
rect 13452 12444 13504 12453
rect 13820 12487 13872 12496
rect 13820 12453 13829 12487
rect 13829 12453 13863 12487
rect 13863 12453 13872 12487
rect 13820 12444 13872 12453
rect 16580 12512 16632 12564
rect 16948 12555 17000 12564
rect 16948 12521 16982 12555
rect 16982 12521 17000 12555
rect 16948 12512 17000 12521
rect 19064 12512 19116 12564
rect 18604 12444 18656 12496
rect 7912 12342 7964 12394
rect 7976 12342 8028 12394
rect 8040 12342 8092 12394
rect 8104 12342 8156 12394
rect 14843 12342 14895 12394
rect 14907 12342 14959 12394
rect 14971 12342 15023 12394
rect 15035 12342 15087 12394
rect 7288 12283 7340 12292
rect 7288 12249 7297 12283
rect 7297 12249 7331 12283
rect 7331 12249 7340 12283
rect 7288 12240 7340 12249
rect 7656 12240 7708 12292
rect 13084 12283 13136 12292
rect 13084 12249 13093 12283
rect 13093 12249 13127 12283
rect 13127 12249 13136 12283
rect 13084 12240 13136 12249
rect 16948 12240 17000 12292
rect 18052 12240 18104 12292
rect 19616 12283 19668 12292
rect 19616 12249 19625 12283
rect 19625 12249 19659 12283
rect 19659 12249 19668 12283
rect 19616 12240 19668 12249
rect 20720 12283 20772 12292
rect 20720 12249 20729 12283
rect 20729 12249 20763 12283
rect 20763 12249 20772 12283
rect 20720 12240 20772 12249
rect 6000 12104 6052 12156
rect 8668 12147 8720 12156
rect 8668 12113 8677 12147
rect 8677 12113 8711 12147
rect 8711 12113 8720 12147
rect 8668 12104 8720 12113
rect 12624 12172 12676 12224
rect 13452 12172 13504 12224
rect 18420 12172 18472 12224
rect 15752 12147 15804 12156
rect 15752 12113 15786 12147
rect 15786 12113 15804 12147
rect 15752 12104 15804 12113
rect 18144 12104 18196 12156
rect 19708 12104 19760 12156
rect 20536 12147 20588 12156
rect 20536 12113 20545 12147
rect 20545 12113 20579 12147
rect 20579 12113 20588 12147
rect 20536 12104 20588 12113
rect 13728 12036 13780 12088
rect 16580 11968 16632 12020
rect 18696 11968 18748 12020
rect 13912 11900 13964 11952
rect 20996 11900 21048 11952
rect 4447 11798 4499 11850
rect 4511 11798 4563 11850
rect 4575 11798 4627 11850
rect 4639 11798 4691 11850
rect 11378 11798 11430 11850
rect 11442 11798 11494 11850
rect 11506 11798 11558 11850
rect 11570 11798 11622 11850
rect 18308 11798 18360 11850
rect 18372 11798 18424 11850
rect 18436 11798 18488 11850
rect 18500 11798 18552 11850
rect 13820 11560 13872 11612
rect 15752 11560 15804 11612
rect 17960 11560 18012 11612
rect 18144 11603 18196 11612
rect 18144 11569 18153 11603
rect 18153 11569 18187 11603
rect 18187 11569 18196 11603
rect 18144 11560 18196 11569
rect 12900 11492 12952 11544
rect 18052 11492 18104 11544
rect 19708 11603 19760 11612
rect 19708 11569 19717 11603
rect 19717 11569 19751 11603
rect 19751 11569 19760 11603
rect 19708 11560 19760 11569
rect 15384 11424 15436 11476
rect 11796 11356 11848 11408
rect 15660 11399 15712 11408
rect 15660 11365 15669 11399
rect 15669 11365 15703 11399
rect 15703 11365 15712 11399
rect 15660 11356 15712 11365
rect 7912 11254 7964 11306
rect 7976 11254 8028 11306
rect 8040 11254 8092 11306
rect 8104 11254 8156 11306
rect 14843 11254 14895 11306
rect 14907 11254 14959 11306
rect 14971 11254 15023 11306
rect 15035 11254 15087 11306
rect 12808 11152 12860 11204
rect 13084 11152 13136 11204
rect 15752 11195 15804 11204
rect 11796 11084 11848 11136
rect 15752 11161 15761 11195
rect 15761 11161 15795 11195
rect 15795 11161 15804 11195
rect 15752 11152 15804 11161
rect 17776 11152 17828 11204
rect 18052 11195 18104 11204
rect 18052 11161 18061 11195
rect 18061 11161 18095 11195
rect 18095 11161 18104 11195
rect 18052 11152 18104 11161
rect 20352 11152 20404 11204
rect 12440 11016 12492 11068
rect 13084 11016 13136 11068
rect 18972 11084 19024 11136
rect 14464 11016 14516 11068
rect 17960 11016 18012 11068
rect 18144 11016 18196 11068
rect 20352 11059 20404 11068
rect 20352 11025 20361 11059
rect 20361 11025 20395 11059
rect 20395 11025 20404 11059
rect 20352 11016 20404 11025
rect 13176 10991 13228 11000
rect 13176 10957 13185 10991
rect 13185 10957 13219 10991
rect 13219 10957 13228 10991
rect 13176 10948 13228 10957
rect 14188 10880 14240 10932
rect 12808 10812 12860 10864
rect 13728 10812 13780 10864
rect 18052 10948 18104 11000
rect 18696 10991 18748 11000
rect 18696 10957 18705 10991
rect 18705 10957 18739 10991
rect 18739 10957 18748 10991
rect 18696 10948 18748 10957
rect 4447 10710 4499 10762
rect 4511 10710 4563 10762
rect 4575 10710 4627 10762
rect 4639 10710 4691 10762
rect 11378 10710 11430 10762
rect 11442 10710 11494 10762
rect 11506 10710 11558 10762
rect 11570 10710 11622 10762
rect 18308 10710 18360 10762
rect 18372 10710 18424 10762
rect 18436 10710 18488 10762
rect 18500 10710 18552 10762
rect 13176 10608 13228 10660
rect 15384 10608 15436 10660
rect 19892 10651 19944 10660
rect 19892 10617 19901 10651
rect 19901 10617 19935 10651
rect 19935 10617 19944 10651
rect 19892 10608 19944 10617
rect 14464 10540 14516 10592
rect 14188 10472 14240 10524
rect 11796 10404 11848 10456
rect 9404 10336 9456 10388
rect 16672 10404 16724 10456
rect 19248 10404 19300 10456
rect 10416 10311 10468 10320
rect 10416 10277 10425 10311
rect 10425 10277 10459 10311
rect 10459 10277 10468 10311
rect 10416 10268 10468 10277
rect 14188 10311 14240 10320
rect 14188 10277 14197 10311
rect 14197 10277 14231 10311
rect 14231 10277 14240 10311
rect 14188 10268 14240 10277
rect 15200 10268 15252 10320
rect 15936 10268 15988 10320
rect 17960 10336 18012 10388
rect 18696 10311 18748 10320
rect 18696 10277 18705 10311
rect 18705 10277 18739 10311
rect 18739 10277 18748 10311
rect 18696 10268 18748 10277
rect 7912 10166 7964 10218
rect 7976 10166 8028 10218
rect 8040 10166 8092 10218
rect 8104 10166 8156 10218
rect 14843 10166 14895 10218
rect 14907 10166 14959 10218
rect 14971 10166 15023 10218
rect 15035 10166 15087 10218
rect 14188 10064 14240 10116
rect 18052 10107 18104 10116
rect 18052 10073 18061 10107
rect 18061 10073 18095 10107
rect 18095 10073 18104 10107
rect 18052 10064 18104 10073
rect 21364 10064 21416 10116
rect 13176 9996 13228 10048
rect 14464 9928 14516 9980
rect 12808 9860 12860 9912
rect 15752 9903 15804 9912
rect 15752 9869 15761 9903
rect 15761 9869 15795 9903
rect 15795 9869 15804 9903
rect 15752 9860 15804 9869
rect 18880 9928 18932 9980
rect 20536 9971 20588 9980
rect 20536 9937 20545 9971
rect 20545 9937 20579 9971
rect 20579 9937 20588 9971
rect 20536 9928 20588 9937
rect 18052 9860 18104 9912
rect 14464 9792 14516 9844
rect 15660 9792 15712 9844
rect 17960 9792 18012 9844
rect 11152 9724 11204 9776
rect 12440 9724 12492 9776
rect 4447 9622 4499 9674
rect 4511 9622 4563 9674
rect 4575 9622 4627 9674
rect 4639 9622 4691 9674
rect 11378 9622 11430 9674
rect 11442 9622 11494 9674
rect 11506 9622 11558 9674
rect 11570 9622 11622 9674
rect 18308 9622 18360 9674
rect 18372 9622 18424 9674
rect 18436 9622 18488 9674
rect 18500 9622 18552 9674
rect 17960 9563 18012 9572
rect 17960 9529 17969 9563
rect 17969 9529 18003 9563
rect 18003 9529 18012 9563
rect 17960 9520 18012 9529
rect 12072 9452 12124 9504
rect 13544 9452 13596 9504
rect 19524 9452 19576 9504
rect 19064 9384 19116 9436
rect 11336 9316 11388 9368
rect 13360 9316 13412 9368
rect 15936 9316 15988 9368
rect 16672 9316 16724 9368
rect 14740 9248 14792 9300
rect 16580 9180 16632 9232
rect 18880 9180 18932 9232
rect 19708 9359 19760 9368
rect 19708 9325 19717 9359
rect 19717 9325 19751 9359
rect 19751 9325 19760 9359
rect 19708 9316 19760 9325
rect 7912 9078 7964 9130
rect 7976 9078 8028 9130
rect 8040 9078 8092 9130
rect 8104 9078 8156 9130
rect 14843 9078 14895 9130
rect 14907 9078 14959 9130
rect 14971 9078 15023 9130
rect 15035 9078 15087 9130
rect 14648 8976 14700 9028
rect 15936 9019 15988 9028
rect 15936 8985 15945 9019
rect 15945 8985 15979 9019
rect 15979 8985 15988 9019
rect 15936 8976 15988 8985
rect 18144 8976 18196 9028
rect 19800 8976 19852 9028
rect 21088 8976 21140 9028
rect 11336 8951 11388 8960
rect 11336 8917 11345 8951
rect 11345 8917 11379 8951
rect 11379 8917 11388 8951
rect 11336 8908 11388 8917
rect 13360 8951 13412 8960
rect 13360 8917 13369 8951
rect 13369 8917 13403 8951
rect 13403 8917 13412 8951
rect 13360 8908 13412 8917
rect 11060 8883 11112 8892
rect 11060 8849 11069 8883
rect 11069 8849 11103 8883
rect 11103 8849 11112 8883
rect 11060 8840 11112 8849
rect 13544 8840 13596 8892
rect 14740 8883 14792 8892
rect 14740 8849 14749 8883
rect 14749 8849 14783 8883
rect 14783 8849 14792 8883
rect 14740 8840 14792 8849
rect 16304 8883 16356 8892
rect 16304 8849 16313 8883
rect 16313 8849 16347 8883
rect 16347 8849 16356 8883
rect 16304 8840 16356 8849
rect 19248 8840 19300 8892
rect 20628 8840 20680 8892
rect 16396 8815 16448 8824
rect 16396 8781 16405 8815
rect 16405 8781 16439 8815
rect 16439 8781 16448 8815
rect 16396 8772 16448 8781
rect 16580 8815 16632 8824
rect 16580 8781 16589 8815
rect 16589 8781 16623 8815
rect 16623 8781 16632 8815
rect 16580 8772 16632 8781
rect 4447 8534 4499 8586
rect 4511 8534 4563 8586
rect 4575 8534 4627 8586
rect 4639 8534 4691 8586
rect 11378 8534 11430 8586
rect 11442 8534 11494 8586
rect 11506 8534 11558 8586
rect 11570 8534 11622 8586
rect 18308 8534 18360 8586
rect 18372 8534 18424 8586
rect 18436 8534 18488 8586
rect 18500 8534 18552 8586
rect 13544 8475 13596 8484
rect 13544 8441 13553 8475
rect 13553 8441 13587 8475
rect 13587 8441 13596 8475
rect 13544 8432 13596 8441
rect 16580 8432 16632 8484
rect 9772 8296 9824 8348
rect 10416 8296 10468 8348
rect 14188 8339 14240 8348
rect 14188 8305 14197 8339
rect 14197 8305 14231 8339
rect 14231 8305 14240 8339
rect 14188 8296 14240 8305
rect 11244 8228 11296 8280
rect 11152 8160 11204 8212
rect 13636 8160 13688 8212
rect 16672 8228 16724 8280
rect 12900 8092 12952 8144
rect 13912 8135 13964 8144
rect 13912 8101 13921 8135
rect 13921 8101 13955 8135
rect 13955 8101 13964 8135
rect 13912 8092 13964 8101
rect 14280 8092 14332 8144
rect 15660 8160 15712 8212
rect 7912 7990 7964 8042
rect 7976 7990 8028 8042
rect 8040 7990 8092 8042
rect 8104 7990 8156 8042
rect 14843 7990 14895 8042
rect 14907 7990 14959 8042
rect 14971 7990 15023 8042
rect 15035 7990 15087 8042
rect 11152 7931 11204 7940
rect 11152 7897 11161 7931
rect 11161 7897 11195 7931
rect 11195 7897 11204 7931
rect 11152 7888 11204 7897
rect 13912 7888 13964 7940
rect 16304 7888 16356 7940
rect 14188 7820 14240 7872
rect 15476 7820 15528 7872
rect 10048 7795 10100 7804
rect 10048 7761 10082 7795
rect 10082 7761 10100 7795
rect 10048 7752 10100 7761
rect 19248 7752 19300 7804
rect 20536 7795 20588 7804
rect 20536 7761 20545 7795
rect 20545 7761 20579 7795
rect 20579 7761 20588 7795
rect 20536 7752 20588 7761
rect 9772 7727 9824 7736
rect 9772 7693 9781 7727
rect 9781 7693 9815 7727
rect 9815 7693 9824 7727
rect 9772 7684 9824 7693
rect 12808 7684 12860 7736
rect 14280 7727 14332 7736
rect 14280 7693 14289 7727
rect 14289 7693 14323 7727
rect 14323 7693 14332 7727
rect 14280 7684 14332 7693
rect 16212 7616 16264 7668
rect 15660 7591 15712 7600
rect 15660 7557 15669 7591
rect 15669 7557 15703 7591
rect 15703 7557 15712 7591
rect 15660 7548 15712 7557
rect 4447 7446 4499 7498
rect 4511 7446 4563 7498
rect 4575 7446 4627 7498
rect 4639 7446 4691 7498
rect 11378 7446 11430 7498
rect 11442 7446 11494 7498
rect 11506 7446 11558 7498
rect 11570 7446 11622 7498
rect 18308 7446 18360 7498
rect 18372 7446 18424 7498
rect 18436 7446 18488 7498
rect 18500 7446 18552 7498
rect 11060 7344 11112 7396
rect 14188 7387 14240 7396
rect 14188 7353 14197 7387
rect 14197 7353 14231 7387
rect 14231 7353 14240 7387
rect 14188 7344 14240 7353
rect 16396 7344 16448 7396
rect 11152 7208 11204 7260
rect 12808 7251 12860 7260
rect 12808 7217 12817 7251
rect 12817 7217 12851 7251
rect 12851 7217 12860 7251
rect 12808 7208 12860 7217
rect 15660 7208 15712 7260
rect 11244 7140 11296 7192
rect 12900 7140 12952 7192
rect 16948 7183 17000 7192
rect 16948 7149 16957 7183
rect 16957 7149 16991 7183
rect 16991 7149 17000 7183
rect 16948 7140 17000 7149
rect 18052 7140 18104 7192
rect 18696 7072 18748 7124
rect 11244 7047 11296 7056
rect 11244 7013 11253 7047
rect 11253 7013 11287 7047
rect 11287 7013 11296 7047
rect 11244 7004 11296 7013
rect 7912 6902 7964 6954
rect 7976 6902 8028 6954
rect 8040 6902 8092 6954
rect 8104 6902 8156 6954
rect 14843 6902 14895 6954
rect 14907 6902 14959 6954
rect 14971 6902 15023 6954
rect 15035 6902 15087 6954
rect 13728 6732 13780 6784
rect 17960 6732 18012 6784
rect 3700 6664 3752 6716
rect 12440 6664 12492 6716
rect 16948 6664 17000 6716
rect 19248 6664 19300 6716
rect 20536 6707 20588 6716
rect 20536 6673 20545 6707
rect 20545 6673 20579 6707
rect 20579 6673 20588 6707
rect 20536 6664 20588 6673
rect 10048 6596 10100 6648
rect 12900 6596 12952 6648
rect 11244 6528 11296 6580
rect 13636 6571 13688 6580
rect 13636 6537 13645 6571
rect 13645 6537 13679 6571
rect 13679 6537 13688 6571
rect 13636 6528 13688 6537
rect 16488 6528 16540 6580
rect 9772 6460 9824 6512
rect 14556 6460 14608 6512
rect 4447 6358 4499 6410
rect 4511 6358 4563 6410
rect 4575 6358 4627 6410
rect 4639 6358 4691 6410
rect 11378 6358 11430 6410
rect 11442 6358 11494 6410
rect 11506 6358 11558 6410
rect 11570 6358 11622 6410
rect 18308 6358 18360 6410
rect 18372 6358 18424 6410
rect 18436 6358 18488 6410
rect 18500 6358 18552 6410
rect 7912 5814 7964 5866
rect 7976 5814 8028 5866
rect 8040 5814 8092 5866
rect 8104 5814 8156 5866
rect 14843 5814 14895 5866
rect 14907 5814 14959 5866
rect 14971 5814 15023 5866
rect 15035 5814 15087 5866
rect 13544 5712 13596 5764
rect 20536 5619 20588 5628
rect 20536 5585 20545 5619
rect 20545 5585 20579 5619
rect 20579 5585 20588 5619
rect 20536 5576 20588 5585
rect 4447 5270 4499 5322
rect 4511 5270 4563 5322
rect 4575 5270 4627 5322
rect 4639 5270 4691 5322
rect 11378 5270 11430 5322
rect 11442 5270 11494 5322
rect 11506 5270 11558 5322
rect 11570 5270 11622 5322
rect 18308 5270 18360 5322
rect 18372 5270 18424 5322
rect 18436 5270 18488 5322
rect 18500 5270 18552 5322
rect 7912 4726 7964 4778
rect 7976 4726 8028 4778
rect 8040 4726 8092 4778
rect 8104 4726 8156 4778
rect 14843 4726 14895 4778
rect 14907 4726 14959 4778
rect 14971 4726 15023 4778
rect 15035 4726 15087 4778
rect 13268 4624 13320 4676
rect 13820 4488 13872 4540
rect 4447 4182 4499 4234
rect 4511 4182 4563 4234
rect 4575 4182 4627 4234
rect 4639 4182 4691 4234
rect 11378 4182 11430 4234
rect 11442 4182 11494 4234
rect 11506 4182 11558 4234
rect 11570 4182 11622 4234
rect 18308 4182 18360 4234
rect 18372 4182 18424 4234
rect 18436 4182 18488 4234
rect 18500 4182 18552 4234
rect 13820 3944 13872 3996
rect 17960 3944 18012 3996
rect 13728 3876 13780 3928
rect 18052 3876 18104 3928
rect 7912 3638 7964 3690
rect 7976 3638 8028 3690
rect 8040 3638 8092 3690
rect 8104 3638 8156 3690
rect 14843 3638 14895 3690
rect 14907 3638 14959 3690
rect 14971 3638 15023 3690
rect 15035 3638 15087 3690
rect 21180 3536 21232 3588
rect 20536 3443 20588 3452
rect 20536 3409 20545 3443
rect 20545 3409 20579 3443
rect 20579 3409 20588 3443
rect 20536 3400 20588 3409
rect 4447 3094 4499 3146
rect 4511 3094 4563 3146
rect 4575 3094 4627 3146
rect 4639 3094 4691 3146
rect 11378 3094 11430 3146
rect 11442 3094 11494 3146
rect 11506 3094 11558 3146
rect 11570 3094 11622 3146
rect 18308 3094 18360 3146
rect 18372 3094 18424 3146
rect 18436 3094 18488 3146
rect 18500 3094 18552 3146
rect 7912 2550 7964 2602
rect 7976 2550 8028 2602
rect 8040 2550 8092 2602
rect 8104 2550 8156 2602
rect 14843 2550 14895 2602
rect 14907 2550 14959 2602
rect 14971 2550 15023 2602
rect 15035 2550 15087 2602
rect 15752 2448 15804 2500
rect 19248 2448 19300 2500
rect 4447 2006 4499 2058
rect 4511 2006 4563 2058
rect 4575 2006 4627 2058
rect 4639 2006 4691 2058
rect 11378 2006 11430 2058
rect 11442 2006 11494 2058
rect 11506 2006 11558 2058
rect 11570 2006 11622 2058
rect 18308 2006 18360 2058
rect 18372 2006 18424 2058
rect 18436 2006 18488 2058
rect 18500 2006 18552 2058
rect 15844 1156 15896 1208
rect 19248 1156 19300 1208
<< metal2 >>
rect 294 22376 350 22856
rect 846 22376 902 22856
rect 1398 22376 1454 22856
rect 1950 22376 2006 22856
rect 2502 22376 2558 22856
rect 3054 22376 3110 22856
rect 3606 22376 3662 22856
rect 4158 22376 4214 22856
rect 4710 22376 4766 22856
rect 5262 22376 5318 22856
rect 5814 22376 5870 22856
rect 6458 22376 6514 22856
rect 7010 22376 7066 22856
rect 7562 22376 7618 22856
rect 8114 22376 8170 22856
rect 8666 22376 8722 22856
rect 9218 22376 9274 22856
rect 9770 22376 9826 22856
rect 10322 22376 10378 22856
rect 10874 22376 10930 22856
rect 11426 22376 11482 22856
rect 12070 22376 12126 22856
rect 12622 22376 12678 22856
rect 13174 22376 13230 22856
rect 13726 22376 13782 22856
rect 14278 22376 14334 22856
rect 14830 22376 14886 22856
rect 15382 22376 15438 22856
rect 15934 22376 15990 22856
rect 16486 22376 16542 22856
rect 17038 22376 17094 22856
rect 17682 22376 17738 22856
rect 18234 22376 18290 22856
rect 18786 22376 18842 22856
rect 19062 22528 19118 22537
rect 19062 22463 19118 22472
rect 308 18554 336 22376
rect 860 18622 888 22376
rect 1412 19098 1440 22376
rect 1400 19092 1452 19098
rect 1400 19034 1452 19040
rect 848 18616 900 18622
rect 848 18558 900 18564
rect 296 18548 348 18554
rect 296 18490 348 18496
rect 1964 18282 1992 22376
rect 2516 18826 2544 22376
rect 2504 18820 2556 18826
rect 2504 18762 2556 18768
rect 1952 18276 2004 18282
rect 1952 18218 2004 18224
rect 3068 17942 3096 22376
rect 3620 19098 3648 22376
rect 3608 19092 3660 19098
rect 3608 19034 3660 19040
rect 4172 18690 4200 22376
rect 4724 20746 4752 22376
rect 4724 20718 4844 20746
rect 4421 20556 4717 20576
rect 4477 20554 4501 20556
rect 4557 20554 4581 20556
rect 4637 20554 4661 20556
rect 4499 20502 4501 20554
rect 4563 20502 4575 20554
rect 4637 20502 4639 20554
rect 4477 20500 4501 20502
rect 4557 20500 4581 20502
rect 4637 20500 4661 20502
rect 4421 20480 4717 20500
rect 4421 19468 4717 19488
rect 4477 19466 4501 19468
rect 4557 19466 4581 19468
rect 4637 19466 4661 19468
rect 4499 19414 4501 19466
rect 4563 19414 4575 19466
rect 4637 19414 4639 19466
rect 4477 19412 4501 19414
rect 4557 19412 4581 19414
rect 4637 19412 4661 19414
rect 4421 19392 4717 19412
rect 4816 18758 4844 20718
rect 4804 18752 4856 18758
rect 4804 18694 4856 18700
rect 4160 18684 4212 18690
rect 4160 18626 4212 18632
rect 4421 18380 4717 18400
rect 4477 18378 4501 18380
rect 4557 18378 4581 18380
rect 4637 18378 4661 18380
rect 4499 18326 4501 18378
rect 4563 18326 4575 18378
rect 4637 18326 4639 18378
rect 4477 18324 4501 18326
rect 4557 18324 4581 18326
rect 4637 18324 4661 18326
rect 4421 18304 4717 18324
rect 3056 17936 3108 17942
rect 3056 17878 3108 17884
rect 4068 17528 4120 17534
rect 4068 17470 4120 17476
rect 4080 17097 4108 17470
rect 4421 17292 4717 17312
rect 4477 17290 4501 17292
rect 4557 17290 4581 17292
rect 4637 17290 4661 17292
rect 4499 17238 4501 17290
rect 4563 17238 4575 17290
rect 4637 17238 4639 17290
rect 4477 17236 4501 17238
rect 4557 17236 4581 17238
rect 4637 17236 4661 17238
rect 4421 17216 4717 17236
rect 4066 17088 4122 17097
rect 4066 17023 4122 17032
rect 5276 16582 5304 22376
rect 5828 20254 5856 22376
rect 5816 20248 5868 20254
rect 5816 20190 5868 20196
rect 6276 19228 6328 19234
rect 6276 19170 6328 19176
rect 5540 18820 5592 18826
rect 5540 18762 5592 18768
rect 5264 16576 5316 16582
rect 5264 16518 5316 16524
rect 4421 16204 4717 16224
rect 4477 16202 4501 16204
rect 4557 16202 4581 16204
rect 4637 16202 4661 16204
rect 4499 16150 4501 16202
rect 4563 16150 4575 16202
rect 4637 16150 4639 16202
rect 4477 16148 4501 16150
rect 4557 16148 4581 16150
rect 4637 16148 4661 16150
rect 4421 16128 4717 16148
rect 4421 15116 4717 15136
rect 4477 15114 4501 15116
rect 4557 15114 4581 15116
rect 4637 15114 4661 15116
rect 4499 15062 4501 15114
rect 4563 15062 4575 15114
rect 4637 15062 4639 15114
rect 4477 15060 4501 15062
rect 4557 15060 4581 15062
rect 4637 15060 4661 15062
rect 4421 15040 4717 15060
rect 4421 14028 4717 14048
rect 4477 14026 4501 14028
rect 4557 14026 4581 14028
rect 4637 14026 4661 14028
rect 4499 13974 4501 14026
rect 4563 13974 4575 14026
rect 4637 13974 4639 14026
rect 4477 13972 4501 13974
rect 4557 13972 4581 13974
rect 4637 13972 4661 13974
rect 4421 13952 4717 13972
rect 5552 13318 5580 18762
rect 6288 18010 6316 19170
rect 6472 18729 6500 22376
rect 6828 19704 6880 19710
rect 6828 19646 6880 19652
rect 6840 19234 6868 19646
rect 6828 19228 6880 19234
rect 6828 19170 6880 19176
rect 6458 18720 6514 18729
rect 6458 18655 6514 18664
rect 6276 18004 6328 18010
rect 6276 17946 6328 17952
rect 6288 16990 6316 17946
rect 7024 17670 7052 22376
rect 7104 20180 7156 20186
rect 7104 20122 7156 20128
rect 7116 18826 7144 20122
rect 7196 20112 7248 20118
rect 7196 20054 7248 20060
rect 7288 20112 7340 20118
rect 7288 20054 7340 20060
rect 7208 19846 7236 20054
rect 7196 19840 7248 19846
rect 7196 19782 7248 19788
rect 7300 19166 7328 20054
rect 7472 19772 7524 19778
rect 7472 19714 7524 19720
rect 7288 19160 7340 19166
rect 7288 19102 7340 19108
rect 7104 18820 7156 18826
rect 7104 18762 7156 18768
rect 7380 18820 7432 18826
rect 7380 18762 7432 18768
rect 7104 18616 7156 18622
rect 7104 18558 7156 18564
rect 7116 18282 7144 18558
rect 7104 18276 7156 18282
rect 7104 18218 7156 18224
rect 7392 18162 7420 18762
rect 7484 18622 7512 19714
rect 7576 18826 7604 22376
rect 8128 20202 8156 22376
rect 8208 20316 8260 20322
rect 8208 20258 8260 20264
rect 7760 20174 8156 20202
rect 7760 18826 7788 20174
rect 7886 20012 8182 20032
rect 7942 20010 7966 20012
rect 8022 20010 8046 20012
rect 8102 20010 8126 20012
rect 7964 19958 7966 20010
rect 8028 19958 8040 20010
rect 8102 19958 8104 20010
rect 7942 19956 7966 19958
rect 8022 19956 8046 19958
rect 8102 19956 8126 19958
rect 7886 19936 8182 19956
rect 8220 19574 8248 20258
rect 8208 19568 8260 19574
rect 8208 19510 8260 19516
rect 8220 19166 8248 19510
rect 8208 19160 8260 19166
rect 8208 19102 8260 19108
rect 8680 19030 8708 22376
rect 9232 19914 9260 22376
rect 9220 19908 9272 19914
rect 9220 19850 9272 19856
rect 8760 19772 8812 19778
rect 8760 19714 8812 19720
rect 9220 19772 9272 19778
rect 9220 19714 9272 19720
rect 8772 19370 8800 19714
rect 9128 19704 9180 19710
rect 9128 19646 9180 19652
rect 8760 19364 8812 19370
rect 8760 19306 8812 19312
rect 9140 19166 9168 19646
rect 9128 19160 9180 19166
rect 9128 19102 9180 19108
rect 8300 19024 8352 19030
rect 8300 18966 8352 18972
rect 8668 19024 8720 19030
rect 8668 18966 8720 18972
rect 7886 18924 8182 18944
rect 7942 18922 7966 18924
rect 8022 18922 8046 18924
rect 8102 18922 8126 18924
rect 7964 18870 7966 18922
rect 8028 18870 8040 18922
rect 8102 18870 8104 18922
rect 7942 18868 7966 18870
rect 8022 18868 8046 18870
rect 8102 18868 8126 18870
rect 7886 18848 8182 18868
rect 7564 18820 7616 18826
rect 7564 18762 7616 18768
rect 7748 18820 7800 18826
rect 7748 18762 7800 18768
rect 7654 18720 7710 18729
rect 7654 18655 7710 18664
rect 7472 18616 7524 18622
rect 7472 18558 7524 18564
rect 7668 18214 7696 18655
rect 7656 18208 7708 18214
rect 7392 18134 7604 18162
rect 7656 18150 7708 18156
rect 7380 18004 7432 18010
rect 7380 17946 7432 17952
rect 7288 17936 7340 17942
rect 7288 17878 7340 17884
rect 7012 17664 7064 17670
rect 7012 17606 7064 17612
rect 7196 17596 7248 17602
rect 7196 17538 7248 17544
rect 6276 16984 6328 16990
rect 6276 16926 6328 16932
rect 7104 16984 7156 16990
rect 7104 16926 7156 16932
rect 6288 15902 6316 16926
rect 7116 16106 7144 16926
rect 7104 16100 7156 16106
rect 7104 16042 7156 16048
rect 6276 15896 6328 15902
rect 6276 15838 6328 15844
rect 6288 14814 6316 15838
rect 6276 14808 6328 14814
rect 6276 14750 6328 14756
rect 7208 13658 7236 17538
rect 7300 15562 7328 17878
rect 7392 16650 7420 17946
rect 7472 17528 7524 17534
rect 7472 17470 7524 17476
rect 7484 16990 7512 17470
rect 7472 16984 7524 16990
rect 7472 16926 7524 16932
rect 7380 16644 7432 16650
rect 7380 16586 7432 16592
rect 7288 15556 7340 15562
rect 7288 15498 7340 15504
rect 7576 15494 7604 18134
rect 7656 18072 7708 18078
rect 7656 18014 7708 18020
rect 7746 18040 7802 18049
rect 7668 17194 7696 18014
rect 7746 17975 7802 17984
rect 7760 17942 7788 17975
rect 8312 17942 8340 18966
rect 8576 18752 8628 18758
rect 8576 18694 8628 18700
rect 8392 18548 8444 18554
rect 8392 18490 8444 18496
rect 8404 18078 8432 18490
rect 8392 18072 8444 18078
rect 8392 18014 8444 18020
rect 8588 18010 8616 18694
rect 8944 18684 8996 18690
rect 8944 18626 8996 18632
rect 8576 18004 8628 18010
rect 8576 17946 8628 17952
rect 7748 17936 7800 17942
rect 7748 17878 7800 17884
rect 8208 17936 8260 17942
rect 8208 17878 8260 17884
rect 8300 17936 8352 17942
rect 8300 17878 8352 17884
rect 7886 17836 8182 17856
rect 7942 17834 7966 17836
rect 8022 17834 8046 17836
rect 8102 17834 8126 17836
rect 7964 17782 7966 17834
rect 8028 17782 8040 17834
rect 8102 17782 8104 17834
rect 7942 17780 7966 17782
rect 8022 17780 8046 17782
rect 8102 17780 8126 17782
rect 7886 17760 8182 17780
rect 8220 17738 8248 17878
rect 8208 17732 8260 17738
rect 8208 17674 8260 17680
rect 8956 17602 8984 18626
rect 8944 17596 8996 17602
rect 8944 17538 8996 17544
rect 7656 17188 7708 17194
rect 7656 17130 7708 17136
rect 9140 16990 9168 19102
rect 9232 18622 9260 19714
rect 9784 19137 9812 22376
rect 9770 19128 9826 19137
rect 9496 19092 9548 19098
rect 9770 19063 9826 19072
rect 10140 19092 10192 19098
rect 9496 19034 9548 19040
rect 10140 19034 10192 19040
rect 9220 18616 9272 18622
rect 9220 18558 9272 18564
rect 9508 17738 9536 19034
rect 10152 18826 10180 19034
rect 10140 18820 10192 18826
rect 10140 18762 10192 18768
rect 10230 18720 10286 18729
rect 10230 18655 10286 18664
rect 9680 18276 9732 18282
rect 9680 18218 9732 18224
rect 9496 17732 9548 17738
rect 9496 17674 9548 17680
rect 9588 17596 9640 17602
rect 9588 17538 9640 17544
rect 9128 16984 9180 16990
rect 9128 16926 9180 16932
rect 7886 16748 8182 16768
rect 7942 16746 7966 16748
rect 8022 16746 8046 16748
rect 8102 16746 8126 16748
rect 7964 16694 7966 16746
rect 8028 16694 8040 16746
rect 8102 16694 8104 16746
rect 7942 16692 7966 16694
rect 8022 16692 8046 16694
rect 8102 16692 8126 16694
rect 7886 16672 8182 16692
rect 9140 16446 9168 16926
rect 9128 16440 9180 16446
rect 9128 16382 9180 16388
rect 8392 16304 8444 16310
rect 8392 16246 8444 16252
rect 7886 15660 8182 15680
rect 7942 15658 7966 15660
rect 8022 15658 8046 15660
rect 8102 15658 8126 15660
rect 7964 15606 7966 15658
rect 8028 15606 8040 15658
rect 8102 15606 8104 15658
rect 7942 15604 7966 15606
rect 8022 15604 8046 15606
rect 8102 15604 8126 15606
rect 7886 15584 8182 15604
rect 7564 15488 7616 15494
rect 7564 15430 7616 15436
rect 8404 15358 8432 16246
rect 9600 15494 9628 17538
rect 9588 15488 9640 15494
rect 9588 15430 9640 15436
rect 8668 15420 8720 15426
rect 8668 15362 8720 15368
rect 7472 15352 7524 15358
rect 7472 15294 7524 15300
rect 8392 15352 8444 15358
rect 8392 15294 8444 15300
rect 7484 14746 7512 15294
rect 7748 15216 7800 15222
rect 7748 15158 7800 15164
rect 7472 14740 7524 14746
rect 7472 14682 7524 14688
rect 7760 14678 7788 15158
rect 8404 14814 8432 15294
rect 8680 14950 8708 15362
rect 8668 14944 8720 14950
rect 8668 14886 8720 14892
rect 8392 14808 8444 14814
rect 8392 14750 8444 14756
rect 8208 14740 8260 14746
rect 8208 14682 8260 14688
rect 7748 14672 7800 14678
rect 7748 14614 7800 14620
rect 7886 14572 8182 14592
rect 7942 14570 7966 14572
rect 8022 14570 8046 14572
rect 8102 14570 8126 14572
rect 7964 14518 7966 14570
rect 8028 14518 8040 14570
rect 8102 14518 8104 14570
rect 7942 14516 7966 14518
rect 8022 14516 8046 14518
rect 8102 14516 8126 14518
rect 7886 14496 8182 14516
rect 8220 14474 8248 14682
rect 8208 14468 8260 14474
rect 8208 14410 8260 14416
rect 8404 14338 8432 14750
rect 7472 14332 7524 14338
rect 7472 14274 7524 14280
rect 8392 14332 8444 14338
rect 8392 14274 8444 14280
rect 7484 13794 7512 14274
rect 8852 13856 8904 13862
rect 8852 13798 8904 13804
rect 7472 13788 7524 13794
rect 7472 13730 7524 13736
rect 7288 13720 7340 13726
rect 7288 13662 7340 13668
rect 7196 13652 7248 13658
rect 7196 13594 7248 13600
rect 5540 13312 5592 13318
rect 5540 13254 5592 13260
rect 7208 13250 7236 13594
rect 7196 13244 7248 13250
rect 7196 13186 7248 13192
rect 4421 12940 4717 12960
rect 4477 12938 4501 12940
rect 4557 12938 4581 12940
rect 4637 12938 4661 12940
rect 4499 12886 4501 12938
rect 4563 12886 4575 12938
rect 4637 12886 4639 12938
rect 4477 12884 4501 12886
rect 4557 12884 4581 12886
rect 4637 12884 4661 12886
rect 4421 12864 4717 12884
rect 6000 12632 6052 12638
rect 6000 12574 6052 12580
rect 6012 12162 6040 12574
rect 7300 12298 7328 13662
rect 7380 13584 7432 13590
rect 7380 13526 7432 13532
rect 7392 13386 7420 13526
rect 7380 13380 7432 13386
rect 7380 13322 7432 13328
rect 7484 12842 7512 13730
rect 7886 13484 8182 13504
rect 7942 13482 7966 13484
rect 8022 13482 8046 13484
rect 8102 13482 8126 13484
rect 7964 13430 7966 13482
rect 8028 13430 8040 13482
rect 8102 13430 8104 13482
rect 7942 13428 7966 13430
rect 8022 13428 8046 13430
rect 8102 13428 8126 13430
rect 7886 13408 8182 13428
rect 8864 13250 8892 13798
rect 9692 13794 9720 18218
rect 10244 18214 10272 18655
rect 10336 18214 10364 22376
rect 10508 19568 10560 19574
rect 10508 19510 10560 19516
rect 10520 19166 10548 19510
rect 10508 19160 10560 19166
rect 10508 19102 10560 19108
rect 10784 19160 10836 19166
rect 10784 19102 10836 19108
rect 10796 18622 10824 19102
rect 10784 18616 10836 18622
rect 10784 18558 10836 18564
rect 10232 18208 10284 18214
rect 10232 18150 10284 18156
rect 10324 18208 10376 18214
rect 10324 18150 10376 18156
rect 9864 18140 9916 18146
rect 9864 18082 9916 18088
rect 9772 17528 9824 17534
rect 9772 17470 9824 17476
rect 9784 16582 9812 17470
rect 9876 17466 9904 18082
rect 10888 18078 10916 22376
rect 11440 20746 11468 22376
rect 11440 20718 11744 20746
rect 11352 20556 11648 20576
rect 11408 20554 11432 20556
rect 11488 20554 11512 20556
rect 11568 20554 11592 20556
rect 11430 20502 11432 20554
rect 11494 20502 11506 20554
rect 11568 20502 11570 20554
rect 11408 20500 11432 20502
rect 11488 20500 11512 20502
rect 11568 20500 11592 20502
rect 11352 20480 11648 20500
rect 11428 20248 11480 20254
rect 11428 20190 11480 20196
rect 11152 20112 11204 20118
rect 11152 20054 11204 20060
rect 11060 19704 11112 19710
rect 11060 19646 11112 19652
rect 10968 19024 11020 19030
rect 10968 18966 11020 18972
rect 10980 18706 11008 18966
rect 11072 18826 11100 19646
rect 11060 18820 11112 18826
rect 11060 18762 11112 18768
rect 10980 18678 11100 18706
rect 11072 18622 11100 18678
rect 11060 18616 11112 18622
rect 11060 18558 11112 18564
rect 10692 18072 10744 18078
rect 10692 18014 10744 18020
rect 10876 18072 10928 18078
rect 10876 18014 10928 18020
rect 10704 17618 10732 18014
rect 11164 17942 11192 20054
rect 11440 19681 11468 20190
rect 11426 19672 11482 19681
rect 11426 19607 11482 19616
rect 11352 19468 11648 19488
rect 11408 19466 11432 19468
rect 11488 19466 11512 19468
rect 11568 19466 11592 19468
rect 11430 19414 11432 19466
rect 11494 19414 11506 19466
rect 11568 19414 11570 19466
rect 11408 19412 11432 19414
rect 11488 19412 11512 19414
rect 11568 19412 11592 19414
rect 11352 19392 11648 19412
rect 11716 18826 11744 20718
rect 11704 18820 11756 18826
rect 11704 18762 11756 18768
rect 11244 18480 11296 18486
rect 11244 18422 11296 18428
rect 11256 17942 11284 18422
rect 11352 18380 11648 18400
rect 11408 18378 11432 18380
rect 11488 18378 11512 18380
rect 11568 18378 11592 18380
rect 11430 18326 11432 18378
rect 11494 18326 11506 18378
rect 11568 18326 11570 18378
rect 11408 18324 11432 18326
rect 11488 18324 11512 18326
rect 11568 18324 11592 18326
rect 11352 18304 11648 18324
rect 11704 18208 11756 18214
rect 11704 18150 11756 18156
rect 10784 17936 10836 17942
rect 11152 17936 11204 17942
rect 10836 17884 11100 17890
rect 10784 17878 11100 17884
rect 11152 17878 11204 17884
rect 11244 17936 11296 17942
rect 11244 17878 11296 17884
rect 10796 17862 11100 17878
rect 11072 17754 11100 17862
rect 11072 17726 11192 17754
rect 10704 17590 11100 17618
rect 9864 17460 9916 17466
rect 9864 17402 9916 17408
rect 10508 17392 10560 17398
rect 10508 17334 10560 17340
rect 9772 16576 9824 16582
rect 9772 16518 9824 16524
rect 9784 15562 9812 16518
rect 10520 15766 10548 17334
rect 10600 16916 10652 16922
rect 10600 16858 10652 16864
rect 10612 16650 10640 16858
rect 10600 16644 10652 16650
rect 10600 16586 10652 16592
rect 10612 15970 10640 16586
rect 11072 16530 11100 17590
rect 10980 16502 11100 16530
rect 10600 15964 10652 15970
rect 10600 15906 10652 15912
rect 10508 15760 10560 15766
rect 10508 15702 10560 15708
rect 10980 15714 11008 16502
rect 11060 16440 11112 16446
rect 11060 16382 11112 16388
rect 11072 15902 11100 16382
rect 11060 15896 11112 15902
rect 11060 15838 11112 15844
rect 10980 15686 11100 15714
rect 9772 15556 9824 15562
rect 9772 15498 9824 15504
rect 10508 15420 10560 15426
rect 10508 15362 10560 15368
rect 9680 13788 9732 13794
rect 9680 13730 9732 13736
rect 10520 13590 10548 15362
rect 10600 15352 10652 15358
rect 10600 15294 10652 15300
rect 10612 14814 10640 15294
rect 10600 14808 10652 14814
rect 10600 14750 10652 14756
rect 11072 14762 11100 15686
rect 11164 14882 11192 17726
rect 11352 17292 11648 17312
rect 11408 17290 11432 17292
rect 11488 17290 11512 17292
rect 11568 17290 11592 17292
rect 11430 17238 11432 17290
rect 11494 17238 11506 17290
rect 11568 17238 11570 17290
rect 11408 17236 11432 17238
rect 11488 17236 11512 17238
rect 11568 17236 11592 17238
rect 11352 17216 11648 17236
rect 11244 16984 11296 16990
rect 11244 16926 11296 16932
rect 11256 16514 11284 16926
rect 11716 16650 11744 18150
rect 11704 16644 11756 16650
rect 11704 16586 11756 16592
rect 11244 16508 11296 16514
rect 11244 16450 11296 16456
rect 11256 15562 11284 16450
rect 11352 16204 11648 16224
rect 11408 16202 11432 16204
rect 11488 16202 11512 16204
rect 11568 16202 11592 16204
rect 11430 16150 11432 16202
rect 11494 16150 11506 16202
rect 11568 16150 11570 16202
rect 11408 16148 11432 16150
rect 11488 16148 11512 16150
rect 11568 16148 11592 16150
rect 11352 16128 11648 16148
rect 11244 15556 11296 15562
rect 11244 15498 11296 15504
rect 11352 15116 11648 15136
rect 11408 15114 11432 15116
rect 11488 15114 11512 15116
rect 11568 15114 11592 15116
rect 11430 15062 11432 15114
rect 11494 15062 11506 15114
rect 11568 15062 11570 15114
rect 11408 15060 11432 15062
rect 11488 15060 11512 15062
rect 11568 15060 11592 15062
rect 11352 15040 11648 15060
rect 11152 14876 11204 14882
rect 11152 14818 11204 14824
rect 11888 14876 11940 14882
rect 11888 14818 11940 14824
rect 11072 14734 11192 14762
rect 10876 14128 10928 14134
rect 10876 14070 10928 14076
rect 10888 13794 10916 14070
rect 10876 13788 10928 13794
rect 10876 13730 10928 13736
rect 10508 13584 10560 13590
rect 10508 13526 10560 13532
rect 10888 13318 10916 13730
rect 10876 13312 10928 13318
rect 9416 13250 9628 13266
rect 10876 13254 10928 13260
rect 8852 13244 8904 13250
rect 8852 13186 8904 13192
rect 9404 13244 9640 13250
rect 9456 13238 9588 13244
rect 9404 13186 9456 13192
rect 9588 13186 9640 13192
rect 7656 13176 7708 13182
rect 7656 13118 7708 13124
rect 9402 13144 9458 13153
rect 7472 12836 7524 12842
rect 7472 12778 7524 12784
rect 7668 12638 7696 13118
rect 9402 13079 9458 13088
rect 9586 13144 9642 13153
rect 9586 13079 9588 13088
rect 7656 12632 7708 12638
rect 7656 12574 7708 12580
rect 7668 12298 7696 12574
rect 9416 12570 9444 13079
rect 9640 13079 9642 13088
rect 9588 13050 9640 13056
rect 8668 12564 8720 12570
rect 8668 12506 8720 12512
rect 9404 12564 9456 12570
rect 9404 12506 9456 12512
rect 7886 12396 8182 12416
rect 7942 12394 7966 12396
rect 8022 12394 8046 12396
rect 8102 12394 8126 12396
rect 7964 12342 7966 12394
rect 8028 12342 8040 12394
rect 8102 12342 8104 12394
rect 7942 12340 7966 12342
rect 8022 12340 8046 12342
rect 8102 12340 8126 12342
rect 7886 12320 8182 12340
rect 7288 12292 7340 12298
rect 7288 12234 7340 12240
rect 7656 12292 7708 12298
rect 7656 12234 7708 12240
rect 8680 12162 8708 12506
rect 6000 12156 6052 12162
rect 6000 12098 6052 12104
rect 8668 12156 8720 12162
rect 8668 12098 8720 12104
rect 4421 11852 4717 11872
rect 4477 11850 4501 11852
rect 4557 11850 4581 11852
rect 4637 11850 4661 11852
rect 4499 11798 4501 11850
rect 4563 11798 4575 11850
rect 4637 11798 4639 11850
rect 4477 11796 4501 11798
rect 4557 11796 4581 11798
rect 4637 11796 4661 11798
rect 4421 11776 4717 11796
rect 7886 11308 8182 11328
rect 7942 11306 7966 11308
rect 8022 11306 8046 11308
rect 8102 11306 8126 11308
rect 7964 11254 7966 11306
rect 8028 11254 8040 11306
rect 8102 11254 8104 11306
rect 7942 11252 7966 11254
rect 8022 11252 8046 11254
rect 8102 11252 8126 11254
rect 7886 11232 8182 11252
rect 4421 10764 4717 10784
rect 4477 10762 4501 10764
rect 4557 10762 4581 10764
rect 4637 10762 4661 10764
rect 4499 10710 4501 10762
rect 4563 10710 4575 10762
rect 4637 10710 4639 10762
rect 4477 10708 4501 10710
rect 4557 10708 4581 10710
rect 4637 10708 4661 10710
rect 4421 10688 4717 10708
rect 9416 10394 9444 12506
rect 9404 10388 9456 10394
rect 9404 10330 9456 10336
rect 10416 10320 10468 10326
rect 10416 10262 10468 10268
rect 7886 10220 8182 10240
rect 7942 10218 7966 10220
rect 8022 10218 8046 10220
rect 8102 10218 8126 10220
rect 7964 10166 7966 10218
rect 8028 10166 8040 10218
rect 8102 10166 8104 10218
rect 7942 10164 7966 10166
rect 8022 10164 8046 10166
rect 8102 10164 8126 10166
rect 7886 10144 8182 10164
rect 4421 9676 4717 9696
rect 4477 9674 4501 9676
rect 4557 9674 4581 9676
rect 4637 9674 4661 9676
rect 4499 9622 4501 9674
rect 4563 9622 4575 9674
rect 4637 9622 4639 9674
rect 4477 9620 4501 9622
rect 4557 9620 4581 9622
rect 4637 9620 4661 9622
rect 4421 9600 4717 9620
rect 7886 9132 8182 9152
rect 7942 9130 7966 9132
rect 8022 9130 8046 9132
rect 8102 9130 8126 9132
rect 7964 9078 7966 9130
rect 8028 9078 8040 9130
rect 8102 9078 8104 9130
rect 7942 9076 7966 9078
rect 8022 9076 8046 9078
rect 8102 9076 8126 9078
rect 7886 9056 8182 9076
rect 4421 8588 4717 8608
rect 4477 8586 4501 8588
rect 4557 8586 4581 8588
rect 4637 8586 4661 8588
rect 4499 8534 4501 8586
rect 4563 8534 4575 8586
rect 4637 8534 4639 8586
rect 4477 8532 4501 8534
rect 4557 8532 4581 8534
rect 4637 8532 4661 8534
rect 4421 8512 4717 8532
rect 10428 8354 10456 10262
rect 11164 9782 11192 14734
rect 11244 14672 11296 14678
rect 11244 14614 11296 14620
rect 11256 13658 11284 14614
rect 11900 14338 11928 14818
rect 11888 14332 11940 14338
rect 11888 14274 11940 14280
rect 11352 14028 11648 14048
rect 11408 14026 11432 14028
rect 11488 14026 11512 14028
rect 11568 14026 11592 14028
rect 11430 13974 11432 14026
rect 11494 13974 11506 14026
rect 11568 13974 11570 14026
rect 11408 13972 11432 13974
rect 11488 13972 11512 13974
rect 11568 13972 11592 13974
rect 11352 13952 11648 13972
rect 11336 13856 11388 13862
rect 11336 13798 11388 13804
rect 11244 13652 11296 13658
rect 11244 13594 11296 13600
rect 11348 13386 11376 13798
rect 11336 13380 11388 13386
rect 11336 13322 11388 13328
rect 11796 13176 11848 13182
rect 11796 13118 11848 13124
rect 11352 12940 11648 12960
rect 11408 12938 11432 12940
rect 11488 12938 11512 12940
rect 11568 12938 11592 12940
rect 11430 12886 11432 12938
rect 11494 12886 11506 12938
rect 11568 12886 11570 12938
rect 11408 12884 11432 12886
rect 11488 12884 11512 12886
rect 11568 12884 11592 12886
rect 11352 12864 11648 12884
rect 11808 12638 11836 13118
rect 11796 12632 11848 12638
rect 11796 12574 11848 12580
rect 11352 11852 11648 11872
rect 11408 11850 11432 11852
rect 11488 11850 11512 11852
rect 11568 11850 11592 11852
rect 11430 11798 11432 11850
rect 11494 11798 11506 11850
rect 11568 11798 11570 11850
rect 11408 11796 11432 11798
rect 11488 11796 11512 11798
rect 11568 11796 11592 11798
rect 11352 11776 11648 11796
rect 11796 11408 11848 11414
rect 11796 11350 11848 11356
rect 11808 11142 11836 11350
rect 11796 11136 11848 11142
rect 11796 11078 11848 11084
rect 11352 10764 11648 10784
rect 11408 10762 11432 10764
rect 11488 10762 11512 10764
rect 11568 10762 11592 10764
rect 11430 10710 11432 10762
rect 11494 10710 11506 10762
rect 11568 10710 11570 10762
rect 11408 10708 11432 10710
rect 11488 10708 11512 10710
rect 11568 10708 11592 10710
rect 11352 10688 11648 10708
rect 11808 10462 11836 11078
rect 11796 10456 11848 10462
rect 11796 10398 11848 10404
rect 11152 9776 11204 9782
rect 11152 9718 11204 9724
rect 11352 9676 11648 9696
rect 11408 9674 11432 9676
rect 11488 9674 11512 9676
rect 11568 9674 11592 9676
rect 11430 9622 11432 9674
rect 11494 9622 11506 9674
rect 11568 9622 11570 9674
rect 11408 9620 11432 9622
rect 11488 9620 11512 9622
rect 11568 9620 11592 9622
rect 11352 9600 11648 9620
rect 12084 9510 12112 22376
rect 12348 19840 12400 19846
rect 12346 19808 12348 19817
rect 12400 19808 12402 19817
rect 12346 19743 12402 19752
rect 12532 19704 12584 19710
rect 12532 19646 12584 19652
rect 12544 19370 12572 19646
rect 12532 19364 12584 19370
rect 12532 19306 12584 19312
rect 12544 19250 12572 19306
rect 12452 19222 12572 19250
rect 12348 19024 12400 19030
rect 12348 18966 12400 18972
rect 12360 18826 12388 18966
rect 12348 18820 12400 18826
rect 12348 18762 12400 18768
rect 12452 18162 12480 19222
rect 12532 18480 12584 18486
rect 12532 18422 12584 18428
rect 12544 18282 12572 18422
rect 12636 18282 12664 22376
rect 13188 20474 13216 22376
rect 13188 20446 13584 20474
rect 13004 20322 13308 20338
rect 13004 20316 13320 20322
rect 13004 20310 13268 20316
rect 13004 19778 13032 20310
rect 13268 20258 13320 20264
rect 13084 20248 13136 20254
rect 13452 20248 13504 20254
rect 13136 20196 13452 20202
rect 13084 20190 13504 20196
rect 13096 20174 13492 20190
rect 12992 19772 13044 19778
rect 12992 19714 13044 19720
rect 13268 19772 13320 19778
rect 13268 19714 13320 19720
rect 13280 19370 13308 19714
rect 13268 19364 13320 19370
rect 13268 19306 13320 19312
rect 12900 19296 12952 19302
rect 12900 19238 12952 19244
rect 12808 19024 12860 19030
rect 12808 18966 12860 18972
rect 12532 18276 12584 18282
rect 12532 18218 12584 18224
rect 12624 18276 12676 18282
rect 12624 18218 12676 18224
rect 12452 18134 12572 18162
rect 12440 17392 12492 17398
rect 12440 17334 12492 17340
rect 12452 15970 12480 17334
rect 12544 16854 12572 18134
rect 12716 17732 12768 17738
rect 12716 17674 12768 17680
rect 12532 16848 12584 16854
rect 12532 16790 12584 16796
rect 12544 16514 12572 16790
rect 12532 16508 12584 16514
rect 12532 16450 12584 16456
rect 12440 15964 12492 15970
rect 12440 15906 12492 15912
rect 12544 14882 12572 16450
rect 12624 16032 12676 16038
rect 12624 15974 12676 15980
rect 12636 15562 12664 15974
rect 12728 15902 12756 17674
rect 12716 15896 12768 15902
rect 12716 15838 12768 15844
rect 12624 15556 12676 15562
rect 12624 15498 12676 15504
rect 12532 14876 12584 14882
rect 12532 14818 12584 14824
rect 12348 13652 12400 13658
rect 12348 13594 12400 13600
rect 12360 13266 12388 13594
rect 12360 13238 12480 13266
rect 12452 11074 12480 13238
rect 12624 12496 12676 12502
rect 12624 12438 12676 12444
rect 12636 12230 12664 12438
rect 12624 12224 12676 12230
rect 12624 12166 12676 12172
rect 12820 11210 12848 18966
rect 12912 18826 12940 19238
rect 12992 19092 13044 19098
rect 12992 19034 13044 19040
rect 12900 18820 12952 18826
rect 12900 18762 12952 18768
rect 13004 18622 13032 19034
rect 13084 18752 13136 18758
rect 13084 18694 13136 18700
rect 12992 18616 13044 18622
rect 12992 18558 13044 18564
rect 13096 17738 13124 18694
rect 13176 18684 13228 18690
rect 13176 18626 13228 18632
rect 13084 17732 13136 17738
rect 13084 17674 13136 17680
rect 13188 17602 13216 18626
rect 13268 18276 13320 18282
rect 13268 18218 13320 18224
rect 13176 17596 13228 17602
rect 13176 17538 13228 17544
rect 12992 17528 13044 17534
rect 12992 17470 13044 17476
rect 13004 17126 13032 17470
rect 12992 17120 13044 17126
rect 12992 17062 13044 17068
rect 13004 16514 13032 17062
rect 12992 16508 13044 16514
rect 12992 16450 13044 16456
rect 13084 15420 13136 15426
rect 13084 15362 13136 15368
rect 13096 13930 13124 15362
rect 13084 13924 13136 13930
rect 13084 13866 13136 13872
rect 13096 13810 13124 13866
rect 12912 13782 13124 13810
rect 12912 11550 12940 13782
rect 13188 13250 13216 17538
rect 13176 13244 13228 13250
rect 13176 13186 13228 13192
rect 13084 13176 13136 13182
rect 13084 13118 13136 13124
rect 12992 13040 13044 13046
rect 12992 12982 13044 12988
rect 13004 12586 13032 12982
rect 13096 12706 13124 13118
rect 13084 12700 13136 12706
rect 13084 12642 13136 12648
rect 13004 12558 13124 12586
rect 13188 12570 13216 13186
rect 13096 12298 13124 12558
rect 13176 12564 13228 12570
rect 13176 12506 13228 12512
rect 13084 12292 13136 12298
rect 13084 12234 13136 12240
rect 12900 11544 12952 11550
rect 12900 11486 12952 11492
rect 12808 11204 12860 11210
rect 12808 11146 12860 11152
rect 13084 11204 13136 11210
rect 13084 11146 13136 11152
rect 13096 11074 13124 11146
rect 12440 11068 12492 11074
rect 12440 11010 12492 11016
rect 13084 11068 13136 11074
rect 13084 11010 13136 11016
rect 13176 11000 13228 11006
rect 13176 10942 13228 10948
rect 12808 10864 12860 10870
rect 12808 10806 12860 10812
rect 12820 9918 12848 10806
rect 13188 10666 13216 10942
rect 13176 10660 13228 10666
rect 13176 10602 13228 10608
rect 13188 10054 13216 10602
rect 13176 10048 13228 10054
rect 13176 9990 13228 9996
rect 12808 9912 12860 9918
rect 12808 9854 12860 9860
rect 12440 9776 12492 9782
rect 12440 9718 12492 9724
rect 12072 9504 12124 9510
rect 12072 9446 12124 9452
rect 11336 9368 11388 9374
rect 11336 9310 11388 9316
rect 11348 8966 11376 9310
rect 11336 8960 11388 8966
rect 11336 8902 11388 8908
rect 11060 8892 11112 8898
rect 11060 8834 11112 8840
rect 9772 8348 9824 8354
rect 9772 8290 9824 8296
rect 10416 8348 10468 8354
rect 10416 8290 10468 8296
rect 7886 8044 8182 8064
rect 7942 8042 7966 8044
rect 8022 8042 8046 8044
rect 8102 8042 8126 8044
rect 7964 7990 7966 8042
rect 8028 7990 8040 8042
rect 8102 7990 8104 8042
rect 7942 7988 7966 7990
rect 8022 7988 8046 7990
rect 8102 7988 8126 7990
rect 7886 7968 8182 7988
rect 9784 7742 9812 8290
rect 10048 7804 10100 7810
rect 10048 7746 10100 7752
rect 9772 7736 9824 7742
rect 9772 7678 9824 7684
rect 4421 7500 4717 7520
rect 4477 7498 4501 7500
rect 4557 7498 4581 7500
rect 4637 7498 4661 7500
rect 4499 7446 4501 7498
rect 4563 7446 4575 7498
rect 4637 7446 4639 7498
rect 4477 7444 4501 7446
rect 4557 7444 4581 7446
rect 4637 7444 4661 7446
rect 4421 7424 4717 7444
rect 7886 6956 8182 6976
rect 7942 6954 7966 6956
rect 8022 6954 8046 6956
rect 8102 6954 8126 6956
rect 7964 6902 7966 6954
rect 8028 6902 8040 6954
rect 8102 6902 8104 6954
rect 7942 6900 7966 6902
rect 8022 6900 8046 6902
rect 8102 6900 8126 6902
rect 7886 6880 8182 6900
rect 3700 6716 3752 6722
rect 3700 6658 3752 6664
rect 3712 5673 3740 6658
rect 9784 6518 9812 7678
rect 10060 6654 10088 7746
rect 11072 7402 11100 8834
rect 11352 8588 11648 8608
rect 11408 8586 11432 8588
rect 11488 8586 11512 8588
rect 11568 8586 11592 8588
rect 11430 8534 11432 8586
rect 11494 8534 11506 8586
rect 11568 8534 11570 8586
rect 11408 8532 11432 8534
rect 11488 8532 11512 8534
rect 11568 8532 11592 8534
rect 11352 8512 11648 8532
rect 11244 8280 11296 8286
rect 11244 8222 11296 8228
rect 11152 8212 11204 8218
rect 11152 8154 11204 8160
rect 11164 7946 11192 8154
rect 11152 7940 11204 7946
rect 11152 7882 11204 7888
rect 11060 7396 11112 7402
rect 11060 7338 11112 7344
rect 11164 7266 11192 7882
rect 11152 7260 11204 7266
rect 11152 7202 11204 7208
rect 11256 7198 11284 8222
rect 11352 7500 11648 7520
rect 11408 7498 11432 7500
rect 11488 7498 11512 7500
rect 11568 7498 11592 7500
rect 11430 7446 11432 7498
rect 11494 7446 11506 7498
rect 11568 7446 11570 7498
rect 11408 7444 11432 7446
rect 11488 7444 11512 7446
rect 11568 7444 11592 7446
rect 11352 7424 11648 7444
rect 11244 7192 11296 7198
rect 11244 7134 11296 7140
rect 11244 7056 11296 7062
rect 11244 6998 11296 7004
rect 10048 6648 10100 6654
rect 10048 6590 10100 6596
rect 11256 6586 11284 6998
rect 12452 6722 12480 9718
rect 12820 7742 12848 9854
rect 12900 8144 12952 8150
rect 12900 8086 12952 8092
rect 12808 7736 12860 7742
rect 12808 7678 12860 7684
rect 12820 7266 12848 7678
rect 12808 7260 12860 7266
rect 12808 7202 12860 7208
rect 12912 7198 12940 8086
rect 12900 7192 12952 7198
rect 12900 7134 12952 7140
rect 12440 6716 12492 6722
rect 12440 6658 12492 6664
rect 12912 6654 12940 7134
rect 12900 6648 12952 6654
rect 12900 6590 12952 6596
rect 11244 6580 11296 6586
rect 11244 6522 11296 6528
rect 9772 6512 9824 6518
rect 9772 6454 9824 6460
rect 4421 6412 4717 6432
rect 4477 6410 4501 6412
rect 4557 6410 4581 6412
rect 4637 6410 4661 6412
rect 4499 6358 4501 6410
rect 4563 6358 4575 6410
rect 4637 6358 4639 6410
rect 4477 6356 4501 6358
rect 4557 6356 4581 6358
rect 4637 6356 4661 6358
rect 4421 6336 4717 6356
rect 11352 6412 11648 6432
rect 11408 6410 11432 6412
rect 11488 6410 11512 6412
rect 11568 6410 11592 6412
rect 11430 6358 11432 6410
rect 11494 6358 11506 6410
rect 11568 6358 11570 6410
rect 11408 6356 11432 6358
rect 11488 6356 11512 6358
rect 11568 6356 11592 6358
rect 11352 6336 11648 6356
rect 7886 5868 8182 5888
rect 7942 5866 7966 5868
rect 8022 5866 8046 5868
rect 8102 5866 8126 5868
rect 7964 5814 7966 5866
rect 8028 5814 8040 5866
rect 8102 5814 8104 5866
rect 7942 5812 7966 5814
rect 8022 5812 8046 5814
rect 8102 5812 8126 5814
rect 7886 5792 8182 5812
rect 3698 5664 3754 5673
rect 3698 5599 3754 5608
rect 4421 5324 4717 5344
rect 4477 5322 4501 5324
rect 4557 5322 4581 5324
rect 4637 5322 4661 5324
rect 4499 5270 4501 5322
rect 4563 5270 4575 5322
rect 4637 5270 4639 5322
rect 4477 5268 4501 5270
rect 4557 5268 4581 5270
rect 4637 5268 4661 5270
rect 4421 5248 4717 5268
rect 11352 5324 11648 5344
rect 11408 5322 11432 5324
rect 11488 5322 11512 5324
rect 11568 5322 11592 5324
rect 11430 5270 11432 5322
rect 11494 5270 11506 5322
rect 11568 5270 11570 5322
rect 11408 5268 11432 5270
rect 11488 5268 11512 5270
rect 11568 5268 11592 5270
rect 11352 5248 11648 5268
rect 7886 4780 8182 4800
rect 7942 4778 7966 4780
rect 8022 4778 8046 4780
rect 8102 4778 8126 4780
rect 7964 4726 7966 4778
rect 8028 4726 8040 4778
rect 8102 4726 8104 4778
rect 7942 4724 7966 4726
rect 8022 4724 8046 4726
rect 8102 4724 8126 4726
rect 7886 4704 8182 4724
rect 13280 4682 13308 18218
rect 13360 18140 13412 18146
rect 13360 18082 13412 18088
rect 13372 17738 13400 18082
rect 13360 17732 13412 17738
rect 13360 17674 13412 17680
rect 13452 15352 13504 15358
rect 13452 15294 13504 15300
rect 13464 15018 13492 15294
rect 13452 15012 13504 15018
rect 13452 14954 13504 14960
rect 13452 12496 13504 12502
rect 13452 12438 13504 12444
rect 13464 12230 13492 12438
rect 13452 12224 13504 12230
rect 13452 12166 13504 12172
rect 13556 9510 13584 20446
rect 13636 20112 13688 20118
rect 13636 20054 13688 20060
rect 13648 19302 13676 20054
rect 13636 19296 13688 19302
rect 13636 19238 13688 19244
rect 13636 18276 13688 18282
rect 13636 18218 13688 18224
rect 13648 18010 13676 18218
rect 13636 18004 13688 18010
rect 13636 17946 13688 17952
rect 13740 17346 13768 22376
rect 13912 19364 13964 19370
rect 13912 19306 13964 19312
rect 13924 18078 13952 19306
rect 14004 18208 14056 18214
rect 14004 18150 14056 18156
rect 13912 18072 13964 18078
rect 13912 18014 13964 18020
rect 14016 17942 14044 18150
rect 14292 18078 14320 22376
rect 14844 20202 14872 22376
rect 14660 20174 14872 20202
rect 14372 19024 14424 19030
rect 14372 18966 14424 18972
rect 14384 18826 14412 18966
rect 14372 18820 14424 18826
rect 14372 18762 14424 18768
rect 14280 18072 14332 18078
rect 14280 18014 14332 18020
rect 14004 17936 14056 17942
rect 14004 17878 14056 17884
rect 13648 17318 13768 17346
rect 13544 9504 13596 9510
rect 13544 9446 13596 9452
rect 13360 9368 13412 9374
rect 13360 9310 13412 9316
rect 13372 8966 13400 9310
rect 13360 8960 13412 8966
rect 13360 8902 13412 8908
rect 13544 8892 13596 8898
rect 13544 8834 13596 8840
rect 13556 8490 13584 8834
rect 13544 8484 13596 8490
rect 13544 8426 13596 8432
rect 13648 8370 13676 17318
rect 13728 16916 13780 16922
rect 13728 16858 13780 16864
rect 13740 16650 13768 16858
rect 13728 16644 13780 16650
rect 13728 16586 13780 16592
rect 13740 15970 13768 16586
rect 13728 15964 13780 15970
rect 13728 15906 13780 15912
rect 14556 15352 14608 15358
rect 14556 15294 14608 15300
rect 13912 15216 13964 15222
rect 13912 15158 13964 15164
rect 13728 14128 13780 14134
rect 13728 14070 13780 14076
rect 13740 12094 13768 14070
rect 13924 13794 13952 15158
rect 14568 14882 14596 15294
rect 14556 14876 14608 14882
rect 14556 14818 14608 14824
rect 14188 14672 14240 14678
rect 14188 14614 14240 14620
rect 14200 14406 14228 14614
rect 14568 14474 14596 14818
rect 14556 14468 14608 14474
rect 14556 14410 14608 14416
rect 14188 14400 14240 14406
rect 14188 14342 14240 14348
rect 14200 13794 14228 14342
rect 13912 13788 13964 13794
rect 13912 13730 13964 13736
rect 14188 13788 14240 13794
rect 14188 13730 14240 13736
rect 13912 13244 13964 13250
rect 13912 13186 13964 13192
rect 13820 12496 13872 12502
rect 13820 12438 13872 12444
rect 13728 12088 13780 12094
rect 13728 12030 13780 12036
rect 13740 10870 13768 12030
rect 13832 11618 13860 12438
rect 13924 11958 13952 13186
rect 13912 11952 13964 11958
rect 13912 11894 13964 11900
rect 13820 11612 13872 11618
rect 13820 11554 13872 11560
rect 14464 11068 14516 11074
rect 14464 11010 14516 11016
rect 14188 10932 14240 10938
rect 14188 10874 14240 10880
rect 13728 10864 13780 10870
rect 13728 10806 13780 10812
rect 14200 10530 14228 10874
rect 14476 10598 14504 11010
rect 14464 10592 14516 10598
rect 14464 10534 14516 10540
rect 14188 10524 14240 10530
rect 14188 10466 14240 10472
rect 14188 10320 14240 10326
rect 14188 10262 14240 10268
rect 14200 10122 14228 10262
rect 14188 10116 14240 10122
rect 14188 10058 14240 10064
rect 14476 9986 14504 10534
rect 14464 9980 14516 9986
rect 14464 9922 14516 9928
rect 14476 9850 14504 9922
rect 14464 9844 14516 9850
rect 14464 9786 14516 9792
rect 14660 9594 14688 20174
rect 14817 20012 15113 20032
rect 14873 20010 14897 20012
rect 14953 20010 14977 20012
rect 15033 20010 15057 20012
rect 14895 19958 14897 20010
rect 14959 19958 14971 20010
rect 15033 19958 15035 20010
rect 14873 19956 14897 19958
rect 14953 19956 14977 19958
rect 15033 19956 15057 19958
rect 14817 19936 15113 19956
rect 15198 19944 15254 19953
rect 15198 19879 15200 19888
rect 15252 19879 15254 19888
rect 15200 19850 15252 19856
rect 15108 19840 15160 19846
rect 15108 19782 15160 19788
rect 15120 19234 15148 19782
rect 15396 19658 15424 22376
rect 15844 19772 15896 19778
rect 15844 19714 15896 19720
rect 15660 19704 15712 19710
rect 15396 19630 15516 19658
rect 15384 19568 15436 19574
rect 15384 19510 15436 19516
rect 15108 19228 15160 19234
rect 15108 19170 15160 19176
rect 15396 19166 15424 19510
rect 15292 19160 15344 19166
rect 15292 19102 15344 19108
rect 15384 19160 15436 19166
rect 15384 19102 15436 19108
rect 15200 19092 15252 19098
rect 15200 19034 15252 19040
rect 15212 19001 15240 19034
rect 15198 18992 15254 19001
rect 14817 18924 15113 18944
rect 15198 18927 15254 18936
rect 14873 18922 14897 18924
rect 14953 18922 14977 18924
rect 15033 18922 15057 18924
rect 14895 18870 14897 18922
rect 14959 18870 14971 18922
rect 15033 18870 15035 18922
rect 14873 18868 14897 18870
rect 14953 18868 14977 18870
rect 15033 18868 15057 18870
rect 14817 18848 15113 18868
rect 15304 18622 15332 19102
rect 15292 18616 15344 18622
rect 14738 18584 14794 18593
rect 15292 18558 15344 18564
rect 14738 18519 14794 18528
rect 14752 18486 14780 18519
rect 14740 18480 14792 18486
rect 14740 18422 14792 18428
rect 14740 18072 14792 18078
rect 14740 18014 14792 18020
rect 13556 8342 13676 8370
rect 14568 9566 14688 9594
rect 14188 8348 14240 8354
rect 13556 5770 13584 8342
rect 14188 8290 14240 8296
rect 13636 8212 13688 8218
rect 13636 8154 13688 8160
rect 13648 6586 13676 8154
rect 13912 8144 13964 8150
rect 13912 8086 13964 8092
rect 13924 7946 13952 8086
rect 13912 7940 13964 7946
rect 13912 7882 13964 7888
rect 14200 7878 14228 8290
rect 14280 8144 14332 8150
rect 14280 8086 14332 8092
rect 14188 7872 14240 7878
rect 14188 7814 14240 7820
rect 14200 7402 14228 7814
rect 14292 7742 14320 8086
rect 14280 7736 14332 7742
rect 14280 7678 14332 7684
rect 14188 7396 14240 7402
rect 14188 7338 14240 7344
rect 13728 6784 13780 6790
rect 13728 6726 13780 6732
rect 13636 6580 13688 6586
rect 13636 6522 13688 6528
rect 13544 5764 13596 5770
rect 13544 5706 13596 5712
rect 13268 4676 13320 4682
rect 13268 4618 13320 4624
rect 4421 4236 4717 4256
rect 4477 4234 4501 4236
rect 4557 4234 4581 4236
rect 4637 4234 4661 4236
rect 4499 4182 4501 4234
rect 4563 4182 4575 4234
rect 4637 4182 4639 4234
rect 4477 4180 4501 4182
rect 4557 4180 4581 4182
rect 4637 4180 4661 4182
rect 4421 4160 4717 4180
rect 11352 4236 11648 4256
rect 11408 4234 11432 4236
rect 11488 4234 11512 4236
rect 11568 4234 11592 4236
rect 11430 4182 11432 4234
rect 11494 4182 11506 4234
rect 11568 4182 11570 4234
rect 11408 4180 11432 4182
rect 11488 4180 11512 4182
rect 11568 4180 11592 4182
rect 11352 4160 11648 4180
rect 13740 3934 13768 6726
rect 14568 6518 14596 9566
rect 14752 9458 14780 18014
rect 14817 17836 15113 17856
rect 14873 17834 14897 17836
rect 14953 17834 14977 17836
rect 15033 17834 15057 17836
rect 14895 17782 14897 17834
rect 14959 17782 14971 17834
rect 15033 17782 15035 17834
rect 14873 17780 14897 17782
rect 14953 17780 14977 17782
rect 15033 17780 15057 17782
rect 14817 17760 15113 17780
rect 15108 17528 15160 17534
rect 15108 17470 15160 17476
rect 15120 17194 15148 17470
rect 15108 17188 15160 17194
rect 15108 17130 15160 17136
rect 15304 16990 15332 18558
rect 15488 18282 15516 19630
rect 15580 19652 15660 19658
rect 15580 19646 15712 19652
rect 15580 19630 15700 19646
rect 15580 19166 15608 19630
rect 15568 19160 15620 19166
rect 15568 19102 15620 19108
rect 15384 18276 15436 18282
rect 15384 18218 15436 18224
rect 15476 18276 15528 18282
rect 15476 18218 15528 18224
rect 15292 16984 15344 16990
rect 15292 16926 15344 16932
rect 15200 16916 15252 16922
rect 15200 16858 15252 16864
rect 14817 16748 15113 16768
rect 14873 16746 14897 16748
rect 14953 16746 14977 16748
rect 15033 16746 15057 16748
rect 14895 16694 14897 16746
rect 14959 16694 14971 16746
rect 15033 16694 15035 16746
rect 14873 16692 14897 16694
rect 14953 16692 14977 16694
rect 15033 16692 15057 16694
rect 14817 16672 15113 16692
rect 15212 16650 15240 16858
rect 15200 16644 15252 16650
rect 15200 16586 15252 16592
rect 15304 16446 15332 16926
rect 15292 16440 15344 16446
rect 15292 16382 15344 16388
rect 14817 15660 15113 15680
rect 14873 15658 14897 15660
rect 14953 15658 14977 15660
rect 15033 15658 15057 15660
rect 14895 15606 14897 15658
rect 14959 15606 14971 15658
rect 15033 15606 15035 15658
rect 14873 15604 14897 15606
rect 14953 15604 14977 15606
rect 15033 15604 15057 15606
rect 14817 15584 15113 15604
rect 15200 15420 15252 15426
rect 15200 15362 15252 15368
rect 14817 14572 15113 14592
rect 14873 14570 14897 14572
rect 14953 14570 14977 14572
rect 15033 14570 15057 14572
rect 14895 14518 14897 14570
rect 14959 14518 14971 14570
rect 15033 14518 15035 14570
rect 14873 14516 14897 14518
rect 14953 14516 14977 14518
rect 15033 14516 15057 14518
rect 14817 14496 15113 14516
rect 14817 13484 15113 13504
rect 14873 13482 14897 13484
rect 14953 13482 14977 13484
rect 15033 13482 15057 13484
rect 14895 13430 14897 13482
rect 14959 13430 14971 13482
rect 15033 13430 15035 13482
rect 14873 13428 14897 13430
rect 14953 13428 14977 13430
rect 15033 13428 15057 13430
rect 14817 13408 15113 13428
rect 14817 12396 15113 12416
rect 14873 12394 14897 12396
rect 14953 12394 14977 12396
rect 15033 12394 15057 12396
rect 14895 12342 14897 12394
rect 14959 12342 14971 12394
rect 15033 12342 15035 12394
rect 14873 12340 14897 12342
rect 14953 12340 14977 12342
rect 15033 12340 15057 12342
rect 14817 12320 15113 12340
rect 14817 11308 15113 11328
rect 14873 11306 14897 11308
rect 14953 11306 14977 11308
rect 15033 11306 15057 11308
rect 14895 11254 14897 11306
rect 14959 11254 14971 11306
rect 15033 11254 15035 11306
rect 14873 11252 14897 11254
rect 14953 11252 14977 11254
rect 15033 11252 15057 11254
rect 14817 11232 15113 11252
rect 15212 10326 15240 15362
rect 15292 14672 15344 14678
rect 15292 14614 15344 14620
rect 15304 13658 15332 14614
rect 15292 13652 15344 13658
rect 15292 13594 15344 13600
rect 15396 13250 15424 18218
rect 15856 17602 15884 19714
rect 15844 17596 15896 17602
rect 15844 17538 15896 17544
rect 15948 17482 15976 22376
rect 16120 20316 16172 20322
rect 16120 20258 16172 20264
rect 16026 19944 16082 19953
rect 16026 19879 16028 19888
rect 16080 19879 16082 19888
rect 16028 19850 16080 19856
rect 16132 19030 16160 20258
rect 16500 20202 16528 22376
rect 16224 20174 16528 20202
rect 16120 19024 16172 19030
rect 16120 18966 16172 18972
rect 16019 18684 16071 18690
rect 16132 18672 16160 18966
rect 16071 18644 16160 18672
rect 16019 18626 16071 18632
rect 16028 17596 16080 17602
rect 16028 17538 16080 17544
rect 15488 17454 15976 17482
rect 15384 13244 15436 13250
rect 15384 13186 15436 13192
rect 15384 11476 15436 11482
rect 15384 11418 15436 11424
rect 15396 10666 15424 11418
rect 15384 10660 15436 10666
rect 15384 10602 15436 10608
rect 15200 10320 15252 10326
rect 15200 10262 15252 10268
rect 14817 10220 15113 10240
rect 14873 10218 14897 10220
rect 14953 10218 14977 10220
rect 15033 10218 15057 10220
rect 14895 10166 14897 10218
rect 14959 10166 14971 10218
rect 15033 10166 15035 10218
rect 14873 10164 14897 10166
rect 14953 10164 14977 10166
rect 15033 10164 15057 10166
rect 14817 10144 15113 10164
rect 14660 9430 14780 9458
rect 14660 9034 14688 9430
rect 14740 9300 14792 9306
rect 14740 9242 14792 9248
rect 14648 9028 14700 9034
rect 14648 8970 14700 8976
rect 14752 8898 14780 9242
rect 14817 9132 15113 9152
rect 14873 9130 14897 9132
rect 14953 9130 14977 9132
rect 15033 9130 15057 9132
rect 14895 9078 14897 9130
rect 14959 9078 14971 9130
rect 15033 9078 15035 9130
rect 14873 9076 14897 9078
rect 14953 9076 14977 9078
rect 15033 9076 15057 9078
rect 14817 9056 15113 9076
rect 14740 8892 14792 8898
rect 14740 8834 14792 8840
rect 14817 8044 15113 8064
rect 14873 8042 14897 8044
rect 14953 8042 14977 8044
rect 15033 8042 15057 8044
rect 14895 7990 14897 8042
rect 14959 7990 14971 8042
rect 15033 7990 15035 8042
rect 14873 7988 14897 7990
rect 14953 7988 14977 7990
rect 15033 7988 15057 7990
rect 14817 7968 15113 7988
rect 15488 7878 15516 17454
rect 15752 17392 15804 17398
rect 16040 17346 16068 17538
rect 15752 17334 15804 17340
rect 15764 15834 15792 17334
rect 15948 17318 16068 17346
rect 15752 15828 15804 15834
rect 15752 15770 15804 15776
rect 15844 15760 15896 15766
rect 15844 15702 15896 15708
rect 15856 15562 15884 15702
rect 15844 15556 15896 15562
rect 15844 15498 15896 15504
rect 15660 14672 15712 14678
rect 15660 14614 15712 14620
rect 15844 14672 15896 14678
rect 15948 14660 15976 17318
rect 16028 16848 16080 16854
rect 16028 16790 16080 16796
rect 16040 16582 16068 16790
rect 16028 16576 16080 16582
rect 16028 16518 16080 16524
rect 16040 15970 16068 16518
rect 16028 15964 16080 15970
rect 16028 15906 16080 15912
rect 15896 14632 15976 14660
rect 15844 14614 15896 14620
rect 15672 14474 15700 14614
rect 15660 14468 15712 14474
rect 15660 14410 15712 14416
rect 15752 13108 15804 13114
rect 15752 13050 15804 13056
rect 15764 12774 15792 13050
rect 15752 12768 15804 12774
rect 15752 12710 15804 12716
rect 15752 12156 15804 12162
rect 15752 12098 15804 12104
rect 15764 11618 15792 12098
rect 15752 11612 15804 11618
rect 15752 11554 15804 11560
rect 15660 11408 15712 11414
rect 15660 11350 15712 11356
rect 15672 9850 15700 11350
rect 15764 11210 15792 11554
rect 15752 11204 15804 11210
rect 15752 11146 15804 11152
rect 15856 10002 15884 14614
rect 15936 13720 15988 13726
rect 15936 13662 15988 13668
rect 15948 13318 15976 13662
rect 15936 13312 15988 13318
rect 15936 13254 15988 13260
rect 15936 10320 15988 10326
rect 15936 10262 15988 10268
rect 15764 9974 15884 10002
rect 15764 9918 15792 9974
rect 15752 9912 15804 9918
rect 15948 9866 15976 10262
rect 15752 9854 15804 9860
rect 15660 9844 15712 9850
rect 15660 9786 15712 9792
rect 15660 8212 15712 8218
rect 15660 8154 15712 8160
rect 15476 7872 15528 7878
rect 15476 7814 15528 7820
rect 15672 7606 15700 8154
rect 15660 7600 15712 7606
rect 15660 7542 15712 7548
rect 15672 7266 15700 7542
rect 15660 7260 15712 7266
rect 15660 7202 15712 7208
rect 14817 6956 15113 6976
rect 14873 6954 14897 6956
rect 14953 6954 14977 6956
rect 15033 6954 15057 6956
rect 14895 6902 14897 6954
rect 14959 6902 14971 6954
rect 15033 6902 15035 6954
rect 14873 6900 14897 6902
rect 14953 6900 14977 6902
rect 15033 6900 15057 6902
rect 14817 6880 15113 6900
rect 14556 6512 14608 6518
rect 14556 6454 14608 6460
rect 14817 5868 15113 5888
rect 14873 5866 14897 5868
rect 14953 5866 14977 5868
rect 15033 5866 15057 5868
rect 14895 5814 14897 5866
rect 14959 5814 14971 5866
rect 15033 5814 15035 5866
rect 14873 5812 14897 5814
rect 14953 5812 14977 5814
rect 15033 5812 15057 5814
rect 14817 5792 15113 5812
rect 14817 4780 15113 4800
rect 14873 4778 14897 4780
rect 14953 4778 14977 4780
rect 15033 4778 15057 4780
rect 14895 4726 14897 4778
rect 14959 4726 14971 4778
rect 15033 4726 15035 4778
rect 14873 4724 14897 4726
rect 14953 4724 14977 4726
rect 15033 4724 15057 4726
rect 14817 4704 15113 4724
rect 13820 4540 13872 4546
rect 13820 4482 13872 4488
rect 13832 4002 13860 4482
rect 13820 3996 13872 4002
rect 13820 3938 13872 3944
rect 13728 3928 13780 3934
rect 13728 3870 13780 3876
rect 7886 3692 8182 3712
rect 7942 3690 7966 3692
rect 8022 3690 8046 3692
rect 8102 3690 8126 3692
rect 7964 3638 7966 3690
rect 8028 3638 8040 3690
rect 8102 3638 8104 3690
rect 7942 3636 7966 3638
rect 8022 3636 8046 3638
rect 8102 3636 8126 3638
rect 7886 3616 8182 3636
rect 14817 3692 15113 3712
rect 14873 3690 14897 3692
rect 14953 3690 14977 3692
rect 15033 3690 15057 3692
rect 14895 3638 14897 3690
rect 14959 3638 14971 3690
rect 15033 3638 15035 3690
rect 14873 3636 14897 3638
rect 14953 3636 14977 3638
rect 15033 3636 15057 3638
rect 14817 3616 15113 3636
rect 4421 3148 4717 3168
rect 4477 3146 4501 3148
rect 4557 3146 4581 3148
rect 4637 3146 4661 3148
rect 4499 3094 4501 3146
rect 4563 3094 4575 3146
rect 4637 3094 4639 3146
rect 4477 3092 4501 3094
rect 4557 3092 4581 3094
rect 4637 3092 4661 3094
rect 4421 3072 4717 3092
rect 11352 3148 11648 3168
rect 11408 3146 11432 3148
rect 11488 3146 11512 3148
rect 11568 3146 11592 3148
rect 11430 3094 11432 3146
rect 11494 3094 11506 3146
rect 11568 3094 11570 3146
rect 11408 3092 11432 3094
rect 11488 3092 11512 3094
rect 11568 3092 11592 3094
rect 11352 3072 11648 3092
rect 7886 2604 8182 2624
rect 7942 2602 7966 2604
rect 8022 2602 8046 2604
rect 8102 2602 8126 2604
rect 7964 2550 7966 2602
rect 8028 2550 8040 2602
rect 8102 2550 8104 2602
rect 7942 2548 7966 2550
rect 8022 2548 8046 2550
rect 8102 2548 8126 2550
rect 7886 2528 8182 2548
rect 14817 2604 15113 2624
rect 14873 2602 14897 2604
rect 14953 2602 14977 2604
rect 15033 2602 15057 2604
rect 14895 2550 14897 2602
rect 14959 2550 14971 2602
rect 15033 2550 15035 2602
rect 14873 2548 14897 2550
rect 14953 2548 14977 2550
rect 15033 2548 15057 2550
rect 14817 2528 15113 2548
rect 15764 2506 15792 9854
rect 15856 9838 15976 9866
rect 15752 2500 15804 2506
rect 15752 2442 15804 2448
rect 4421 2060 4717 2080
rect 4477 2058 4501 2060
rect 4557 2058 4581 2060
rect 4637 2058 4661 2060
rect 4499 2006 4501 2058
rect 4563 2006 4575 2058
rect 4637 2006 4639 2058
rect 4477 2004 4501 2006
rect 4557 2004 4581 2006
rect 4637 2004 4661 2006
rect 4421 1984 4717 2004
rect 11352 2060 11648 2080
rect 11408 2058 11432 2060
rect 11488 2058 11512 2060
rect 11568 2058 11592 2060
rect 11430 2006 11432 2058
rect 11494 2006 11506 2058
rect 11568 2006 11570 2058
rect 11408 2004 11432 2006
rect 11488 2004 11512 2006
rect 11568 2004 11592 2006
rect 11352 1984 11648 2004
rect 15856 1214 15884 9838
rect 15936 9368 15988 9374
rect 15936 9310 15988 9316
rect 15948 9034 15976 9310
rect 15936 9028 15988 9034
rect 15936 8970 15988 8976
rect 16224 7674 16252 20174
rect 16304 20112 16356 20118
rect 16304 20054 16356 20060
rect 16488 20112 16540 20118
rect 16488 20054 16540 20060
rect 16316 19778 16344 20054
rect 16396 19908 16448 19914
rect 16396 19850 16448 19856
rect 16408 19817 16436 19850
rect 16394 19808 16450 19817
rect 16304 19772 16356 19778
rect 16394 19743 16450 19752
rect 16304 19714 16356 19720
rect 16396 19704 16448 19710
rect 16396 19646 16448 19652
rect 16408 19370 16436 19646
rect 16500 19642 16528 20054
rect 16488 19636 16540 19642
rect 16488 19578 16540 19584
rect 16396 19364 16448 19370
rect 16396 19306 16448 19312
rect 16764 19092 16816 19098
rect 16764 19034 16816 19040
rect 16776 19001 16804 19034
rect 17052 19030 17080 22376
rect 17590 19808 17646 19817
rect 17590 19743 17646 19752
rect 17500 19228 17552 19234
rect 17500 19170 17552 19176
rect 17040 19024 17092 19030
rect 16762 18992 16818 19001
rect 17040 18966 17092 18972
rect 16762 18927 16818 18936
rect 17512 18729 17540 19170
rect 17604 18826 17632 19743
rect 17696 19250 17724 22376
rect 18142 21984 18198 21993
rect 18142 21919 18198 21928
rect 17866 21032 17922 21041
rect 17866 20967 17922 20976
rect 17880 20458 17908 20967
rect 17868 20452 17920 20458
rect 17868 20394 17920 20400
rect 18050 19672 18106 19681
rect 18050 19607 18106 19616
rect 17960 19296 18012 19302
rect 17696 19222 17908 19250
rect 17960 19238 18012 19244
rect 17682 19128 17738 19137
rect 17682 19063 17738 19072
rect 17592 18820 17644 18826
rect 17592 18762 17644 18768
rect 17498 18720 17554 18729
rect 17498 18655 17554 18664
rect 17500 18616 17552 18622
rect 17500 18558 17552 18564
rect 16488 18208 16540 18214
rect 16488 18150 16540 18156
rect 16304 8892 16356 8898
rect 16304 8834 16356 8840
rect 16316 7946 16344 8834
rect 16396 8824 16448 8830
rect 16396 8766 16448 8772
rect 16304 7940 16356 7946
rect 16304 7882 16356 7888
rect 16212 7668 16264 7674
rect 16212 7610 16264 7616
rect 16408 7402 16436 8766
rect 16396 7396 16448 7402
rect 16396 7338 16448 7344
rect 16500 6586 16528 18150
rect 17040 18072 17092 18078
rect 17040 18014 17092 18020
rect 17224 18072 17276 18078
rect 17224 18014 17276 18020
rect 17052 17670 17080 18014
rect 17040 17664 17092 17670
rect 17040 17606 17092 17612
rect 16856 17596 16908 17602
rect 16856 17538 16908 17544
rect 16868 17058 16896 17538
rect 16856 17052 16908 17058
rect 16856 16994 16908 17000
rect 16580 16644 16632 16650
rect 16580 16586 16632 16592
rect 16592 16038 16620 16586
rect 17236 16394 17264 18014
rect 17512 18010 17540 18558
rect 17696 18486 17724 19063
rect 17880 18690 17908 19222
rect 17868 18684 17920 18690
rect 17868 18626 17920 18632
rect 17684 18480 17736 18486
rect 17684 18422 17736 18428
rect 17776 18480 17828 18486
rect 17776 18422 17828 18428
rect 17316 18004 17368 18010
rect 17316 17946 17368 17952
rect 17500 18004 17552 18010
rect 17500 17946 17552 17952
rect 17684 18004 17736 18010
rect 17684 17946 17736 17952
rect 17328 17890 17356 17946
rect 17696 17890 17724 17946
rect 17328 17862 17724 17890
rect 17236 16366 17356 16394
rect 17328 16310 17356 16366
rect 17592 16372 17644 16378
rect 17592 16314 17644 16320
rect 17316 16304 17368 16310
rect 17316 16246 17368 16252
rect 16580 16032 16632 16038
rect 16580 15974 16632 15980
rect 17328 15902 17356 16246
rect 17604 15902 17632 16314
rect 17316 15896 17368 15902
rect 17316 15838 17368 15844
rect 17592 15896 17644 15902
rect 17592 15838 17644 15844
rect 17328 14134 17356 15838
rect 17684 15828 17736 15834
rect 17684 15770 17736 15776
rect 17696 15426 17724 15770
rect 17684 15420 17736 15426
rect 17684 15362 17736 15368
rect 17408 14808 17460 14814
rect 17408 14750 17460 14756
rect 17316 14128 17368 14134
rect 17316 14070 17368 14076
rect 17224 13720 17276 13726
rect 17224 13662 17276 13668
rect 16672 13584 16724 13590
rect 16672 13526 16724 13532
rect 16684 13250 16712 13526
rect 17236 13386 17264 13662
rect 17224 13380 17276 13386
rect 17224 13322 17276 13328
rect 17420 13318 17448 14750
rect 17408 13312 17460 13318
rect 17408 13254 17460 13260
rect 16672 13244 16724 13250
rect 16672 13186 16724 13192
rect 16948 13176 17000 13182
rect 16948 13118 17000 13124
rect 16672 12632 16724 12638
rect 16672 12574 16724 12580
rect 16580 12564 16632 12570
rect 16580 12506 16632 12512
rect 16592 12026 16620 12506
rect 16580 12020 16632 12026
rect 16580 11962 16632 11968
rect 16684 10462 16712 12574
rect 16960 12570 16988 13118
rect 16948 12564 17000 12570
rect 16948 12506 17000 12512
rect 16960 12298 16988 12506
rect 16948 12292 17000 12298
rect 16948 12234 17000 12240
rect 17788 11210 17816 18422
rect 17972 18185 18000 19238
rect 18064 19234 18092 19607
rect 18156 19250 18184 21919
rect 18248 20746 18276 22376
rect 18248 20718 18644 20746
rect 18282 20556 18578 20576
rect 18338 20554 18362 20556
rect 18418 20554 18442 20556
rect 18498 20554 18522 20556
rect 18360 20502 18362 20554
rect 18424 20502 18436 20554
rect 18498 20502 18500 20554
rect 18338 20500 18362 20502
rect 18418 20500 18442 20502
rect 18498 20500 18522 20502
rect 18282 20480 18578 20500
rect 18282 19468 18578 19488
rect 18338 19466 18362 19468
rect 18418 19466 18442 19468
rect 18498 19466 18522 19468
rect 18360 19414 18362 19466
rect 18424 19414 18436 19466
rect 18498 19414 18500 19466
rect 18338 19412 18362 19414
rect 18418 19412 18442 19414
rect 18498 19412 18522 19414
rect 18282 19392 18578 19412
rect 18052 19228 18104 19234
rect 18156 19222 18276 19250
rect 18052 19170 18104 19176
rect 18144 19160 18196 19166
rect 18144 19102 18196 19108
rect 18052 18820 18104 18826
rect 18052 18762 18104 18768
rect 17958 18176 18014 18185
rect 17958 18111 18014 18120
rect 18064 17738 18092 18762
rect 18052 17732 18104 17738
rect 18052 17674 18104 17680
rect 17868 17596 17920 17602
rect 17868 17538 17920 17544
rect 17880 17466 17908 17538
rect 18156 17466 18184 19102
rect 18248 18593 18276 19222
rect 18510 18992 18566 19001
rect 18510 18927 18566 18936
rect 18524 18826 18552 18927
rect 18616 18826 18644 20718
rect 18696 20180 18748 20186
rect 18696 20122 18748 20128
rect 18512 18820 18564 18826
rect 18512 18762 18564 18768
rect 18604 18820 18656 18826
rect 18604 18762 18656 18768
rect 18418 18720 18474 18729
rect 18418 18655 18420 18664
rect 18472 18655 18474 18664
rect 18420 18626 18472 18632
rect 18234 18584 18290 18593
rect 18234 18519 18290 18528
rect 18602 18584 18658 18593
rect 18602 18519 18658 18528
rect 18282 18380 18578 18400
rect 18338 18378 18362 18380
rect 18418 18378 18442 18380
rect 18498 18378 18522 18380
rect 18360 18326 18362 18378
rect 18424 18326 18436 18378
rect 18498 18326 18500 18378
rect 18338 18324 18362 18326
rect 18418 18324 18442 18326
rect 18498 18324 18522 18326
rect 18282 18304 18578 18324
rect 18616 18282 18644 18519
rect 18604 18276 18656 18282
rect 18604 18218 18656 18224
rect 18236 18208 18288 18214
rect 18236 18150 18288 18156
rect 18248 17942 18276 18150
rect 18708 18010 18736 20122
rect 18696 18004 18748 18010
rect 18696 17946 18748 17952
rect 18236 17936 18288 17942
rect 18236 17878 18288 17884
rect 18604 17936 18656 17942
rect 18604 17878 18656 17884
rect 18616 17534 18644 17878
rect 18604 17528 18656 17534
rect 18604 17470 18656 17476
rect 17868 17460 17920 17466
rect 17868 17402 17920 17408
rect 18144 17460 18196 17466
rect 18144 17402 18196 17408
rect 17960 17392 18012 17398
rect 17960 17334 18012 17340
rect 17972 16689 18000 17334
rect 18282 17292 18578 17312
rect 18338 17290 18362 17292
rect 18418 17290 18442 17292
rect 18498 17290 18522 17292
rect 18360 17238 18362 17290
rect 18424 17238 18436 17290
rect 18498 17238 18500 17290
rect 18338 17236 18362 17238
rect 18418 17236 18442 17238
rect 18498 17236 18522 17238
rect 18282 17216 18578 17236
rect 18800 17194 18828 22376
rect 18970 20624 19026 20633
rect 18970 20559 19026 20568
rect 18878 20080 18934 20089
rect 18878 20015 18934 20024
rect 18892 18214 18920 20015
rect 18880 18208 18932 18214
rect 18880 18150 18932 18156
rect 18984 18146 19012 20559
rect 19076 18146 19104 22463
rect 19338 22376 19394 22856
rect 19890 22376 19946 22856
rect 20442 22376 20498 22856
rect 20994 22376 21050 22856
rect 21546 22376 21602 22856
rect 22098 22376 22154 22856
rect 22650 22376 22706 22856
rect 19154 21576 19210 21585
rect 19154 21511 19210 21520
rect 18972 18140 19024 18146
rect 18972 18082 19024 18088
rect 19064 18140 19116 18146
rect 19064 18082 19116 18088
rect 18880 18072 18932 18078
rect 19168 18026 19196 21511
rect 19248 20112 19300 20118
rect 19248 20054 19300 20060
rect 18880 18014 18932 18020
rect 18144 17188 18196 17194
rect 18144 17130 18196 17136
rect 18788 17188 18840 17194
rect 18788 17130 18840 17136
rect 18050 17088 18106 17097
rect 18050 17023 18106 17032
rect 17958 16680 18014 16689
rect 17958 16615 18014 16624
rect 18064 16394 18092 17023
rect 17972 16366 18092 16394
rect 17972 15562 18000 16366
rect 18052 16304 18104 16310
rect 18052 16246 18104 16252
rect 18064 15562 18092 16246
rect 17960 15556 18012 15562
rect 17960 15498 18012 15504
rect 18052 15556 18104 15562
rect 18052 15498 18104 15504
rect 17958 14232 18014 14241
rect 17958 14167 18014 14176
rect 17972 13930 18000 14167
rect 17960 13924 18012 13930
rect 17960 13866 18012 13872
rect 18156 13674 18184 17130
rect 18602 16952 18658 16961
rect 18602 16887 18658 16896
rect 18512 16440 18564 16446
rect 18616 16428 18644 16887
rect 18564 16400 18644 16428
rect 18512 16382 18564 16388
rect 18282 16204 18578 16224
rect 18338 16202 18362 16204
rect 18418 16202 18442 16204
rect 18498 16202 18522 16204
rect 18360 16150 18362 16202
rect 18424 16150 18436 16202
rect 18498 16150 18500 16202
rect 18338 16148 18362 16150
rect 18418 16148 18442 16150
rect 18498 16148 18522 16150
rect 18282 16128 18578 16148
rect 18282 15116 18578 15136
rect 18338 15114 18362 15116
rect 18418 15114 18442 15116
rect 18498 15114 18522 15116
rect 18360 15062 18362 15114
rect 18424 15062 18436 15114
rect 18498 15062 18500 15114
rect 18338 15060 18362 15062
rect 18418 15060 18442 15062
rect 18498 15060 18522 15062
rect 18282 15040 18578 15060
rect 18616 14898 18644 16400
rect 18788 15760 18840 15766
rect 18788 15702 18840 15708
rect 18800 15358 18828 15702
rect 18892 15442 18920 18014
rect 18984 17998 19196 18026
rect 18984 16922 19012 17998
rect 19156 17936 19208 17942
rect 19156 17878 19208 17884
rect 19064 16984 19116 16990
rect 19064 16926 19116 16932
rect 18972 16916 19024 16922
rect 18972 16858 19024 16864
rect 18892 15414 19012 15442
rect 18788 15352 18840 15358
rect 18788 15294 18840 15300
rect 18880 15352 18932 15358
rect 18880 15294 18932 15300
rect 18694 15184 18750 15193
rect 18694 15119 18750 15128
rect 18708 15018 18736 15119
rect 18696 15012 18748 15018
rect 18696 14954 18748 14960
rect 18616 14870 18736 14898
rect 18892 14882 18920 15294
rect 18604 14672 18656 14678
rect 18602 14640 18604 14649
rect 18656 14640 18658 14649
rect 18602 14575 18658 14584
rect 18282 14028 18578 14048
rect 18338 14026 18362 14028
rect 18418 14026 18442 14028
rect 18498 14026 18522 14028
rect 18360 13974 18362 14026
rect 18424 13974 18436 14026
rect 18498 13974 18500 14026
rect 18338 13972 18362 13974
rect 18418 13972 18442 13974
rect 18498 13972 18522 13974
rect 18282 13952 18578 13972
rect 18064 13646 18184 13674
rect 17960 13244 18012 13250
rect 17960 13186 18012 13192
rect 17972 11618 18000 13186
rect 18064 12298 18092 13646
rect 18144 13584 18196 13590
rect 18144 13526 18196 13532
rect 18604 13584 18656 13590
rect 18604 13526 18656 13532
rect 18156 12706 18184 13526
rect 18282 12940 18578 12960
rect 18338 12938 18362 12940
rect 18418 12938 18442 12940
rect 18498 12938 18522 12940
rect 18360 12886 18362 12938
rect 18424 12886 18436 12938
rect 18498 12886 18500 12938
rect 18338 12884 18362 12886
rect 18418 12884 18442 12886
rect 18498 12884 18522 12886
rect 18282 12864 18578 12884
rect 18144 12700 18196 12706
rect 18144 12642 18196 12648
rect 18616 12502 18644 13526
rect 18708 13386 18736 14870
rect 18880 14876 18932 14882
rect 18880 14818 18932 14824
rect 18984 13862 19012 15414
rect 19076 14882 19104 16926
rect 19168 16145 19196 17878
rect 19260 17641 19288 20054
rect 19246 17632 19302 17641
rect 19246 17567 19302 17576
rect 19248 16848 19300 16854
rect 19248 16790 19300 16796
rect 19154 16136 19210 16145
rect 19154 16071 19210 16080
rect 19260 15737 19288 16790
rect 19246 15728 19302 15737
rect 19246 15663 19302 15672
rect 19248 15420 19300 15426
rect 19248 15362 19300 15368
rect 19064 14876 19116 14882
rect 19064 14818 19116 14824
rect 19064 14468 19116 14474
rect 19064 14410 19116 14416
rect 18972 13856 19024 13862
rect 18972 13798 19024 13804
rect 18696 13380 18748 13386
rect 18696 13322 18748 13328
rect 18972 13380 19024 13386
rect 18972 13322 19024 13328
rect 18880 13176 18932 13182
rect 18880 13118 18932 13124
rect 18604 12496 18656 12502
rect 18604 12438 18656 12444
rect 18052 12292 18104 12298
rect 18052 12234 18104 12240
rect 18420 12224 18472 12230
rect 18418 12192 18420 12201
rect 18472 12192 18474 12201
rect 18144 12156 18196 12162
rect 18418 12127 18474 12136
rect 18144 12098 18196 12104
rect 18156 11618 18184 12098
rect 18282 11852 18578 11872
rect 18338 11850 18362 11852
rect 18418 11850 18442 11852
rect 18498 11850 18522 11852
rect 18360 11798 18362 11850
rect 18424 11798 18436 11850
rect 18498 11798 18500 11850
rect 18338 11796 18362 11798
rect 18418 11796 18442 11798
rect 18498 11796 18522 11798
rect 18282 11776 18578 11796
rect 17960 11612 18012 11618
rect 17960 11554 18012 11560
rect 18144 11612 18196 11618
rect 18144 11554 18196 11560
rect 18052 11544 18104 11550
rect 18052 11486 18104 11492
rect 17958 11240 18014 11249
rect 17776 11204 17828 11210
rect 18064 11210 18092 11486
rect 17958 11175 18014 11184
rect 18052 11204 18104 11210
rect 17776 11146 17828 11152
rect 17972 11074 18000 11175
rect 18052 11146 18104 11152
rect 17960 11068 18012 11074
rect 17960 11010 18012 11016
rect 18144 11068 18196 11074
rect 18144 11010 18196 11016
rect 18052 11000 18104 11006
rect 18052 10942 18104 10948
rect 16672 10456 16724 10462
rect 16672 10398 16724 10404
rect 16684 9374 16712 10398
rect 17960 10388 18012 10394
rect 17960 10330 18012 10336
rect 17972 9850 18000 10330
rect 18064 10122 18092 10942
rect 18052 10116 18104 10122
rect 18052 10058 18104 10064
rect 18052 9912 18104 9918
rect 18052 9854 18104 9860
rect 17960 9844 18012 9850
rect 17960 9786 18012 9792
rect 17972 9578 18000 9786
rect 17960 9572 18012 9578
rect 17960 9514 18012 9520
rect 16672 9368 16724 9374
rect 16672 9310 16724 9316
rect 16580 9232 16632 9238
rect 16580 9174 16632 9180
rect 16592 8830 16620 9174
rect 16580 8824 16632 8830
rect 16580 8766 16632 8772
rect 16592 8490 16620 8766
rect 16580 8484 16632 8490
rect 16580 8426 16632 8432
rect 16684 8286 16712 9310
rect 16672 8280 16724 8286
rect 16672 8222 16724 8228
rect 18064 7198 18092 9854
rect 18156 9034 18184 11010
rect 18282 10764 18578 10784
rect 18338 10762 18362 10764
rect 18418 10762 18442 10764
rect 18498 10762 18522 10764
rect 18360 10710 18362 10762
rect 18424 10710 18436 10762
rect 18498 10710 18500 10762
rect 18338 10708 18362 10710
rect 18418 10708 18442 10710
rect 18498 10708 18522 10710
rect 18282 10688 18578 10708
rect 18282 9676 18578 9696
rect 18338 9674 18362 9676
rect 18418 9674 18442 9676
rect 18498 9674 18522 9676
rect 18360 9622 18362 9674
rect 18424 9622 18436 9674
rect 18498 9622 18500 9674
rect 18338 9620 18362 9622
rect 18418 9620 18442 9622
rect 18498 9620 18522 9622
rect 18282 9600 18578 9620
rect 18144 9028 18196 9034
rect 18144 8970 18196 8976
rect 18282 8588 18578 8608
rect 18338 8586 18362 8588
rect 18418 8586 18442 8588
rect 18498 8586 18522 8588
rect 18360 8534 18362 8586
rect 18424 8534 18436 8586
rect 18498 8534 18500 8586
rect 18338 8532 18362 8534
rect 18418 8532 18442 8534
rect 18498 8532 18522 8534
rect 18282 8512 18578 8532
rect 18282 7500 18578 7520
rect 18338 7498 18362 7500
rect 18418 7498 18442 7500
rect 18498 7498 18522 7500
rect 18360 7446 18362 7498
rect 18424 7446 18436 7498
rect 18498 7446 18500 7498
rect 18338 7444 18362 7446
rect 18418 7444 18442 7446
rect 18498 7444 18522 7446
rect 18282 7424 18578 7444
rect 16948 7192 17000 7198
rect 16948 7134 17000 7140
rect 18052 7192 18104 7198
rect 18052 7134 18104 7140
rect 16960 6722 16988 7134
rect 17960 6784 18012 6790
rect 17960 6726 18012 6732
rect 16948 6716 17000 6722
rect 16948 6658 17000 6664
rect 16488 6580 16540 6586
rect 16488 6522 16540 6528
rect 17972 4449 18000 6726
rect 18282 6412 18578 6432
rect 18338 6410 18362 6412
rect 18418 6410 18442 6412
rect 18498 6410 18522 6412
rect 18360 6358 18362 6410
rect 18424 6358 18436 6410
rect 18498 6358 18500 6410
rect 18338 6356 18362 6358
rect 18418 6356 18442 6358
rect 18498 6356 18522 6358
rect 18282 6336 18578 6356
rect 18282 5324 18578 5344
rect 18338 5322 18362 5324
rect 18418 5322 18442 5324
rect 18498 5322 18522 5324
rect 18360 5270 18362 5322
rect 18424 5270 18436 5322
rect 18498 5270 18500 5322
rect 18338 5268 18362 5270
rect 18418 5268 18442 5270
rect 18498 5268 18522 5270
rect 18282 5248 18578 5268
rect 17958 4440 18014 4449
rect 17958 4375 18014 4384
rect 18282 4236 18578 4256
rect 18338 4234 18362 4236
rect 18418 4234 18442 4236
rect 18498 4234 18522 4236
rect 18360 4182 18362 4234
rect 18424 4182 18436 4234
rect 18498 4182 18500 4234
rect 18338 4180 18362 4182
rect 18418 4180 18442 4182
rect 18498 4180 18522 4182
rect 18282 4160 18578 4180
rect 17960 3996 18012 4002
rect 17960 3938 18012 3944
rect 17972 3905 18000 3938
rect 18052 3928 18104 3934
rect 17958 3896 18014 3905
rect 18052 3870 18104 3876
rect 17958 3831 18014 3840
rect 18064 3497 18092 3870
rect 18050 3488 18106 3497
rect 18050 3423 18106 3432
rect 18282 3148 18578 3168
rect 18338 3146 18362 3148
rect 18418 3146 18442 3148
rect 18498 3146 18522 3148
rect 18360 3094 18362 3146
rect 18424 3094 18436 3146
rect 18498 3094 18500 3146
rect 18338 3092 18362 3094
rect 18418 3092 18442 3094
rect 18498 3092 18522 3094
rect 18282 3072 18578 3092
rect 18282 2060 18578 2080
rect 18338 2058 18362 2060
rect 18418 2058 18442 2060
rect 18498 2058 18522 2060
rect 18360 2006 18362 2058
rect 18424 2006 18436 2058
rect 18498 2006 18500 2058
rect 18338 2004 18362 2006
rect 18418 2004 18442 2006
rect 18498 2004 18522 2006
rect 18282 1984 18578 2004
rect 18616 1457 18644 12438
rect 18892 12314 18920 13118
rect 18984 12638 19012 13322
rect 18972 12632 19024 12638
rect 18972 12574 19024 12580
rect 18984 12450 19012 12574
rect 19076 12570 19104 14410
rect 19156 14332 19208 14338
rect 19156 14274 19208 14280
rect 19168 13794 19196 14274
rect 19156 13788 19208 13794
rect 19156 13730 19208 13736
rect 19168 13182 19196 13730
rect 19260 13658 19288 15362
rect 19352 15222 19380 22376
rect 19432 19908 19484 19914
rect 19432 19850 19484 19856
rect 19444 18690 19472 19850
rect 19432 18684 19484 18690
rect 19432 18626 19484 18632
rect 19800 18616 19852 18622
rect 19800 18558 19852 18564
rect 19708 18072 19760 18078
rect 19708 18014 19760 18020
rect 19616 18004 19668 18010
rect 19616 17946 19668 17952
rect 19524 16984 19576 16990
rect 19524 16926 19576 16932
rect 19536 16106 19564 16926
rect 19524 16100 19576 16106
rect 19524 16042 19576 16048
rect 19524 15896 19576 15902
rect 19524 15838 19576 15844
rect 19432 15488 19484 15494
rect 19432 15430 19484 15436
rect 19340 15216 19392 15222
rect 19340 15158 19392 15164
rect 19444 15018 19472 15430
rect 19536 15290 19564 15838
rect 19524 15284 19576 15290
rect 19524 15226 19576 15232
rect 19628 15170 19656 17946
rect 19720 16582 19748 18014
rect 19708 16576 19760 16582
rect 19708 16518 19760 16524
rect 19536 15142 19656 15170
rect 19432 15012 19484 15018
rect 19432 14954 19484 14960
rect 19430 14912 19486 14921
rect 19430 14847 19432 14856
rect 19484 14847 19486 14856
rect 19432 14818 19484 14824
rect 19338 14776 19394 14785
rect 19338 14711 19340 14720
rect 19392 14711 19394 14720
rect 19340 14682 19392 14688
rect 19248 13652 19300 13658
rect 19248 13594 19300 13600
rect 19156 13176 19208 13182
rect 19156 13118 19208 13124
rect 19168 12774 19196 13118
rect 19248 13040 19300 13046
rect 19248 12982 19300 12988
rect 19156 12768 19208 12774
rect 19156 12710 19208 12716
rect 19260 12638 19288 12982
rect 19248 12632 19300 12638
rect 19248 12574 19300 12580
rect 19064 12564 19116 12570
rect 19064 12506 19116 12512
rect 18984 12422 19196 12450
rect 18892 12286 19104 12314
rect 18696 12020 18748 12026
rect 18696 11962 18748 11968
rect 18708 11793 18736 11962
rect 18694 11784 18750 11793
rect 18694 11719 18750 11728
rect 18972 11136 19024 11142
rect 18972 11078 19024 11084
rect 18696 11000 18748 11006
rect 18696 10942 18748 10948
rect 18708 10326 18736 10942
rect 18696 10320 18748 10326
rect 18696 10262 18748 10268
rect 18880 9980 18932 9986
rect 18880 9922 18932 9928
rect 18892 9345 18920 9922
rect 18878 9336 18934 9345
rect 18878 9271 18934 9280
rect 18880 9232 18932 9238
rect 18880 9174 18932 9180
rect 18696 7124 18748 7130
rect 18696 7066 18748 7072
rect 18708 5401 18736 7066
rect 18694 5392 18750 5401
rect 18694 5327 18750 5336
rect 18602 1448 18658 1457
rect 18602 1383 18658 1392
rect 15844 1208 15896 1214
rect 15844 1150 15896 1156
rect 18892 505 18920 9174
rect 18878 496 18934 505
rect 18878 431 18934 440
rect 18984 97 19012 11078
rect 19076 9442 19104 12286
rect 19064 9436 19116 9442
rect 19064 9378 19116 9384
rect 19168 2409 19196 12422
rect 19248 10456 19300 10462
rect 19248 10398 19300 10404
rect 19260 9753 19288 10398
rect 19246 9744 19302 9753
rect 19246 9679 19302 9688
rect 19536 9510 19564 15142
rect 19706 14912 19762 14921
rect 19706 14847 19708 14856
rect 19760 14847 19762 14856
rect 19708 14818 19760 14824
rect 19614 12736 19670 12745
rect 19614 12671 19670 12680
rect 19628 12298 19656 12671
rect 19616 12292 19668 12298
rect 19616 12234 19668 12240
rect 19708 12156 19760 12162
rect 19708 12098 19760 12104
rect 19720 11618 19748 12098
rect 19708 11612 19760 11618
rect 19708 11554 19760 11560
rect 19706 10832 19762 10841
rect 19706 10767 19762 10776
rect 19524 9504 19576 9510
rect 19524 9446 19576 9452
rect 19720 9374 19748 10767
rect 19708 9368 19760 9374
rect 19708 9310 19760 9316
rect 19812 9034 19840 18558
rect 19904 18146 19932 22376
rect 19984 19704 20036 19710
rect 19984 19646 20036 19652
rect 19996 19098 20024 19646
rect 19984 19092 20036 19098
rect 19984 19034 20036 19040
rect 19892 18140 19944 18146
rect 19892 18082 19944 18088
rect 20352 18140 20404 18146
rect 20352 18082 20404 18088
rect 19890 18040 19946 18049
rect 19890 17975 19946 17984
rect 19904 17602 19932 17975
rect 19892 17596 19944 17602
rect 19892 17538 19944 17544
rect 19984 15420 20036 15426
rect 19984 15362 20036 15368
rect 19892 15216 19944 15222
rect 19892 15158 19944 15164
rect 19904 10666 19932 15158
rect 19996 14785 20024 15362
rect 19982 14776 20038 14785
rect 19982 14711 20038 14720
rect 20168 13244 20220 13250
rect 20168 13186 20220 13192
rect 20180 12842 20208 13186
rect 20168 12836 20220 12842
rect 20168 12778 20220 12784
rect 20364 11210 20392 18082
rect 20456 18010 20484 22376
rect 21008 18486 21036 22376
rect 21088 19024 21140 19030
rect 21088 18966 21140 18972
rect 20996 18480 21048 18486
rect 20996 18422 21048 18428
rect 20444 18004 20496 18010
rect 20444 17946 20496 17952
rect 20996 17392 21048 17398
rect 20996 17334 21048 17340
rect 20444 14332 20496 14338
rect 20444 14274 20496 14280
rect 20456 13318 20484 14274
rect 20628 14128 20680 14134
rect 20628 14070 20680 14076
rect 20536 13720 20588 13726
rect 20536 13662 20588 13668
rect 20444 13312 20496 13318
rect 20444 13254 20496 13260
rect 20548 12162 20576 13662
rect 20640 13289 20668 14070
rect 20718 13688 20774 13697
rect 20718 13623 20774 13632
rect 20626 13280 20682 13289
rect 20626 13215 20682 13224
rect 20732 12298 20760 13623
rect 20720 12292 20772 12298
rect 20720 12234 20772 12240
rect 20536 12156 20588 12162
rect 20536 12098 20588 12104
rect 21008 11958 21036 17334
rect 20996 11952 21048 11958
rect 20996 11894 21048 11900
rect 20352 11204 20404 11210
rect 20352 11146 20404 11152
rect 20352 11068 20404 11074
rect 20352 11010 20404 11016
rect 19892 10660 19944 10666
rect 19892 10602 19944 10608
rect 20364 10297 20392 11010
rect 20350 10288 20406 10297
rect 20350 10223 20406 10232
rect 20536 9980 20588 9986
rect 20536 9922 20588 9928
rect 19800 9028 19852 9034
rect 19800 8970 19852 8976
rect 19248 8892 19300 8898
rect 19248 8834 19300 8840
rect 19260 8393 19288 8834
rect 20548 8801 20576 9922
rect 21100 9034 21128 18966
rect 21364 18820 21416 18826
rect 21364 18762 21416 18768
rect 21180 17936 21232 17942
rect 21180 17878 21232 17884
rect 21088 9028 21140 9034
rect 21088 8970 21140 8976
rect 20628 8892 20680 8898
rect 20628 8834 20680 8840
rect 20534 8792 20590 8801
rect 20534 8727 20590 8736
rect 19246 8384 19302 8393
rect 19246 8319 19302 8328
rect 20640 7849 20668 8834
rect 20626 7840 20682 7849
rect 19248 7804 19300 7810
rect 19248 7746 19300 7752
rect 20536 7804 20588 7810
rect 20626 7775 20682 7784
rect 20536 7746 20588 7752
rect 19260 7305 19288 7746
rect 19246 7296 19302 7305
rect 19246 7231 19302 7240
rect 20548 6897 20576 7746
rect 20534 6888 20590 6897
rect 20534 6823 20590 6832
rect 19248 6716 19300 6722
rect 19248 6658 19300 6664
rect 20536 6716 20588 6722
rect 20536 6658 20588 6664
rect 19260 6353 19288 6658
rect 19246 6344 19302 6353
rect 19246 6279 19302 6288
rect 20548 5945 20576 6658
rect 20534 5936 20590 5945
rect 20534 5871 20590 5880
rect 20536 5628 20588 5634
rect 20536 5570 20588 5576
rect 20548 4857 20576 5570
rect 20534 4848 20590 4857
rect 20534 4783 20590 4792
rect 21192 3594 21220 17878
rect 21376 10122 21404 18762
rect 21560 13114 21588 22376
rect 22112 17398 22140 22376
rect 22664 17942 22692 22376
rect 22652 17936 22704 17942
rect 22652 17878 22704 17884
rect 22100 17392 22152 17398
rect 22100 17334 22152 17340
rect 21548 13108 21600 13114
rect 21548 13050 21600 13056
rect 21364 10116 21416 10122
rect 21364 10058 21416 10064
rect 21180 3588 21232 3594
rect 21180 3530 21232 3536
rect 20536 3452 20588 3458
rect 20536 3394 20588 3400
rect 20548 2953 20576 3394
rect 20534 2944 20590 2953
rect 20534 2879 20590 2888
rect 19248 2500 19300 2506
rect 19248 2442 19300 2448
rect 19154 2400 19210 2409
rect 19154 2335 19210 2344
rect 19260 2001 19288 2442
rect 19246 1992 19302 2001
rect 19246 1927 19302 1936
rect 19248 1208 19300 1214
rect 19248 1150 19300 1156
rect 19260 1049 19288 1150
rect 19246 1040 19302 1049
rect 19246 975 19302 984
rect 18970 88 19026 97
rect 18970 23 19026 32
<< via2 >>
rect 19062 22472 19118 22528
rect 4421 20554 4477 20556
rect 4501 20554 4557 20556
rect 4581 20554 4637 20556
rect 4661 20554 4717 20556
rect 4421 20502 4447 20554
rect 4447 20502 4477 20554
rect 4501 20502 4511 20554
rect 4511 20502 4557 20554
rect 4581 20502 4627 20554
rect 4627 20502 4637 20554
rect 4661 20502 4691 20554
rect 4691 20502 4717 20554
rect 4421 20500 4477 20502
rect 4501 20500 4557 20502
rect 4581 20500 4637 20502
rect 4661 20500 4717 20502
rect 4421 19466 4477 19468
rect 4501 19466 4557 19468
rect 4581 19466 4637 19468
rect 4661 19466 4717 19468
rect 4421 19414 4447 19466
rect 4447 19414 4477 19466
rect 4501 19414 4511 19466
rect 4511 19414 4557 19466
rect 4581 19414 4627 19466
rect 4627 19414 4637 19466
rect 4661 19414 4691 19466
rect 4691 19414 4717 19466
rect 4421 19412 4477 19414
rect 4501 19412 4557 19414
rect 4581 19412 4637 19414
rect 4661 19412 4717 19414
rect 4421 18378 4477 18380
rect 4501 18378 4557 18380
rect 4581 18378 4637 18380
rect 4661 18378 4717 18380
rect 4421 18326 4447 18378
rect 4447 18326 4477 18378
rect 4501 18326 4511 18378
rect 4511 18326 4557 18378
rect 4581 18326 4627 18378
rect 4627 18326 4637 18378
rect 4661 18326 4691 18378
rect 4691 18326 4717 18378
rect 4421 18324 4477 18326
rect 4501 18324 4557 18326
rect 4581 18324 4637 18326
rect 4661 18324 4717 18326
rect 4421 17290 4477 17292
rect 4501 17290 4557 17292
rect 4581 17290 4637 17292
rect 4661 17290 4717 17292
rect 4421 17238 4447 17290
rect 4447 17238 4477 17290
rect 4501 17238 4511 17290
rect 4511 17238 4557 17290
rect 4581 17238 4627 17290
rect 4627 17238 4637 17290
rect 4661 17238 4691 17290
rect 4691 17238 4717 17290
rect 4421 17236 4477 17238
rect 4501 17236 4557 17238
rect 4581 17236 4637 17238
rect 4661 17236 4717 17238
rect 4066 17032 4122 17088
rect 4421 16202 4477 16204
rect 4501 16202 4557 16204
rect 4581 16202 4637 16204
rect 4661 16202 4717 16204
rect 4421 16150 4447 16202
rect 4447 16150 4477 16202
rect 4501 16150 4511 16202
rect 4511 16150 4557 16202
rect 4581 16150 4627 16202
rect 4627 16150 4637 16202
rect 4661 16150 4691 16202
rect 4691 16150 4717 16202
rect 4421 16148 4477 16150
rect 4501 16148 4557 16150
rect 4581 16148 4637 16150
rect 4661 16148 4717 16150
rect 4421 15114 4477 15116
rect 4501 15114 4557 15116
rect 4581 15114 4637 15116
rect 4661 15114 4717 15116
rect 4421 15062 4447 15114
rect 4447 15062 4477 15114
rect 4501 15062 4511 15114
rect 4511 15062 4557 15114
rect 4581 15062 4627 15114
rect 4627 15062 4637 15114
rect 4661 15062 4691 15114
rect 4691 15062 4717 15114
rect 4421 15060 4477 15062
rect 4501 15060 4557 15062
rect 4581 15060 4637 15062
rect 4661 15060 4717 15062
rect 4421 14026 4477 14028
rect 4501 14026 4557 14028
rect 4581 14026 4637 14028
rect 4661 14026 4717 14028
rect 4421 13974 4447 14026
rect 4447 13974 4477 14026
rect 4501 13974 4511 14026
rect 4511 13974 4557 14026
rect 4581 13974 4627 14026
rect 4627 13974 4637 14026
rect 4661 13974 4691 14026
rect 4691 13974 4717 14026
rect 4421 13972 4477 13974
rect 4501 13972 4557 13974
rect 4581 13972 4637 13974
rect 4661 13972 4717 13974
rect 6458 18664 6514 18720
rect 7886 20010 7942 20012
rect 7966 20010 8022 20012
rect 8046 20010 8102 20012
rect 8126 20010 8182 20012
rect 7886 19958 7912 20010
rect 7912 19958 7942 20010
rect 7966 19958 7976 20010
rect 7976 19958 8022 20010
rect 8046 19958 8092 20010
rect 8092 19958 8102 20010
rect 8126 19958 8156 20010
rect 8156 19958 8182 20010
rect 7886 19956 7942 19958
rect 7966 19956 8022 19958
rect 8046 19956 8102 19958
rect 8126 19956 8182 19958
rect 7886 18922 7942 18924
rect 7966 18922 8022 18924
rect 8046 18922 8102 18924
rect 8126 18922 8182 18924
rect 7886 18870 7912 18922
rect 7912 18870 7942 18922
rect 7966 18870 7976 18922
rect 7976 18870 8022 18922
rect 8046 18870 8092 18922
rect 8092 18870 8102 18922
rect 8126 18870 8156 18922
rect 8156 18870 8182 18922
rect 7886 18868 7942 18870
rect 7966 18868 8022 18870
rect 8046 18868 8102 18870
rect 8126 18868 8182 18870
rect 7654 18664 7710 18720
rect 7746 17984 7802 18040
rect 7886 17834 7942 17836
rect 7966 17834 8022 17836
rect 8046 17834 8102 17836
rect 8126 17834 8182 17836
rect 7886 17782 7912 17834
rect 7912 17782 7942 17834
rect 7966 17782 7976 17834
rect 7976 17782 8022 17834
rect 8046 17782 8092 17834
rect 8092 17782 8102 17834
rect 8126 17782 8156 17834
rect 8156 17782 8182 17834
rect 7886 17780 7942 17782
rect 7966 17780 8022 17782
rect 8046 17780 8102 17782
rect 8126 17780 8182 17782
rect 9770 19072 9826 19128
rect 10230 18664 10286 18720
rect 7886 16746 7942 16748
rect 7966 16746 8022 16748
rect 8046 16746 8102 16748
rect 8126 16746 8182 16748
rect 7886 16694 7912 16746
rect 7912 16694 7942 16746
rect 7966 16694 7976 16746
rect 7976 16694 8022 16746
rect 8046 16694 8092 16746
rect 8092 16694 8102 16746
rect 8126 16694 8156 16746
rect 8156 16694 8182 16746
rect 7886 16692 7942 16694
rect 7966 16692 8022 16694
rect 8046 16692 8102 16694
rect 8126 16692 8182 16694
rect 7886 15658 7942 15660
rect 7966 15658 8022 15660
rect 8046 15658 8102 15660
rect 8126 15658 8182 15660
rect 7886 15606 7912 15658
rect 7912 15606 7942 15658
rect 7966 15606 7976 15658
rect 7976 15606 8022 15658
rect 8046 15606 8092 15658
rect 8092 15606 8102 15658
rect 8126 15606 8156 15658
rect 8156 15606 8182 15658
rect 7886 15604 7942 15606
rect 7966 15604 8022 15606
rect 8046 15604 8102 15606
rect 8126 15604 8182 15606
rect 7886 14570 7942 14572
rect 7966 14570 8022 14572
rect 8046 14570 8102 14572
rect 8126 14570 8182 14572
rect 7886 14518 7912 14570
rect 7912 14518 7942 14570
rect 7966 14518 7976 14570
rect 7976 14518 8022 14570
rect 8046 14518 8092 14570
rect 8092 14518 8102 14570
rect 8126 14518 8156 14570
rect 8156 14518 8182 14570
rect 7886 14516 7942 14518
rect 7966 14516 8022 14518
rect 8046 14516 8102 14518
rect 8126 14516 8182 14518
rect 4421 12938 4477 12940
rect 4501 12938 4557 12940
rect 4581 12938 4637 12940
rect 4661 12938 4717 12940
rect 4421 12886 4447 12938
rect 4447 12886 4477 12938
rect 4501 12886 4511 12938
rect 4511 12886 4557 12938
rect 4581 12886 4627 12938
rect 4627 12886 4637 12938
rect 4661 12886 4691 12938
rect 4691 12886 4717 12938
rect 4421 12884 4477 12886
rect 4501 12884 4557 12886
rect 4581 12884 4637 12886
rect 4661 12884 4717 12886
rect 7886 13482 7942 13484
rect 7966 13482 8022 13484
rect 8046 13482 8102 13484
rect 8126 13482 8182 13484
rect 7886 13430 7912 13482
rect 7912 13430 7942 13482
rect 7966 13430 7976 13482
rect 7976 13430 8022 13482
rect 8046 13430 8092 13482
rect 8092 13430 8102 13482
rect 8126 13430 8156 13482
rect 8156 13430 8182 13482
rect 7886 13428 7942 13430
rect 7966 13428 8022 13430
rect 8046 13428 8102 13430
rect 8126 13428 8182 13430
rect 11352 20554 11408 20556
rect 11432 20554 11488 20556
rect 11512 20554 11568 20556
rect 11592 20554 11648 20556
rect 11352 20502 11378 20554
rect 11378 20502 11408 20554
rect 11432 20502 11442 20554
rect 11442 20502 11488 20554
rect 11512 20502 11558 20554
rect 11558 20502 11568 20554
rect 11592 20502 11622 20554
rect 11622 20502 11648 20554
rect 11352 20500 11408 20502
rect 11432 20500 11488 20502
rect 11512 20500 11568 20502
rect 11592 20500 11648 20502
rect 11426 19616 11482 19672
rect 11352 19466 11408 19468
rect 11432 19466 11488 19468
rect 11512 19466 11568 19468
rect 11592 19466 11648 19468
rect 11352 19414 11378 19466
rect 11378 19414 11408 19466
rect 11432 19414 11442 19466
rect 11442 19414 11488 19466
rect 11512 19414 11558 19466
rect 11558 19414 11568 19466
rect 11592 19414 11622 19466
rect 11622 19414 11648 19466
rect 11352 19412 11408 19414
rect 11432 19412 11488 19414
rect 11512 19412 11568 19414
rect 11592 19412 11648 19414
rect 11352 18378 11408 18380
rect 11432 18378 11488 18380
rect 11512 18378 11568 18380
rect 11592 18378 11648 18380
rect 11352 18326 11378 18378
rect 11378 18326 11408 18378
rect 11432 18326 11442 18378
rect 11442 18326 11488 18378
rect 11512 18326 11558 18378
rect 11558 18326 11568 18378
rect 11592 18326 11622 18378
rect 11622 18326 11648 18378
rect 11352 18324 11408 18326
rect 11432 18324 11488 18326
rect 11512 18324 11568 18326
rect 11592 18324 11648 18326
rect 11352 17290 11408 17292
rect 11432 17290 11488 17292
rect 11512 17290 11568 17292
rect 11592 17290 11648 17292
rect 11352 17238 11378 17290
rect 11378 17238 11408 17290
rect 11432 17238 11442 17290
rect 11442 17238 11488 17290
rect 11512 17238 11558 17290
rect 11558 17238 11568 17290
rect 11592 17238 11622 17290
rect 11622 17238 11648 17290
rect 11352 17236 11408 17238
rect 11432 17236 11488 17238
rect 11512 17236 11568 17238
rect 11592 17236 11648 17238
rect 11352 16202 11408 16204
rect 11432 16202 11488 16204
rect 11512 16202 11568 16204
rect 11592 16202 11648 16204
rect 11352 16150 11378 16202
rect 11378 16150 11408 16202
rect 11432 16150 11442 16202
rect 11442 16150 11488 16202
rect 11512 16150 11558 16202
rect 11558 16150 11568 16202
rect 11592 16150 11622 16202
rect 11622 16150 11648 16202
rect 11352 16148 11408 16150
rect 11432 16148 11488 16150
rect 11512 16148 11568 16150
rect 11592 16148 11648 16150
rect 11352 15114 11408 15116
rect 11432 15114 11488 15116
rect 11512 15114 11568 15116
rect 11592 15114 11648 15116
rect 11352 15062 11378 15114
rect 11378 15062 11408 15114
rect 11432 15062 11442 15114
rect 11442 15062 11488 15114
rect 11512 15062 11558 15114
rect 11558 15062 11568 15114
rect 11592 15062 11622 15114
rect 11622 15062 11648 15114
rect 11352 15060 11408 15062
rect 11432 15060 11488 15062
rect 11512 15060 11568 15062
rect 11592 15060 11648 15062
rect 9402 13088 9458 13144
rect 9586 13108 9642 13144
rect 9586 13088 9588 13108
rect 9588 13088 9640 13108
rect 9640 13088 9642 13108
rect 7886 12394 7942 12396
rect 7966 12394 8022 12396
rect 8046 12394 8102 12396
rect 8126 12394 8182 12396
rect 7886 12342 7912 12394
rect 7912 12342 7942 12394
rect 7966 12342 7976 12394
rect 7976 12342 8022 12394
rect 8046 12342 8092 12394
rect 8092 12342 8102 12394
rect 8126 12342 8156 12394
rect 8156 12342 8182 12394
rect 7886 12340 7942 12342
rect 7966 12340 8022 12342
rect 8046 12340 8102 12342
rect 8126 12340 8182 12342
rect 4421 11850 4477 11852
rect 4501 11850 4557 11852
rect 4581 11850 4637 11852
rect 4661 11850 4717 11852
rect 4421 11798 4447 11850
rect 4447 11798 4477 11850
rect 4501 11798 4511 11850
rect 4511 11798 4557 11850
rect 4581 11798 4627 11850
rect 4627 11798 4637 11850
rect 4661 11798 4691 11850
rect 4691 11798 4717 11850
rect 4421 11796 4477 11798
rect 4501 11796 4557 11798
rect 4581 11796 4637 11798
rect 4661 11796 4717 11798
rect 7886 11306 7942 11308
rect 7966 11306 8022 11308
rect 8046 11306 8102 11308
rect 8126 11306 8182 11308
rect 7886 11254 7912 11306
rect 7912 11254 7942 11306
rect 7966 11254 7976 11306
rect 7976 11254 8022 11306
rect 8046 11254 8092 11306
rect 8092 11254 8102 11306
rect 8126 11254 8156 11306
rect 8156 11254 8182 11306
rect 7886 11252 7942 11254
rect 7966 11252 8022 11254
rect 8046 11252 8102 11254
rect 8126 11252 8182 11254
rect 4421 10762 4477 10764
rect 4501 10762 4557 10764
rect 4581 10762 4637 10764
rect 4661 10762 4717 10764
rect 4421 10710 4447 10762
rect 4447 10710 4477 10762
rect 4501 10710 4511 10762
rect 4511 10710 4557 10762
rect 4581 10710 4627 10762
rect 4627 10710 4637 10762
rect 4661 10710 4691 10762
rect 4691 10710 4717 10762
rect 4421 10708 4477 10710
rect 4501 10708 4557 10710
rect 4581 10708 4637 10710
rect 4661 10708 4717 10710
rect 7886 10218 7942 10220
rect 7966 10218 8022 10220
rect 8046 10218 8102 10220
rect 8126 10218 8182 10220
rect 7886 10166 7912 10218
rect 7912 10166 7942 10218
rect 7966 10166 7976 10218
rect 7976 10166 8022 10218
rect 8046 10166 8092 10218
rect 8092 10166 8102 10218
rect 8126 10166 8156 10218
rect 8156 10166 8182 10218
rect 7886 10164 7942 10166
rect 7966 10164 8022 10166
rect 8046 10164 8102 10166
rect 8126 10164 8182 10166
rect 4421 9674 4477 9676
rect 4501 9674 4557 9676
rect 4581 9674 4637 9676
rect 4661 9674 4717 9676
rect 4421 9622 4447 9674
rect 4447 9622 4477 9674
rect 4501 9622 4511 9674
rect 4511 9622 4557 9674
rect 4581 9622 4627 9674
rect 4627 9622 4637 9674
rect 4661 9622 4691 9674
rect 4691 9622 4717 9674
rect 4421 9620 4477 9622
rect 4501 9620 4557 9622
rect 4581 9620 4637 9622
rect 4661 9620 4717 9622
rect 7886 9130 7942 9132
rect 7966 9130 8022 9132
rect 8046 9130 8102 9132
rect 8126 9130 8182 9132
rect 7886 9078 7912 9130
rect 7912 9078 7942 9130
rect 7966 9078 7976 9130
rect 7976 9078 8022 9130
rect 8046 9078 8092 9130
rect 8092 9078 8102 9130
rect 8126 9078 8156 9130
rect 8156 9078 8182 9130
rect 7886 9076 7942 9078
rect 7966 9076 8022 9078
rect 8046 9076 8102 9078
rect 8126 9076 8182 9078
rect 4421 8586 4477 8588
rect 4501 8586 4557 8588
rect 4581 8586 4637 8588
rect 4661 8586 4717 8588
rect 4421 8534 4447 8586
rect 4447 8534 4477 8586
rect 4501 8534 4511 8586
rect 4511 8534 4557 8586
rect 4581 8534 4627 8586
rect 4627 8534 4637 8586
rect 4661 8534 4691 8586
rect 4691 8534 4717 8586
rect 4421 8532 4477 8534
rect 4501 8532 4557 8534
rect 4581 8532 4637 8534
rect 4661 8532 4717 8534
rect 11352 14026 11408 14028
rect 11432 14026 11488 14028
rect 11512 14026 11568 14028
rect 11592 14026 11648 14028
rect 11352 13974 11378 14026
rect 11378 13974 11408 14026
rect 11432 13974 11442 14026
rect 11442 13974 11488 14026
rect 11512 13974 11558 14026
rect 11558 13974 11568 14026
rect 11592 13974 11622 14026
rect 11622 13974 11648 14026
rect 11352 13972 11408 13974
rect 11432 13972 11488 13974
rect 11512 13972 11568 13974
rect 11592 13972 11648 13974
rect 11352 12938 11408 12940
rect 11432 12938 11488 12940
rect 11512 12938 11568 12940
rect 11592 12938 11648 12940
rect 11352 12886 11378 12938
rect 11378 12886 11408 12938
rect 11432 12886 11442 12938
rect 11442 12886 11488 12938
rect 11512 12886 11558 12938
rect 11558 12886 11568 12938
rect 11592 12886 11622 12938
rect 11622 12886 11648 12938
rect 11352 12884 11408 12886
rect 11432 12884 11488 12886
rect 11512 12884 11568 12886
rect 11592 12884 11648 12886
rect 11352 11850 11408 11852
rect 11432 11850 11488 11852
rect 11512 11850 11568 11852
rect 11592 11850 11648 11852
rect 11352 11798 11378 11850
rect 11378 11798 11408 11850
rect 11432 11798 11442 11850
rect 11442 11798 11488 11850
rect 11512 11798 11558 11850
rect 11558 11798 11568 11850
rect 11592 11798 11622 11850
rect 11622 11798 11648 11850
rect 11352 11796 11408 11798
rect 11432 11796 11488 11798
rect 11512 11796 11568 11798
rect 11592 11796 11648 11798
rect 11352 10762 11408 10764
rect 11432 10762 11488 10764
rect 11512 10762 11568 10764
rect 11592 10762 11648 10764
rect 11352 10710 11378 10762
rect 11378 10710 11408 10762
rect 11432 10710 11442 10762
rect 11442 10710 11488 10762
rect 11512 10710 11558 10762
rect 11558 10710 11568 10762
rect 11592 10710 11622 10762
rect 11622 10710 11648 10762
rect 11352 10708 11408 10710
rect 11432 10708 11488 10710
rect 11512 10708 11568 10710
rect 11592 10708 11648 10710
rect 11352 9674 11408 9676
rect 11432 9674 11488 9676
rect 11512 9674 11568 9676
rect 11592 9674 11648 9676
rect 11352 9622 11378 9674
rect 11378 9622 11408 9674
rect 11432 9622 11442 9674
rect 11442 9622 11488 9674
rect 11512 9622 11558 9674
rect 11558 9622 11568 9674
rect 11592 9622 11622 9674
rect 11622 9622 11648 9674
rect 11352 9620 11408 9622
rect 11432 9620 11488 9622
rect 11512 9620 11568 9622
rect 11592 9620 11648 9622
rect 12346 19788 12348 19808
rect 12348 19788 12400 19808
rect 12400 19788 12402 19808
rect 12346 19752 12402 19788
rect 7886 8042 7942 8044
rect 7966 8042 8022 8044
rect 8046 8042 8102 8044
rect 8126 8042 8182 8044
rect 7886 7990 7912 8042
rect 7912 7990 7942 8042
rect 7966 7990 7976 8042
rect 7976 7990 8022 8042
rect 8046 7990 8092 8042
rect 8092 7990 8102 8042
rect 8126 7990 8156 8042
rect 8156 7990 8182 8042
rect 7886 7988 7942 7990
rect 7966 7988 8022 7990
rect 8046 7988 8102 7990
rect 8126 7988 8182 7990
rect 4421 7498 4477 7500
rect 4501 7498 4557 7500
rect 4581 7498 4637 7500
rect 4661 7498 4717 7500
rect 4421 7446 4447 7498
rect 4447 7446 4477 7498
rect 4501 7446 4511 7498
rect 4511 7446 4557 7498
rect 4581 7446 4627 7498
rect 4627 7446 4637 7498
rect 4661 7446 4691 7498
rect 4691 7446 4717 7498
rect 4421 7444 4477 7446
rect 4501 7444 4557 7446
rect 4581 7444 4637 7446
rect 4661 7444 4717 7446
rect 7886 6954 7942 6956
rect 7966 6954 8022 6956
rect 8046 6954 8102 6956
rect 8126 6954 8182 6956
rect 7886 6902 7912 6954
rect 7912 6902 7942 6954
rect 7966 6902 7976 6954
rect 7976 6902 8022 6954
rect 8046 6902 8092 6954
rect 8092 6902 8102 6954
rect 8126 6902 8156 6954
rect 8156 6902 8182 6954
rect 7886 6900 7942 6902
rect 7966 6900 8022 6902
rect 8046 6900 8102 6902
rect 8126 6900 8182 6902
rect 11352 8586 11408 8588
rect 11432 8586 11488 8588
rect 11512 8586 11568 8588
rect 11592 8586 11648 8588
rect 11352 8534 11378 8586
rect 11378 8534 11408 8586
rect 11432 8534 11442 8586
rect 11442 8534 11488 8586
rect 11512 8534 11558 8586
rect 11558 8534 11568 8586
rect 11592 8534 11622 8586
rect 11622 8534 11648 8586
rect 11352 8532 11408 8534
rect 11432 8532 11488 8534
rect 11512 8532 11568 8534
rect 11592 8532 11648 8534
rect 11352 7498 11408 7500
rect 11432 7498 11488 7500
rect 11512 7498 11568 7500
rect 11592 7498 11648 7500
rect 11352 7446 11378 7498
rect 11378 7446 11408 7498
rect 11432 7446 11442 7498
rect 11442 7446 11488 7498
rect 11512 7446 11558 7498
rect 11558 7446 11568 7498
rect 11592 7446 11622 7498
rect 11622 7446 11648 7498
rect 11352 7444 11408 7446
rect 11432 7444 11488 7446
rect 11512 7444 11568 7446
rect 11592 7444 11648 7446
rect 4421 6410 4477 6412
rect 4501 6410 4557 6412
rect 4581 6410 4637 6412
rect 4661 6410 4717 6412
rect 4421 6358 4447 6410
rect 4447 6358 4477 6410
rect 4501 6358 4511 6410
rect 4511 6358 4557 6410
rect 4581 6358 4627 6410
rect 4627 6358 4637 6410
rect 4661 6358 4691 6410
rect 4691 6358 4717 6410
rect 4421 6356 4477 6358
rect 4501 6356 4557 6358
rect 4581 6356 4637 6358
rect 4661 6356 4717 6358
rect 11352 6410 11408 6412
rect 11432 6410 11488 6412
rect 11512 6410 11568 6412
rect 11592 6410 11648 6412
rect 11352 6358 11378 6410
rect 11378 6358 11408 6410
rect 11432 6358 11442 6410
rect 11442 6358 11488 6410
rect 11512 6358 11558 6410
rect 11558 6358 11568 6410
rect 11592 6358 11622 6410
rect 11622 6358 11648 6410
rect 11352 6356 11408 6358
rect 11432 6356 11488 6358
rect 11512 6356 11568 6358
rect 11592 6356 11648 6358
rect 7886 5866 7942 5868
rect 7966 5866 8022 5868
rect 8046 5866 8102 5868
rect 8126 5866 8182 5868
rect 7886 5814 7912 5866
rect 7912 5814 7942 5866
rect 7966 5814 7976 5866
rect 7976 5814 8022 5866
rect 8046 5814 8092 5866
rect 8092 5814 8102 5866
rect 8126 5814 8156 5866
rect 8156 5814 8182 5866
rect 7886 5812 7942 5814
rect 7966 5812 8022 5814
rect 8046 5812 8102 5814
rect 8126 5812 8182 5814
rect 3698 5608 3754 5664
rect 4421 5322 4477 5324
rect 4501 5322 4557 5324
rect 4581 5322 4637 5324
rect 4661 5322 4717 5324
rect 4421 5270 4447 5322
rect 4447 5270 4477 5322
rect 4501 5270 4511 5322
rect 4511 5270 4557 5322
rect 4581 5270 4627 5322
rect 4627 5270 4637 5322
rect 4661 5270 4691 5322
rect 4691 5270 4717 5322
rect 4421 5268 4477 5270
rect 4501 5268 4557 5270
rect 4581 5268 4637 5270
rect 4661 5268 4717 5270
rect 11352 5322 11408 5324
rect 11432 5322 11488 5324
rect 11512 5322 11568 5324
rect 11592 5322 11648 5324
rect 11352 5270 11378 5322
rect 11378 5270 11408 5322
rect 11432 5270 11442 5322
rect 11442 5270 11488 5322
rect 11512 5270 11558 5322
rect 11558 5270 11568 5322
rect 11592 5270 11622 5322
rect 11622 5270 11648 5322
rect 11352 5268 11408 5270
rect 11432 5268 11488 5270
rect 11512 5268 11568 5270
rect 11592 5268 11648 5270
rect 7886 4778 7942 4780
rect 7966 4778 8022 4780
rect 8046 4778 8102 4780
rect 8126 4778 8182 4780
rect 7886 4726 7912 4778
rect 7912 4726 7942 4778
rect 7966 4726 7976 4778
rect 7976 4726 8022 4778
rect 8046 4726 8092 4778
rect 8092 4726 8102 4778
rect 8126 4726 8156 4778
rect 8156 4726 8182 4778
rect 7886 4724 7942 4726
rect 7966 4724 8022 4726
rect 8046 4724 8102 4726
rect 8126 4724 8182 4726
rect 14817 20010 14873 20012
rect 14897 20010 14953 20012
rect 14977 20010 15033 20012
rect 15057 20010 15113 20012
rect 14817 19958 14843 20010
rect 14843 19958 14873 20010
rect 14897 19958 14907 20010
rect 14907 19958 14953 20010
rect 14977 19958 15023 20010
rect 15023 19958 15033 20010
rect 15057 19958 15087 20010
rect 15087 19958 15113 20010
rect 14817 19956 14873 19958
rect 14897 19956 14953 19958
rect 14977 19956 15033 19958
rect 15057 19956 15113 19958
rect 15198 19908 15254 19944
rect 15198 19888 15200 19908
rect 15200 19888 15252 19908
rect 15252 19888 15254 19908
rect 15198 18936 15254 18992
rect 14817 18922 14873 18924
rect 14897 18922 14953 18924
rect 14977 18922 15033 18924
rect 15057 18922 15113 18924
rect 14817 18870 14843 18922
rect 14843 18870 14873 18922
rect 14897 18870 14907 18922
rect 14907 18870 14953 18922
rect 14977 18870 15023 18922
rect 15023 18870 15033 18922
rect 15057 18870 15087 18922
rect 15087 18870 15113 18922
rect 14817 18868 14873 18870
rect 14897 18868 14953 18870
rect 14977 18868 15033 18870
rect 15057 18868 15113 18870
rect 14738 18528 14794 18584
rect 4421 4234 4477 4236
rect 4501 4234 4557 4236
rect 4581 4234 4637 4236
rect 4661 4234 4717 4236
rect 4421 4182 4447 4234
rect 4447 4182 4477 4234
rect 4501 4182 4511 4234
rect 4511 4182 4557 4234
rect 4581 4182 4627 4234
rect 4627 4182 4637 4234
rect 4661 4182 4691 4234
rect 4691 4182 4717 4234
rect 4421 4180 4477 4182
rect 4501 4180 4557 4182
rect 4581 4180 4637 4182
rect 4661 4180 4717 4182
rect 11352 4234 11408 4236
rect 11432 4234 11488 4236
rect 11512 4234 11568 4236
rect 11592 4234 11648 4236
rect 11352 4182 11378 4234
rect 11378 4182 11408 4234
rect 11432 4182 11442 4234
rect 11442 4182 11488 4234
rect 11512 4182 11558 4234
rect 11558 4182 11568 4234
rect 11592 4182 11622 4234
rect 11622 4182 11648 4234
rect 11352 4180 11408 4182
rect 11432 4180 11488 4182
rect 11512 4180 11568 4182
rect 11592 4180 11648 4182
rect 14817 17834 14873 17836
rect 14897 17834 14953 17836
rect 14977 17834 15033 17836
rect 15057 17834 15113 17836
rect 14817 17782 14843 17834
rect 14843 17782 14873 17834
rect 14897 17782 14907 17834
rect 14907 17782 14953 17834
rect 14977 17782 15023 17834
rect 15023 17782 15033 17834
rect 15057 17782 15087 17834
rect 15087 17782 15113 17834
rect 14817 17780 14873 17782
rect 14897 17780 14953 17782
rect 14977 17780 15033 17782
rect 15057 17780 15113 17782
rect 14817 16746 14873 16748
rect 14897 16746 14953 16748
rect 14977 16746 15033 16748
rect 15057 16746 15113 16748
rect 14817 16694 14843 16746
rect 14843 16694 14873 16746
rect 14897 16694 14907 16746
rect 14907 16694 14953 16746
rect 14977 16694 15023 16746
rect 15023 16694 15033 16746
rect 15057 16694 15087 16746
rect 15087 16694 15113 16746
rect 14817 16692 14873 16694
rect 14897 16692 14953 16694
rect 14977 16692 15033 16694
rect 15057 16692 15113 16694
rect 14817 15658 14873 15660
rect 14897 15658 14953 15660
rect 14977 15658 15033 15660
rect 15057 15658 15113 15660
rect 14817 15606 14843 15658
rect 14843 15606 14873 15658
rect 14897 15606 14907 15658
rect 14907 15606 14953 15658
rect 14977 15606 15023 15658
rect 15023 15606 15033 15658
rect 15057 15606 15087 15658
rect 15087 15606 15113 15658
rect 14817 15604 14873 15606
rect 14897 15604 14953 15606
rect 14977 15604 15033 15606
rect 15057 15604 15113 15606
rect 14817 14570 14873 14572
rect 14897 14570 14953 14572
rect 14977 14570 15033 14572
rect 15057 14570 15113 14572
rect 14817 14518 14843 14570
rect 14843 14518 14873 14570
rect 14897 14518 14907 14570
rect 14907 14518 14953 14570
rect 14977 14518 15023 14570
rect 15023 14518 15033 14570
rect 15057 14518 15087 14570
rect 15087 14518 15113 14570
rect 14817 14516 14873 14518
rect 14897 14516 14953 14518
rect 14977 14516 15033 14518
rect 15057 14516 15113 14518
rect 14817 13482 14873 13484
rect 14897 13482 14953 13484
rect 14977 13482 15033 13484
rect 15057 13482 15113 13484
rect 14817 13430 14843 13482
rect 14843 13430 14873 13482
rect 14897 13430 14907 13482
rect 14907 13430 14953 13482
rect 14977 13430 15023 13482
rect 15023 13430 15033 13482
rect 15057 13430 15087 13482
rect 15087 13430 15113 13482
rect 14817 13428 14873 13430
rect 14897 13428 14953 13430
rect 14977 13428 15033 13430
rect 15057 13428 15113 13430
rect 14817 12394 14873 12396
rect 14897 12394 14953 12396
rect 14977 12394 15033 12396
rect 15057 12394 15113 12396
rect 14817 12342 14843 12394
rect 14843 12342 14873 12394
rect 14897 12342 14907 12394
rect 14907 12342 14953 12394
rect 14977 12342 15023 12394
rect 15023 12342 15033 12394
rect 15057 12342 15087 12394
rect 15087 12342 15113 12394
rect 14817 12340 14873 12342
rect 14897 12340 14953 12342
rect 14977 12340 15033 12342
rect 15057 12340 15113 12342
rect 14817 11306 14873 11308
rect 14897 11306 14953 11308
rect 14977 11306 15033 11308
rect 15057 11306 15113 11308
rect 14817 11254 14843 11306
rect 14843 11254 14873 11306
rect 14897 11254 14907 11306
rect 14907 11254 14953 11306
rect 14977 11254 15023 11306
rect 15023 11254 15033 11306
rect 15057 11254 15087 11306
rect 15087 11254 15113 11306
rect 14817 11252 14873 11254
rect 14897 11252 14953 11254
rect 14977 11252 15033 11254
rect 15057 11252 15113 11254
rect 16026 19908 16082 19944
rect 16026 19888 16028 19908
rect 16028 19888 16080 19908
rect 16080 19888 16082 19908
rect 14817 10218 14873 10220
rect 14897 10218 14953 10220
rect 14977 10218 15033 10220
rect 15057 10218 15113 10220
rect 14817 10166 14843 10218
rect 14843 10166 14873 10218
rect 14897 10166 14907 10218
rect 14907 10166 14953 10218
rect 14977 10166 15023 10218
rect 15023 10166 15033 10218
rect 15057 10166 15087 10218
rect 15087 10166 15113 10218
rect 14817 10164 14873 10166
rect 14897 10164 14953 10166
rect 14977 10164 15033 10166
rect 15057 10164 15113 10166
rect 14817 9130 14873 9132
rect 14897 9130 14953 9132
rect 14977 9130 15033 9132
rect 15057 9130 15113 9132
rect 14817 9078 14843 9130
rect 14843 9078 14873 9130
rect 14897 9078 14907 9130
rect 14907 9078 14953 9130
rect 14977 9078 15023 9130
rect 15023 9078 15033 9130
rect 15057 9078 15087 9130
rect 15087 9078 15113 9130
rect 14817 9076 14873 9078
rect 14897 9076 14953 9078
rect 14977 9076 15033 9078
rect 15057 9076 15113 9078
rect 14817 8042 14873 8044
rect 14897 8042 14953 8044
rect 14977 8042 15033 8044
rect 15057 8042 15113 8044
rect 14817 7990 14843 8042
rect 14843 7990 14873 8042
rect 14897 7990 14907 8042
rect 14907 7990 14953 8042
rect 14977 7990 15023 8042
rect 15023 7990 15033 8042
rect 15057 7990 15087 8042
rect 15087 7990 15113 8042
rect 14817 7988 14873 7990
rect 14897 7988 14953 7990
rect 14977 7988 15033 7990
rect 15057 7988 15113 7990
rect 14817 6954 14873 6956
rect 14897 6954 14953 6956
rect 14977 6954 15033 6956
rect 15057 6954 15113 6956
rect 14817 6902 14843 6954
rect 14843 6902 14873 6954
rect 14897 6902 14907 6954
rect 14907 6902 14953 6954
rect 14977 6902 15023 6954
rect 15023 6902 15033 6954
rect 15057 6902 15087 6954
rect 15087 6902 15113 6954
rect 14817 6900 14873 6902
rect 14897 6900 14953 6902
rect 14977 6900 15033 6902
rect 15057 6900 15113 6902
rect 14817 5866 14873 5868
rect 14897 5866 14953 5868
rect 14977 5866 15033 5868
rect 15057 5866 15113 5868
rect 14817 5814 14843 5866
rect 14843 5814 14873 5866
rect 14897 5814 14907 5866
rect 14907 5814 14953 5866
rect 14977 5814 15023 5866
rect 15023 5814 15033 5866
rect 15057 5814 15087 5866
rect 15087 5814 15113 5866
rect 14817 5812 14873 5814
rect 14897 5812 14953 5814
rect 14977 5812 15033 5814
rect 15057 5812 15113 5814
rect 14817 4778 14873 4780
rect 14897 4778 14953 4780
rect 14977 4778 15033 4780
rect 15057 4778 15113 4780
rect 14817 4726 14843 4778
rect 14843 4726 14873 4778
rect 14897 4726 14907 4778
rect 14907 4726 14953 4778
rect 14977 4726 15023 4778
rect 15023 4726 15033 4778
rect 15057 4726 15087 4778
rect 15087 4726 15113 4778
rect 14817 4724 14873 4726
rect 14897 4724 14953 4726
rect 14977 4724 15033 4726
rect 15057 4724 15113 4726
rect 7886 3690 7942 3692
rect 7966 3690 8022 3692
rect 8046 3690 8102 3692
rect 8126 3690 8182 3692
rect 7886 3638 7912 3690
rect 7912 3638 7942 3690
rect 7966 3638 7976 3690
rect 7976 3638 8022 3690
rect 8046 3638 8092 3690
rect 8092 3638 8102 3690
rect 8126 3638 8156 3690
rect 8156 3638 8182 3690
rect 7886 3636 7942 3638
rect 7966 3636 8022 3638
rect 8046 3636 8102 3638
rect 8126 3636 8182 3638
rect 14817 3690 14873 3692
rect 14897 3690 14953 3692
rect 14977 3690 15033 3692
rect 15057 3690 15113 3692
rect 14817 3638 14843 3690
rect 14843 3638 14873 3690
rect 14897 3638 14907 3690
rect 14907 3638 14953 3690
rect 14977 3638 15023 3690
rect 15023 3638 15033 3690
rect 15057 3638 15087 3690
rect 15087 3638 15113 3690
rect 14817 3636 14873 3638
rect 14897 3636 14953 3638
rect 14977 3636 15033 3638
rect 15057 3636 15113 3638
rect 4421 3146 4477 3148
rect 4501 3146 4557 3148
rect 4581 3146 4637 3148
rect 4661 3146 4717 3148
rect 4421 3094 4447 3146
rect 4447 3094 4477 3146
rect 4501 3094 4511 3146
rect 4511 3094 4557 3146
rect 4581 3094 4627 3146
rect 4627 3094 4637 3146
rect 4661 3094 4691 3146
rect 4691 3094 4717 3146
rect 4421 3092 4477 3094
rect 4501 3092 4557 3094
rect 4581 3092 4637 3094
rect 4661 3092 4717 3094
rect 11352 3146 11408 3148
rect 11432 3146 11488 3148
rect 11512 3146 11568 3148
rect 11592 3146 11648 3148
rect 11352 3094 11378 3146
rect 11378 3094 11408 3146
rect 11432 3094 11442 3146
rect 11442 3094 11488 3146
rect 11512 3094 11558 3146
rect 11558 3094 11568 3146
rect 11592 3094 11622 3146
rect 11622 3094 11648 3146
rect 11352 3092 11408 3094
rect 11432 3092 11488 3094
rect 11512 3092 11568 3094
rect 11592 3092 11648 3094
rect 7886 2602 7942 2604
rect 7966 2602 8022 2604
rect 8046 2602 8102 2604
rect 8126 2602 8182 2604
rect 7886 2550 7912 2602
rect 7912 2550 7942 2602
rect 7966 2550 7976 2602
rect 7976 2550 8022 2602
rect 8046 2550 8092 2602
rect 8092 2550 8102 2602
rect 8126 2550 8156 2602
rect 8156 2550 8182 2602
rect 7886 2548 7942 2550
rect 7966 2548 8022 2550
rect 8046 2548 8102 2550
rect 8126 2548 8182 2550
rect 14817 2602 14873 2604
rect 14897 2602 14953 2604
rect 14977 2602 15033 2604
rect 15057 2602 15113 2604
rect 14817 2550 14843 2602
rect 14843 2550 14873 2602
rect 14897 2550 14907 2602
rect 14907 2550 14953 2602
rect 14977 2550 15023 2602
rect 15023 2550 15033 2602
rect 15057 2550 15087 2602
rect 15087 2550 15113 2602
rect 14817 2548 14873 2550
rect 14897 2548 14953 2550
rect 14977 2548 15033 2550
rect 15057 2548 15113 2550
rect 4421 2058 4477 2060
rect 4501 2058 4557 2060
rect 4581 2058 4637 2060
rect 4661 2058 4717 2060
rect 4421 2006 4447 2058
rect 4447 2006 4477 2058
rect 4501 2006 4511 2058
rect 4511 2006 4557 2058
rect 4581 2006 4627 2058
rect 4627 2006 4637 2058
rect 4661 2006 4691 2058
rect 4691 2006 4717 2058
rect 4421 2004 4477 2006
rect 4501 2004 4557 2006
rect 4581 2004 4637 2006
rect 4661 2004 4717 2006
rect 11352 2058 11408 2060
rect 11432 2058 11488 2060
rect 11512 2058 11568 2060
rect 11592 2058 11648 2060
rect 11352 2006 11378 2058
rect 11378 2006 11408 2058
rect 11432 2006 11442 2058
rect 11442 2006 11488 2058
rect 11512 2006 11558 2058
rect 11558 2006 11568 2058
rect 11592 2006 11622 2058
rect 11622 2006 11648 2058
rect 11352 2004 11408 2006
rect 11432 2004 11488 2006
rect 11512 2004 11568 2006
rect 11592 2004 11648 2006
rect 16394 19752 16450 19808
rect 17590 19752 17646 19808
rect 16762 18936 16818 18992
rect 18142 21928 18198 21984
rect 17866 20976 17922 21032
rect 18050 19616 18106 19672
rect 17682 19072 17738 19128
rect 17498 18664 17554 18720
rect 18282 20554 18338 20556
rect 18362 20554 18418 20556
rect 18442 20554 18498 20556
rect 18522 20554 18578 20556
rect 18282 20502 18308 20554
rect 18308 20502 18338 20554
rect 18362 20502 18372 20554
rect 18372 20502 18418 20554
rect 18442 20502 18488 20554
rect 18488 20502 18498 20554
rect 18522 20502 18552 20554
rect 18552 20502 18578 20554
rect 18282 20500 18338 20502
rect 18362 20500 18418 20502
rect 18442 20500 18498 20502
rect 18522 20500 18578 20502
rect 18282 19466 18338 19468
rect 18362 19466 18418 19468
rect 18442 19466 18498 19468
rect 18522 19466 18578 19468
rect 18282 19414 18308 19466
rect 18308 19414 18338 19466
rect 18362 19414 18372 19466
rect 18372 19414 18418 19466
rect 18442 19414 18488 19466
rect 18488 19414 18498 19466
rect 18522 19414 18552 19466
rect 18552 19414 18578 19466
rect 18282 19412 18338 19414
rect 18362 19412 18418 19414
rect 18442 19412 18498 19414
rect 18522 19412 18578 19414
rect 17958 18120 18014 18176
rect 18510 18936 18566 18992
rect 18418 18684 18474 18720
rect 18418 18664 18420 18684
rect 18420 18664 18472 18684
rect 18472 18664 18474 18684
rect 18234 18528 18290 18584
rect 18602 18528 18658 18584
rect 18282 18378 18338 18380
rect 18362 18378 18418 18380
rect 18442 18378 18498 18380
rect 18522 18378 18578 18380
rect 18282 18326 18308 18378
rect 18308 18326 18338 18378
rect 18362 18326 18372 18378
rect 18372 18326 18418 18378
rect 18442 18326 18488 18378
rect 18488 18326 18498 18378
rect 18522 18326 18552 18378
rect 18552 18326 18578 18378
rect 18282 18324 18338 18326
rect 18362 18324 18418 18326
rect 18442 18324 18498 18326
rect 18522 18324 18578 18326
rect 18282 17290 18338 17292
rect 18362 17290 18418 17292
rect 18442 17290 18498 17292
rect 18522 17290 18578 17292
rect 18282 17238 18308 17290
rect 18308 17238 18338 17290
rect 18362 17238 18372 17290
rect 18372 17238 18418 17290
rect 18442 17238 18488 17290
rect 18488 17238 18498 17290
rect 18522 17238 18552 17290
rect 18552 17238 18578 17290
rect 18282 17236 18338 17238
rect 18362 17236 18418 17238
rect 18442 17236 18498 17238
rect 18522 17236 18578 17238
rect 18970 20568 19026 20624
rect 18878 20024 18934 20080
rect 19154 21520 19210 21576
rect 18050 17032 18106 17088
rect 17958 16624 18014 16680
rect 17958 14176 18014 14232
rect 18602 16896 18658 16952
rect 18282 16202 18338 16204
rect 18362 16202 18418 16204
rect 18442 16202 18498 16204
rect 18522 16202 18578 16204
rect 18282 16150 18308 16202
rect 18308 16150 18338 16202
rect 18362 16150 18372 16202
rect 18372 16150 18418 16202
rect 18442 16150 18488 16202
rect 18488 16150 18498 16202
rect 18522 16150 18552 16202
rect 18552 16150 18578 16202
rect 18282 16148 18338 16150
rect 18362 16148 18418 16150
rect 18442 16148 18498 16150
rect 18522 16148 18578 16150
rect 18282 15114 18338 15116
rect 18362 15114 18418 15116
rect 18442 15114 18498 15116
rect 18522 15114 18578 15116
rect 18282 15062 18308 15114
rect 18308 15062 18338 15114
rect 18362 15062 18372 15114
rect 18372 15062 18418 15114
rect 18442 15062 18488 15114
rect 18488 15062 18498 15114
rect 18522 15062 18552 15114
rect 18552 15062 18578 15114
rect 18282 15060 18338 15062
rect 18362 15060 18418 15062
rect 18442 15060 18498 15062
rect 18522 15060 18578 15062
rect 18694 15128 18750 15184
rect 18602 14620 18604 14640
rect 18604 14620 18656 14640
rect 18656 14620 18658 14640
rect 18602 14584 18658 14620
rect 18282 14026 18338 14028
rect 18362 14026 18418 14028
rect 18442 14026 18498 14028
rect 18522 14026 18578 14028
rect 18282 13974 18308 14026
rect 18308 13974 18338 14026
rect 18362 13974 18372 14026
rect 18372 13974 18418 14026
rect 18442 13974 18488 14026
rect 18488 13974 18498 14026
rect 18522 13974 18552 14026
rect 18552 13974 18578 14026
rect 18282 13972 18338 13974
rect 18362 13972 18418 13974
rect 18442 13972 18498 13974
rect 18522 13972 18578 13974
rect 18282 12938 18338 12940
rect 18362 12938 18418 12940
rect 18442 12938 18498 12940
rect 18522 12938 18578 12940
rect 18282 12886 18308 12938
rect 18308 12886 18338 12938
rect 18362 12886 18372 12938
rect 18372 12886 18418 12938
rect 18442 12886 18488 12938
rect 18488 12886 18498 12938
rect 18522 12886 18552 12938
rect 18552 12886 18578 12938
rect 18282 12884 18338 12886
rect 18362 12884 18418 12886
rect 18442 12884 18498 12886
rect 18522 12884 18578 12886
rect 19246 17576 19302 17632
rect 19154 16080 19210 16136
rect 19246 15672 19302 15728
rect 18418 12172 18420 12192
rect 18420 12172 18472 12192
rect 18472 12172 18474 12192
rect 18418 12136 18474 12172
rect 18282 11850 18338 11852
rect 18362 11850 18418 11852
rect 18442 11850 18498 11852
rect 18522 11850 18578 11852
rect 18282 11798 18308 11850
rect 18308 11798 18338 11850
rect 18362 11798 18372 11850
rect 18372 11798 18418 11850
rect 18442 11798 18488 11850
rect 18488 11798 18498 11850
rect 18522 11798 18552 11850
rect 18552 11798 18578 11850
rect 18282 11796 18338 11798
rect 18362 11796 18418 11798
rect 18442 11796 18498 11798
rect 18522 11796 18578 11798
rect 17958 11184 18014 11240
rect 18282 10762 18338 10764
rect 18362 10762 18418 10764
rect 18442 10762 18498 10764
rect 18522 10762 18578 10764
rect 18282 10710 18308 10762
rect 18308 10710 18338 10762
rect 18362 10710 18372 10762
rect 18372 10710 18418 10762
rect 18442 10710 18488 10762
rect 18488 10710 18498 10762
rect 18522 10710 18552 10762
rect 18552 10710 18578 10762
rect 18282 10708 18338 10710
rect 18362 10708 18418 10710
rect 18442 10708 18498 10710
rect 18522 10708 18578 10710
rect 18282 9674 18338 9676
rect 18362 9674 18418 9676
rect 18442 9674 18498 9676
rect 18522 9674 18578 9676
rect 18282 9622 18308 9674
rect 18308 9622 18338 9674
rect 18362 9622 18372 9674
rect 18372 9622 18418 9674
rect 18442 9622 18488 9674
rect 18488 9622 18498 9674
rect 18522 9622 18552 9674
rect 18552 9622 18578 9674
rect 18282 9620 18338 9622
rect 18362 9620 18418 9622
rect 18442 9620 18498 9622
rect 18522 9620 18578 9622
rect 18282 8586 18338 8588
rect 18362 8586 18418 8588
rect 18442 8586 18498 8588
rect 18522 8586 18578 8588
rect 18282 8534 18308 8586
rect 18308 8534 18338 8586
rect 18362 8534 18372 8586
rect 18372 8534 18418 8586
rect 18442 8534 18488 8586
rect 18488 8534 18498 8586
rect 18522 8534 18552 8586
rect 18552 8534 18578 8586
rect 18282 8532 18338 8534
rect 18362 8532 18418 8534
rect 18442 8532 18498 8534
rect 18522 8532 18578 8534
rect 18282 7498 18338 7500
rect 18362 7498 18418 7500
rect 18442 7498 18498 7500
rect 18522 7498 18578 7500
rect 18282 7446 18308 7498
rect 18308 7446 18338 7498
rect 18362 7446 18372 7498
rect 18372 7446 18418 7498
rect 18442 7446 18488 7498
rect 18488 7446 18498 7498
rect 18522 7446 18552 7498
rect 18552 7446 18578 7498
rect 18282 7444 18338 7446
rect 18362 7444 18418 7446
rect 18442 7444 18498 7446
rect 18522 7444 18578 7446
rect 18282 6410 18338 6412
rect 18362 6410 18418 6412
rect 18442 6410 18498 6412
rect 18522 6410 18578 6412
rect 18282 6358 18308 6410
rect 18308 6358 18338 6410
rect 18362 6358 18372 6410
rect 18372 6358 18418 6410
rect 18442 6358 18488 6410
rect 18488 6358 18498 6410
rect 18522 6358 18552 6410
rect 18552 6358 18578 6410
rect 18282 6356 18338 6358
rect 18362 6356 18418 6358
rect 18442 6356 18498 6358
rect 18522 6356 18578 6358
rect 18282 5322 18338 5324
rect 18362 5322 18418 5324
rect 18442 5322 18498 5324
rect 18522 5322 18578 5324
rect 18282 5270 18308 5322
rect 18308 5270 18338 5322
rect 18362 5270 18372 5322
rect 18372 5270 18418 5322
rect 18442 5270 18488 5322
rect 18488 5270 18498 5322
rect 18522 5270 18552 5322
rect 18552 5270 18578 5322
rect 18282 5268 18338 5270
rect 18362 5268 18418 5270
rect 18442 5268 18498 5270
rect 18522 5268 18578 5270
rect 17958 4384 18014 4440
rect 18282 4234 18338 4236
rect 18362 4234 18418 4236
rect 18442 4234 18498 4236
rect 18522 4234 18578 4236
rect 18282 4182 18308 4234
rect 18308 4182 18338 4234
rect 18362 4182 18372 4234
rect 18372 4182 18418 4234
rect 18442 4182 18488 4234
rect 18488 4182 18498 4234
rect 18522 4182 18552 4234
rect 18552 4182 18578 4234
rect 18282 4180 18338 4182
rect 18362 4180 18418 4182
rect 18442 4180 18498 4182
rect 18522 4180 18578 4182
rect 17958 3840 18014 3896
rect 18050 3432 18106 3488
rect 18282 3146 18338 3148
rect 18362 3146 18418 3148
rect 18442 3146 18498 3148
rect 18522 3146 18578 3148
rect 18282 3094 18308 3146
rect 18308 3094 18338 3146
rect 18362 3094 18372 3146
rect 18372 3094 18418 3146
rect 18442 3094 18488 3146
rect 18488 3094 18498 3146
rect 18522 3094 18552 3146
rect 18552 3094 18578 3146
rect 18282 3092 18338 3094
rect 18362 3092 18418 3094
rect 18442 3092 18498 3094
rect 18522 3092 18578 3094
rect 18282 2058 18338 2060
rect 18362 2058 18418 2060
rect 18442 2058 18498 2060
rect 18522 2058 18578 2060
rect 18282 2006 18308 2058
rect 18308 2006 18338 2058
rect 18362 2006 18372 2058
rect 18372 2006 18418 2058
rect 18442 2006 18488 2058
rect 18488 2006 18498 2058
rect 18522 2006 18552 2058
rect 18552 2006 18578 2058
rect 18282 2004 18338 2006
rect 18362 2004 18418 2006
rect 18442 2004 18498 2006
rect 18522 2004 18578 2006
rect 19430 14876 19486 14912
rect 19430 14856 19432 14876
rect 19432 14856 19484 14876
rect 19484 14856 19486 14876
rect 19338 14740 19394 14776
rect 19338 14720 19340 14740
rect 19340 14720 19392 14740
rect 19392 14720 19394 14740
rect 18694 11728 18750 11784
rect 18878 9280 18934 9336
rect 18694 5336 18750 5392
rect 18602 1392 18658 1448
rect 18878 440 18934 496
rect 19246 9688 19302 9744
rect 19706 14876 19762 14912
rect 19706 14856 19708 14876
rect 19708 14856 19760 14876
rect 19760 14856 19762 14876
rect 19614 12680 19670 12736
rect 19706 10776 19762 10832
rect 19890 17984 19946 18040
rect 19982 14720 20038 14776
rect 20718 13632 20774 13688
rect 20626 13224 20682 13280
rect 20350 10232 20406 10288
rect 20534 8736 20590 8792
rect 19246 8328 19302 8384
rect 20626 7784 20682 7840
rect 19246 7240 19302 7296
rect 20534 6832 20590 6888
rect 19246 6288 19302 6344
rect 20534 5880 20590 5936
rect 20534 4792 20590 4848
rect 20534 2888 20590 2944
rect 19154 2344 19210 2400
rect 19246 1936 19302 1992
rect 19246 984 19302 1040
rect 18970 32 19026 88
<< metal3 >>
rect 19057 22530 19123 22533
rect 22520 22530 23000 22560
rect 19057 22528 23000 22530
rect 19057 22472 19062 22528
rect 19118 22472 23000 22528
rect 19057 22470 23000 22472
rect 19057 22467 19123 22470
rect 22520 22440 23000 22470
rect 18137 21986 18203 21989
rect 22520 21986 23000 22016
rect 18137 21984 23000 21986
rect 18137 21928 18142 21984
rect 18198 21928 23000 21984
rect 18137 21926 23000 21928
rect 18137 21923 18203 21926
rect 22520 21896 23000 21926
rect 19149 21578 19215 21581
rect 22520 21578 23000 21608
rect 19149 21576 23000 21578
rect 19149 21520 19154 21576
rect 19210 21520 23000 21576
rect 19149 21518 23000 21520
rect 19149 21515 19215 21518
rect 22520 21488 23000 21518
rect 17861 21034 17927 21037
rect 22520 21034 23000 21064
rect 17861 21032 23000 21034
rect 17861 20976 17866 21032
rect 17922 20976 23000 21032
rect 17861 20974 23000 20976
rect 17861 20971 17927 20974
rect 22520 20944 23000 20974
rect 18965 20626 19031 20629
rect 22520 20626 23000 20656
rect 18965 20624 23000 20626
rect 18965 20568 18970 20624
rect 19026 20568 23000 20624
rect 18965 20566 23000 20568
rect 18965 20563 19031 20566
rect 4409 20560 4729 20561
rect 4409 20496 4417 20560
rect 4481 20496 4497 20560
rect 4561 20496 4577 20560
rect 4641 20496 4657 20560
rect 4721 20496 4729 20560
rect 4409 20495 4729 20496
rect 11340 20560 11660 20561
rect 11340 20496 11348 20560
rect 11412 20496 11428 20560
rect 11492 20496 11508 20560
rect 11572 20496 11588 20560
rect 11652 20496 11660 20560
rect 11340 20495 11660 20496
rect 18270 20560 18590 20561
rect 18270 20496 18278 20560
rect 18342 20496 18358 20560
rect 18422 20496 18438 20560
rect 18502 20496 18518 20560
rect 18582 20496 18590 20560
rect 22520 20536 23000 20566
rect 18270 20495 18590 20496
rect 18873 20082 18939 20085
rect 22520 20082 23000 20112
rect 18873 20080 23000 20082
rect 18873 20024 18878 20080
rect 18934 20024 23000 20080
rect 18873 20022 23000 20024
rect 18873 20019 18939 20022
rect 7874 20016 8194 20017
rect 7874 19952 7882 20016
rect 7946 19952 7962 20016
rect 8026 19952 8042 20016
rect 8106 19952 8122 20016
rect 8186 19952 8194 20016
rect 7874 19951 8194 19952
rect 14805 20016 15125 20017
rect 14805 19952 14813 20016
rect 14877 19952 14893 20016
rect 14957 19952 14973 20016
rect 15037 19952 15053 20016
rect 15117 19952 15125 20016
rect 22520 19992 23000 20022
rect 14805 19951 15125 19952
rect 15193 19946 15259 19949
rect 16021 19946 16087 19949
rect 15193 19944 16087 19946
rect 15193 19888 15198 19944
rect 15254 19888 16026 19944
rect 16082 19888 16087 19944
rect 15193 19886 16087 19888
rect 15193 19883 15259 19886
rect 16021 19883 16087 19886
rect 12341 19810 12407 19813
rect 16389 19810 16455 19813
rect 12341 19808 16455 19810
rect 12341 19752 12346 19808
rect 12402 19752 16394 19808
rect 16450 19752 16455 19808
rect 12341 19750 16455 19752
rect 12341 19747 12407 19750
rect 16389 19747 16455 19750
rect 17585 19810 17651 19813
rect 17585 19808 18844 19810
rect 17585 19752 17590 19808
rect 17646 19752 18844 19808
rect 17585 19750 18844 19752
rect 17585 19747 17651 19750
rect 11421 19674 11487 19677
rect 18045 19674 18111 19677
rect 11421 19672 18111 19674
rect 11421 19616 11426 19672
rect 11482 19616 18050 19672
rect 18106 19616 18111 19672
rect 11421 19614 18111 19616
rect 11421 19611 11487 19614
rect 18045 19611 18111 19614
rect 18784 19538 18844 19750
rect 22520 19538 23000 19568
rect 18784 19478 23000 19538
rect 4409 19472 4729 19473
rect 4409 19408 4417 19472
rect 4481 19408 4497 19472
rect 4561 19408 4577 19472
rect 4641 19408 4657 19472
rect 4721 19408 4729 19472
rect 4409 19407 4729 19408
rect 11340 19472 11660 19473
rect 11340 19408 11348 19472
rect 11412 19408 11428 19472
rect 11492 19408 11508 19472
rect 11572 19408 11588 19472
rect 11652 19408 11660 19472
rect 11340 19407 11660 19408
rect 18270 19472 18590 19473
rect 18270 19408 18278 19472
rect 18342 19408 18358 19472
rect 18422 19408 18438 19472
rect 18502 19408 18518 19472
rect 18582 19408 18590 19472
rect 22520 19448 23000 19478
rect 18270 19407 18590 19408
rect 9765 19130 9831 19133
rect 17677 19130 17743 19133
rect 22520 19130 23000 19160
rect 9765 19128 17602 19130
rect 9765 19072 9770 19128
rect 9826 19072 17602 19128
rect 9765 19070 17602 19072
rect 9765 19067 9831 19070
rect 15193 18994 15259 18997
rect 16757 18994 16823 18997
rect 15193 18992 16823 18994
rect 15193 18936 15198 18992
rect 15254 18936 16762 18992
rect 16818 18936 16823 18992
rect 15193 18934 16823 18936
rect 17542 18994 17602 19070
rect 17677 19128 23000 19130
rect 17677 19072 17682 19128
rect 17738 19072 23000 19128
rect 17677 19070 23000 19072
rect 17677 19067 17743 19070
rect 22520 19040 23000 19070
rect 18505 18994 18571 18997
rect 17542 18992 18571 18994
rect 17542 18936 18510 18992
rect 18566 18936 18571 18992
rect 17542 18934 18571 18936
rect 15193 18931 15259 18934
rect 16757 18931 16823 18934
rect 18505 18931 18571 18934
rect 7874 18928 8194 18929
rect 7874 18864 7882 18928
rect 7946 18864 7962 18928
rect 8026 18864 8042 18928
rect 8106 18864 8122 18928
rect 8186 18864 8194 18928
rect 7874 18863 8194 18864
rect 14805 18928 15125 18929
rect 14805 18864 14813 18928
rect 14877 18864 14893 18928
rect 14957 18864 14973 18928
rect 15037 18864 15053 18928
rect 15117 18864 15125 18928
rect 14805 18863 15125 18864
rect 6453 18722 6519 18725
rect 7649 18722 7715 18725
rect 6453 18720 7715 18722
rect 6453 18664 6458 18720
rect 6514 18664 7654 18720
rect 7710 18664 7715 18720
rect 6453 18662 7715 18664
rect 6453 18659 6519 18662
rect 7649 18659 7715 18662
rect 10225 18722 10291 18725
rect 17493 18722 17559 18725
rect 10225 18720 17559 18722
rect 10225 18664 10230 18720
rect 10286 18664 17498 18720
rect 17554 18664 17559 18720
rect 10225 18662 17559 18664
rect 10225 18659 10291 18662
rect 17493 18659 17559 18662
rect 18413 18722 18479 18725
rect 18822 18722 18828 18724
rect 18413 18720 18828 18722
rect 18413 18664 18418 18720
rect 18474 18664 18828 18720
rect 18413 18662 18828 18664
rect 18413 18659 18479 18662
rect 18822 18660 18828 18662
rect 18892 18660 18898 18724
rect 14733 18586 14799 18589
rect 18229 18586 18295 18589
rect 14733 18584 18295 18586
rect 14733 18528 14738 18584
rect 14794 18528 18234 18584
rect 18290 18528 18295 18584
rect 14733 18526 18295 18528
rect 14733 18523 14799 18526
rect 18229 18523 18295 18526
rect 18597 18586 18663 18589
rect 22520 18586 23000 18616
rect 18597 18584 23000 18586
rect 18597 18528 18602 18584
rect 18658 18528 23000 18584
rect 18597 18526 23000 18528
rect 18597 18523 18663 18526
rect 22520 18496 23000 18526
rect 4409 18384 4729 18385
rect 4409 18320 4417 18384
rect 4481 18320 4497 18384
rect 4561 18320 4577 18384
rect 4641 18320 4657 18384
rect 4721 18320 4729 18384
rect 4409 18319 4729 18320
rect 11340 18384 11660 18385
rect 11340 18320 11348 18384
rect 11412 18320 11428 18384
rect 11492 18320 11508 18384
rect 11572 18320 11588 18384
rect 11652 18320 11660 18384
rect 11340 18319 11660 18320
rect 18270 18384 18590 18385
rect 18270 18320 18278 18384
rect 18342 18320 18358 18384
rect 18422 18320 18438 18384
rect 18502 18320 18518 18384
rect 18582 18320 18590 18384
rect 18270 18319 18590 18320
rect 17953 18178 18019 18181
rect 22520 18178 23000 18208
rect 17953 18176 23000 18178
rect 17953 18120 17958 18176
rect 18014 18120 23000 18176
rect 17953 18118 23000 18120
rect 17953 18115 18019 18118
rect 22520 18088 23000 18118
rect 7741 18042 7807 18045
rect 19885 18042 19951 18045
rect 7741 18040 19951 18042
rect 7741 17984 7746 18040
rect 7802 17984 19890 18040
rect 19946 17984 19951 18040
rect 7741 17982 19951 17984
rect 7741 17979 7807 17982
rect 19885 17979 19951 17982
rect 7874 17840 8194 17841
rect 7874 17776 7882 17840
rect 7946 17776 7962 17840
rect 8026 17776 8042 17840
rect 8106 17776 8122 17840
rect 8186 17776 8194 17840
rect 7874 17775 8194 17776
rect 14805 17840 15125 17841
rect 14805 17776 14813 17840
rect 14877 17776 14893 17840
rect 14957 17776 14973 17840
rect 15037 17776 15053 17840
rect 15117 17776 15125 17840
rect 14805 17775 15125 17776
rect 19241 17634 19307 17637
rect 22520 17634 23000 17664
rect 19241 17632 23000 17634
rect 19241 17576 19246 17632
rect 19302 17576 23000 17632
rect 19241 17574 23000 17576
rect 19241 17571 19307 17574
rect 22520 17544 23000 17574
rect 4409 17296 4729 17297
rect 4409 17232 4417 17296
rect 4481 17232 4497 17296
rect 4561 17232 4577 17296
rect 4641 17232 4657 17296
rect 4721 17232 4729 17296
rect 4409 17231 4729 17232
rect 11340 17296 11660 17297
rect 11340 17232 11348 17296
rect 11412 17232 11428 17296
rect 11492 17232 11508 17296
rect 11572 17232 11588 17296
rect 11652 17232 11660 17296
rect 11340 17231 11660 17232
rect 18270 17296 18590 17297
rect 18270 17232 18278 17296
rect 18342 17232 18358 17296
rect 18422 17232 18438 17296
rect 18502 17232 18518 17296
rect 18582 17232 18590 17296
rect 18270 17231 18590 17232
rect 0 17090 480 17120
rect 4061 17090 4127 17093
rect 0 17088 4127 17090
rect 0 17032 4066 17088
rect 4122 17032 4127 17088
rect 0 17030 4127 17032
rect 0 17000 480 17030
rect 4061 17027 4127 17030
rect 18045 17090 18111 17093
rect 22520 17090 23000 17120
rect 18045 17088 23000 17090
rect 18045 17032 18050 17088
rect 18106 17032 23000 17088
rect 18045 17030 23000 17032
rect 18045 17027 18111 17030
rect 22520 17000 23000 17030
rect 18597 16954 18663 16957
rect 18822 16954 18828 16956
rect 18597 16952 18828 16954
rect 18597 16896 18602 16952
rect 18658 16896 18828 16952
rect 18597 16894 18828 16896
rect 18597 16891 18663 16894
rect 18822 16892 18828 16894
rect 18892 16892 18898 16956
rect 7874 16752 8194 16753
rect 7874 16688 7882 16752
rect 7946 16688 7962 16752
rect 8026 16688 8042 16752
rect 8106 16688 8122 16752
rect 8186 16688 8194 16752
rect 7874 16687 8194 16688
rect 14805 16752 15125 16753
rect 14805 16688 14813 16752
rect 14877 16688 14893 16752
rect 14957 16688 14973 16752
rect 15037 16688 15053 16752
rect 15117 16688 15125 16752
rect 14805 16687 15125 16688
rect 17953 16682 18019 16685
rect 22520 16682 23000 16712
rect 17953 16680 23000 16682
rect 17953 16624 17958 16680
rect 18014 16624 23000 16680
rect 17953 16622 23000 16624
rect 17953 16619 18019 16622
rect 22520 16592 23000 16622
rect 4409 16208 4729 16209
rect 4409 16144 4417 16208
rect 4481 16144 4497 16208
rect 4561 16144 4577 16208
rect 4641 16144 4657 16208
rect 4721 16144 4729 16208
rect 4409 16143 4729 16144
rect 11340 16208 11660 16209
rect 11340 16144 11348 16208
rect 11412 16144 11428 16208
rect 11492 16144 11508 16208
rect 11572 16144 11588 16208
rect 11652 16144 11660 16208
rect 11340 16143 11660 16144
rect 18270 16208 18590 16209
rect 18270 16144 18278 16208
rect 18342 16144 18358 16208
rect 18422 16144 18438 16208
rect 18502 16144 18518 16208
rect 18582 16144 18590 16208
rect 18270 16143 18590 16144
rect 19149 16138 19215 16141
rect 22520 16138 23000 16168
rect 19149 16136 23000 16138
rect 19149 16080 19154 16136
rect 19210 16080 23000 16136
rect 19149 16078 23000 16080
rect 19149 16075 19215 16078
rect 22520 16048 23000 16078
rect 19241 15730 19307 15733
rect 22520 15730 23000 15760
rect 19241 15728 23000 15730
rect 19241 15672 19246 15728
rect 19302 15672 23000 15728
rect 19241 15670 23000 15672
rect 19241 15667 19307 15670
rect 7874 15664 8194 15665
rect 7874 15600 7882 15664
rect 7946 15600 7962 15664
rect 8026 15600 8042 15664
rect 8106 15600 8122 15664
rect 8186 15600 8194 15664
rect 7874 15599 8194 15600
rect 14805 15664 15125 15665
rect 14805 15600 14813 15664
rect 14877 15600 14893 15664
rect 14957 15600 14973 15664
rect 15037 15600 15053 15664
rect 15117 15600 15125 15664
rect 22520 15640 23000 15670
rect 14805 15599 15125 15600
rect 18689 15186 18755 15189
rect 22520 15186 23000 15216
rect 18689 15184 23000 15186
rect 18689 15128 18694 15184
rect 18750 15128 23000 15184
rect 18689 15126 23000 15128
rect 18689 15123 18755 15126
rect 4409 15120 4729 15121
rect 4409 15056 4417 15120
rect 4481 15056 4497 15120
rect 4561 15056 4577 15120
rect 4641 15056 4657 15120
rect 4721 15056 4729 15120
rect 4409 15055 4729 15056
rect 11340 15120 11660 15121
rect 11340 15056 11348 15120
rect 11412 15056 11428 15120
rect 11492 15056 11508 15120
rect 11572 15056 11588 15120
rect 11652 15056 11660 15120
rect 11340 15055 11660 15056
rect 18270 15120 18590 15121
rect 18270 15056 18278 15120
rect 18342 15056 18358 15120
rect 18422 15056 18438 15120
rect 18502 15056 18518 15120
rect 18582 15056 18590 15120
rect 22520 15096 23000 15126
rect 18270 15055 18590 15056
rect 19425 14914 19491 14917
rect 19701 14914 19767 14917
rect 19425 14912 19767 14914
rect 19425 14856 19430 14912
rect 19486 14856 19706 14912
rect 19762 14856 19767 14912
rect 19425 14854 19767 14856
rect 19425 14851 19491 14854
rect 19701 14851 19767 14854
rect 19333 14778 19399 14781
rect 19977 14778 20043 14781
rect 19333 14776 20043 14778
rect 19333 14720 19338 14776
rect 19394 14720 19982 14776
rect 20038 14720 20043 14776
rect 19333 14718 20043 14720
rect 19333 14715 19399 14718
rect 19977 14715 20043 14718
rect 18597 14642 18663 14645
rect 22520 14642 23000 14672
rect 18597 14640 23000 14642
rect 18597 14584 18602 14640
rect 18658 14584 23000 14640
rect 18597 14582 23000 14584
rect 18597 14579 18663 14582
rect 7874 14576 8194 14577
rect 7874 14512 7882 14576
rect 7946 14512 7962 14576
rect 8026 14512 8042 14576
rect 8106 14512 8122 14576
rect 8186 14512 8194 14576
rect 7874 14511 8194 14512
rect 14805 14576 15125 14577
rect 14805 14512 14813 14576
rect 14877 14512 14893 14576
rect 14957 14512 14973 14576
rect 15037 14512 15053 14576
rect 15117 14512 15125 14576
rect 22520 14552 23000 14582
rect 14805 14511 15125 14512
rect 17953 14234 18019 14237
rect 22520 14234 23000 14264
rect 17953 14232 23000 14234
rect 17953 14176 17958 14232
rect 18014 14176 23000 14232
rect 17953 14174 23000 14176
rect 17953 14171 18019 14174
rect 22520 14144 23000 14174
rect 4409 14032 4729 14033
rect 4409 13968 4417 14032
rect 4481 13968 4497 14032
rect 4561 13968 4577 14032
rect 4641 13968 4657 14032
rect 4721 13968 4729 14032
rect 4409 13967 4729 13968
rect 11340 14032 11660 14033
rect 11340 13968 11348 14032
rect 11412 13968 11428 14032
rect 11492 13968 11508 14032
rect 11572 13968 11588 14032
rect 11652 13968 11660 14032
rect 11340 13967 11660 13968
rect 18270 14032 18590 14033
rect 18270 13968 18278 14032
rect 18342 13968 18358 14032
rect 18422 13968 18438 14032
rect 18502 13968 18518 14032
rect 18582 13968 18590 14032
rect 18270 13967 18590 13968
rect 20713 13690 20779 13693
rect 22520 13690 23000 13720
rect 20713 13688 23000 13690
rect 20713 13632 20718 13688
rect 20774 13632 23000 13688
rect 20713 13630 23000 13632
rect 20713 13627 20779 13630
rect 22520 13600 23000 13630
rect 7874 13488 8194 13489
rect 7874 13424 7882 13488
rect 7946 13424 7962 13488
rect 8026 13424 8042 13488
rect 8106 13424 8122 13488
rect 8186 13424 8194 13488
rect 7874 13423 8194 13424
rect 14805 13488 15125 13489
rect 14805 13424 14813 13488
rect 14877 13424 14893 13488
rect 14957 13424 14973 13488
rect 15037 13424 15053 13488
rect 15117 13424 15125 13488
rect 14805 13423 15125 13424
rect 20621 13282 20687 13285
rect 22520 13282 23000 13312
rect 20621 13280 23000 13282
rect 20621 13224 20626 13280
rect 20682 13224 23000 13280
rect 20621 13222 23000 13224
rect 20621 13219 20687 13222
rect 22520 13192 23000 13222
rect 9397 13146 9463 13149
rect 9581 13146 9647 13149
rect 9397 13144 9647 13146
rect 9397 13088 9402 13144
rect 9458 13088 9586 13144
rect 9642 13088 9647 13144
rect 9397 13086 9647 13088
rect 9397 13083 9463 13086
rect 9581 13083 9647 13086
rect 4409 12944 4729 12945
rect 4409 12880 4417 12944
rect 4481 12880 4497 12944
rect 4561 12880 4577 12944
rect 4641 12880 4657 12944
rect 4721 12880 4729 12944
rect 4409 12879 4729 12880
rect 11340 12944 11660 12945
rect 11340 12880 11348 12944
rect 11412 12880 11428 12944
rect 11492 12880 11508 12944
rect 11572 12880 11588 12944
rect 11652 12880 11660 12944
rect 11340 12879 11660 12880
rect 18270 12944 18590 12945
rect 18270 12880 18278 12944
rect 18342 12880 18358 12944
rect 18422 12880 18438 12944
rect 18502 12880 18518 12944
rect 18582 12880 18590 12944
rect 18270 12879 18590 12880
rect 19609 12738 19675 12741
rect 22520 12738 23000 12768
rect 19609 12736 23000 12738
rect 19609 12680 19614 12736
rect 19670 12680 23000 12736
rect 19609 12678 23000 12680
rect 19609 12675 19675 12678
rect 22520 12648 23000 12678
rect 7874 12400 8194 12401
rect 7874 12336 7882 12400
rect 7946 12336 7962 12400
rect 8026 12336 8042 12400
rect 8106 12336 8122 12400
rect 8186 12336 8194 12400
rect 7874 12335 8194 12336
rect 14805 12400 15125 12401
rect 14805 12336 14813 12400
rect 14877 12336 14893 12400
rect 14957 12336 14973 12400
rect 15037 12336 15053 12400
rect 15117 12336 15125 12400
rect 14805 12335 15125 12336
rect 18413 12194 18479 12197
rect 22520 12194 23000 12224
rect 18413 12192 23000 12194
rect 18413 12136 18418 12192
rect 18474 12136 23000 12192
rect 18413 12134 23000 12136
rect 18413 12131 18479 12134
rect 22520 12104 23000 12134
rect 4409 11856 4729 11857
rect 4409 11792 4417 11856
rect 4481 11792 4497 11856
rect 4561 11792 4577 11856
rect 4641 11792 4657 11856
rect 4721 11792 4729 11856
rect 4409 11791 4729 11792
rect 11340 11856 11660 11857
rect 11340 11792 11348 11856
rect 11412 11792 11428 11856
rect 11492 11792 11508 11856
rect 11572 11792 11588 11856
rect 11652 11792 11660 11856
rect 11340 11791 11660 11792
rect 18270 11856 18590 11857
rect 18270 11792 18278 11856
rect 18342 11792 18358 11856
rect 18422 11792 18438 11856
rect 18502 11792 18518 11856
rect 18582 11792 18590 11856
rect 18270 11791 18590 11792
rect 18689 11786 18755 11789
rect 22520 11786 23000 11816
rect 18689 11784 23000 11786
rect 18689 11728 18694 11784
rect 18750 11728 23000 11784
rect 18689 11726 23000 11728
rect 18689 11723 18755 11726
rect 22520 11696 23000 11726
rect 7874 11312 8194 11313
rect 7874 11248 7882 11312
rect 7946 11248 7962 11312
rect 8026 11248 8042 11312
rect 8106 11248 8122 11312
rect 8186 11248 8194 11312
rect 7874 11247 8194 11248
rect 14805 11312 15125 11313
rect 14805 11248 14813 11312
rect 14877 11248 14893 11312
rect 14957 11248 14973 11312
rect 15037 11248 15053 11312
rect 15117 11248 15125 11312
rect 14805 11247 15125 11248
rect 17953 11242 18019 11245
rect 22520 11242 23000 11272
rect 17953 11240 23000 11242
rect 17953 11184 17958 11240
rect 18014 11184 23000 11240
rect 17953 11182 23000 11184
rect 17953 11179 18019 11182
rect 22520 11152 23000 11182
rect 19701 10834 19767 10837
rect 22520 10834 23000 10864
rect 19701 10832 23000 10834
rect 19701 10776 19706 10832
rect 19762 10776 23000 10832
rect 19701 10774 23000 10776
rect 19701 10771 19767 10774
rect 4409 10768 4729 10769
rect 4409 10704 4417 10768
rect 4481 10704 4497 10768
rect 4561 10704 4577 10768
rect 4641 10704 4657 10768
rect 4721 10704 4729 10768
rect 4409 10703 4729 10704
rect 11340 10768 11660 10769
rect 11340 10704 11348 10768
rect 11412 10704 11428 10768
rect 11492 10704 11508 10768
rect 11572 10704 11588 10768
rect 11652 10704 11660 10768
rect 11340 10703 11660 10704
rect 18270 10768 18590 10769
rect 18270 10704 18278 10768
rect 18342 10704 18358 10768
rect 18422 10704 18438 10768
rect 18502 10704 18518 10768
rect 18582 10704 18590 10768
rect 22520 10744 23000 10774
rect 18270 10703 18590 10704
rect 20345 10290 20411 10293
rect 22520 10290 23000 10320
rect 20345 10288 23000 10290
rect 20345 10232 20350 10288
rect 20406 10232 23000 10288
rect 20345 10230 23000 10232
rect 20345 10227 20411 10230
rect 7874 10224 8194 10225
rect 7874 10160 7882 10224
rect 7946 10160 7962 10224
rect 8026 10160 8042 10224
rect 8106 10160 8122 10224
rect 8186 10160 8194 10224
rect 7874 10159 8194 10160
rect 14805 10224 15125 10225
rect 14805 10160 14813 10224
rect 14877 10160 14893 10224
rect 14957 10160 14973 10224
rect 15037 10160 15053 10224
rect 15117 10160 15125 10224
rect 22520 10200 23000 10230
rect 14805 10159 15125 10160
rect 19241 9746 19307 9749
rect 22520 9746 23000 9776
rect 19241 9744 23000 9746
rect 19241 9688 19246 9744
rect 19302 9688 23000 9744
rect 19241 9686 23000 9688
rect 19241 9683 19307 9686
rect 4409 9680 4729 9681
rect 4409 9616 4417 9680
rect 4481 9616 4497 9680
rect 4561 9616 4577 9680
rect 4641 9616 4657 9680
rect 4721 9616 4729 9680
rect 4409 9615 4729 9616
rect 11340 9680 11660 9681
rect 11340 9616 11348 9680
rect 11412 9616 11428 9680
rect 11492 9616 11508 9680
rect 11572 9616 11588 9680
rect 11652 9616 11660 9680
rect 11340 9615 11660 9616
rect 18270 9680 18590 9681
rect 18270 9616 18278 9680
rect 18342 9616 18358 9680
rect 18422 9616 18438 9680
rect 18502 9616 18518 9680
rect 18582 9616 18590 9680
rect 22520 9656 23000 9686
rect 18270 9615 18590 9616
rect 18873 9338 18939 9341
rect 22520 9338 23000 9368
rect 18873 9336 23000 9338
rect 18873 9280 18878 9336
rect 18934 9280 23000 9336
rect 18873 9278 23000 9280
rect 18873 9275 18939 9278
rect 22520 9248 23000 9278
rect 7874 9136 8194 9137
rect 7874 9072 7882 9136
rect 7946 9072 7962 9136
rect 8026 9072 8042 9136
rect 8106 9072 8122 9136
rect 8186 9072 8194 9136
rect 7874 9071 8194 9072
rect 14805 9136 15125 9137
rect 14805 9072 14813 9136
rect 14877 9072 14893 9136
rect 14957 9072 14973 9136
rect 15037 9072 15053 9136
rect 15117 9072 15125 9136
rect 14805 9071 15125 9072
rect 20529 8794 20595 8797
rect 22520 8794 23000 8824
rect 20529 8792 23000 8794
rect 20529 8736 20534 8792
rect 20590 8736 23000 8792
rect 20529 8734 23000 8736
rect 20529 8731 20595 8734
rect 22520 8704 23000 8734
rect 4409 8592 4729 8593
rect 4409 8528 4417 8592
rect 4481 8528 4497 8592
rect 4561 8528 4577 8592
rect 4641 8528 4657 8592
rect 4721 8528 4729 8592
rect 4409 8527 4729 8528
rect 11340 8592 11660 8593
rect 11340 8528 11348 8592
rect 11412 8528 11428 8592
rect 11492 8528 11508 8592
rect 11572 8528 11588 8592
rect 11652 8528 11660 8592
rect 11340 8527 11660 8528
rect 18270 8592 18590 8593
rect 18270 8528 18278 8592
rect 18342 8528 18358 8592
rect 18422 8528 18438 8592
rect 18502 8528 18518 8592
rect 18582 8528 18590 8592
rect 18270 8527 18590 8528
rect 19241 8386 19307 8389
rect 22520 8386 23000 8416
rect 19241 8384 23000 8386
rect 19241 8328 19246 8384
rect 19302 8328 23000 8384
rect 19241 8326 23000 8328
rect 19241 8323 19307 8326
rect 22520 8296 23000 8326
rect 7874 8048 8194 8049
rect 7874 7984 7882 8048
rect 7946 7984 7962 8048
rect 8026 7984 8042 8048
rect 8106 7984 8122 8048
rect 8186 7984 8194 8048
rect 7874 7983 8194 7984
rect 14805 8048 15125 8049
rect 14805 7984 14813 8048
rect 14877 7984 14893 8048
rect 14957 7984 14973 8048
rect 15037 7984 15053 8048
rect 15117 7984 15125 8048
rect 14805 7983 15125 7984
rect 20621 7842 20687 7845
rect 22520 7842 23000 7872
rect 20621 7840 23000 7842
rect 20621 7784 20626 7840
rect 20682 7784 23000 7840
rect 20621 7782 23000 7784
rect 20621 7779 20687 7782
rect 22520 7752 23000 7782
rect 4409 7504 4729 7505
rect 4409 7440 4417 7504
rect 4481 7440 4497 7504
rect 4561 7440 4577 7504
rect 4641 7440 4657 7504
rect 4721 7440 4729 7504
rect 4409 7439 4729 7440
rect 11340 7504 11660 7505
rect 11340 7440 11348 7504
rect 11412 7440 11428 7504
rect 11492 7440 11508 7504
rect 11572 7440 11588 7504
rect 11652 7440 11660 7504
rect 11340 7439 11660 7440
rect 18270 7504 18590 7505
rect 18270 7440 18278 7504
rect 18342 7440 18358 7504
rect 18422 7440 18438 7504
rect 18502 7440 18518 7504
rect 18582 7440 18590 7504
rect 18270 7439 18590 7440
rect 19241 7298 19307 7301
rect 22520 7298 23000 7328
rect 19241 7296 23000 7298
rect 19241 7240 19246 7296
rect 19302 7240 23000 7296
rect 19241 7238 23000 7240
rect 19241 7235 19307 7238
rect 22520 7208 23000 7238
rect 7874 6960 8194 6961
rect 7874 6896 7882 6960
rect 7946 6896 7962 6960
rect 8026 6896 8042 6960
rect 8106 6896 8122 6960
rect 8186 6896 8194 6960
rect 7874 6895 8194 6896
rect 14805 6960 15125 6961
rect 14805 6896 14813 6960
rect 14877 6896 14893 6960
rect 14957 6896 14973 6960
rect 15037 6896 15053 6960
rect 15117 6896 15125 6960
rect 14805 6895 15125 6896
rect 20529 6890 20595 6893
rect 22520 6890 23000 6920
rect 20529 6888 23000 6890
rect 20529 6832 20534 6888
rect 20590 6832 23000 6888
rect 20529 6830 23000 6832
rect 20529 6827 20595 6830
rect 22520 6800 23000 6830
rect 4409 6416 4729 6417
rect 4409 6352 4417 6416
rect 4481 6352 4497 6416
rect 4561 6352 4577 6416
rect 4641 6352 4657 6416
rect 4721 6352 4729 6416
rect 4409 6351 4729 6352
rect 11340 6416 11660 6417
rect 11340 6352 11348 6416
rect 11412 6352 11428 6416
rect 11492 6352 11508 6416
rect 11572 6352 11588 6416
rect 11652 6352 11660 6416
rect 11340 6351 11660 6352
rect 18270 6416 18590 6417
rect 18270 6352 18278 6416
rect 18342 6352 18358 6416
rect 18422 6352 18438 6416
rect 18502 6352 18518 6416
rect 18582 6352 18590 6416
rect 18270 6351 18590 6352
rect 19241 6346 19307 6349
rect 22520 6346 23000 6376
rect 19241 6344 23000 6346
rect 19241 6288 19246 6344
rect 19302 6288 23000 6344
rect 19241 6286 23000 6288
rect 19241 6283 19307 6286
rect 22520 6256 23000 6286
rect 20529 5938 20595 5941
rect 22520 5938 23000 5968
rect 20529 5936 23000 5938
rect 20529 5880 20534 5936
rect 20590 5880 23000 5936
rect 20529 5878 23000 5880
rect 20529 5875 20595 5878
rect 7874 5872 8194 5873
rect 7874 5808 7882 5872
rect 7946 5808 7962 5872
rect 8026 5808 8042 5872
rect 8106 5808 8122 5872
rect 8186 5808 8194 5872
rect 7874 5807 8194 5808
rect 14805 5872 15125 5873
rect 14805 5808 14813 5872
rect 14877 5808 14893 5872
rect 14957 5808 14973 5872
rect 15037 5808 15053 5872
rect 15117 5808 15125 5872
rect 22520 5848 23000 5878
rect 14805 5807 15125 5808
rect 0 5666 480 5696
rect 3693 5666 3759 5669
rect 0 5664 3759 5666
rect 0 5608 3698 5664
rect 3754 5608 3759 5664
rect 0 5606 3759 5608
rect 0 5576 480 5606
rect 3693 5603 3759 5606
rect 18689 5394 18755 5397
rect 22520 5394 23000 5424
rect 18689 5392 23000 5394
rect 18689 5336 18694 5392
rect 18750 5336 23000 5392
rect 18689 5334 23000 5336
rect 18689 5331 18755 5334
rect 4409 5328 4729 5329
rect 4409 5264 4417 5328
rect 4481 5264 4497 5328
rect 4561 5264 4577 5328
rect 4641 5264 4657 5328
rect 4721 5264 4729 5328
rect 4409 5263 4729 5264
rect 11340 5328 11660 5329
rect 11340 5264 11348 5328
rect 11412 5264 11428 5328
rect 11492 5264 11508 5328
rect 11572 5264 11588 5328
rect 11652 5264 11660 5328
rect 11340 5263 11660 5264
rect 18270 5328 18590 5329
rect 18270 5264 18278 5328
rect 18342 5264 18358 5328
rect 18422 5264 18438 5328
rect 18502 5264 18518 5328
rect 18582 5264 18590 5328
rect 22520 5304 23000 5334
rect 18270 5263 18590 5264
rect 20529 4850 20595 4853
rect 22520 4850 23000 4880
rect 20529 4848 23000 4850
rect 20529 4792 20534 4848
rect 20590 4792 23000 4848
rect 20529 4790 23000 4792
rect 20529 4787 20595 4790
rect 7874 4784 8194 4785
rect 7874 4720 7882 4784
rect 7946 4720 7962 4784
rect 8026 4720 8042 4784
rect 8106 4720 8122 4784
rect 8186 4720 8194 4784
rect 7874 4719 8194 4720
rect 14805 4784 15125 4785
rect 14805 4720 14813 4784
rect 14877 4720 14893 4784
rect 14957 4720 14973 4784
rect 15037 4720 15053 4784
rect 15117 4720 15125 4784
rect 22520 4760 23000 4790
rect 14805 4719 15125 4720
rect 17953 4442 18019 4445
rect 22520 4442 23000 4472
rect 17953 4440 23000 4442
rect 17953 4384 17958 4440
rect 18014 4384 23000 4440
rect 17953 4382 23000 4384
rect 17953 4379 18019 4382
rect 22520 4352 23000 4382
rect 4409 4240 4729 4241
rect 4409 4176 4417 4240
rect 4481 4176 4497 4240
rect 4561 4176 4577 4240
rect 4641 4176 4657 4240
rect 4721 4176 4729 4240
rect 4409 4175 4729 4176
rect 11340 4240 11660 4241
rect 11340 4176 11348 4240
rect 11412 4176 11428 4240
rect 11492 4176 11508 4240
rect 11572 4176 11588 4240
rect 11652 4176 11660 4240
rect 11340 4175 11660 4176
rect 18270 4240 18590 4241
rect 18270 4176 18278 4240
rect 18342 4176 18358 4240
rect 18422 4176 18438 4240
rect 18502 4176 18518 4240
rect 18582 4176 18590 4240
rect 18270 4175 18590 4176
rect 17953 3898 18019 3901
rect 22520 3898 23000 3928
rect 17953 3896 23000 3898
rect 17953 3840 17958 3896
rect 18014 3840 23000 3896
rect 17953 3838 23000 3840
rect 17953 3835 18019 3838
rect 22520 3808 23000 3838
rect 7874 3696 8194 3697
rect 7874 3632 7882 3696
rect 7946 3632 7962 3696
rect 8026 3632 8042 3696
rect 8106 3632 8122 3696
rect 8186 3632 8194 3696
rect 7874 3631 8194 3632
rect 14805 3696 15125 3697
rect 14805 3632 14813 3696
rect 14877 3632 14893 3696
rect 14957 3632 14973 3696
rect 15037 3632 15053 3696
rect 15117 3632 15125 3696
rect 14805 3631 15125 3632
rect 18045 3490 18111 3493
rect 22520 3490 23000 3520
rect 18045 3488 23000 3490
rect 18045 3432 18050 3488
rect 18106 3432 23000 3488
rect 18045 3430 23000 3432
rect 18045 3427 18111 3430
rect 22520 3400 23000 3430
rect 4409 3152 4729 3153
rect 4409 3088 4417 3152
rect 4481 3088 4497 3152
rect 4561 3088 4577 3152
rect 4641 3088 4657 3152
rect 4721 3088 4729 3152
rect 4409 3087 4729 3088
rect 11340 3152 11660 3153
rect 11340 3088 11348 3152
rect 11412 3088 11428 3152
rect 11492 3088 11508 3152
rect 11572 3088 11588 3152
rect 11652 3088 11660 3152
rect 11340 3087 11660 3088
rect 18270 3152 18590 3153
rect 18270 3088 18278 3152
rect 18342 3088 18358 3152
rect 18422 3088 18438 3152
rect 18502 3088 18518 3152
rect 18582 3088 18590 3152
rect 18270 3087 18590 3088
rect 20529 2946 20595 2949
rect 22520 2946 23000 2976
rect 20529 2944 23000 2946
rect 20529 2888 20534 2944
rect 20590 2888 23000 2944
rect 20529 2886 23000 2888
rect 20529 2883 20595 2886
rect 22520 2856 23000 2886
rect 7874 2608 8194 2609
rect 7874 2544 7882 2608
rect 7946 2544 7962 2608
rect 8026 2544 8042 2608
rect 8106 2544 8122 2608
rect 8186 2544 8194 2608
rect 7874 2543 8194 2544
rect 14805 2608 15125 2609
rect 14805 2544 14813 2608
rect 14877 2544 14893 2608
rect 14957 2544 14973 2608
rect 15037 2544 15053 2608
rect 15117 2544 15125 2608
rect 14805 2543 15125 2544
rect 19149 2402 19215 2405
rect 22520 2402 23000 2432
rect 19149 2400 23000 2402
rect 19149 2344 19154 2400
rect 19210 2344 23000 2400
rect 19149 2342 23000 2344
rect 19149 2339 19215 2342
rect 22520 2312 23000 2342
rect 4409 2064 4729 2065
rect 4409 2000 4417 2064
rect 4481 2000 4497 2064
rect 4561 2000 4577 2064
rect 4641 2000 4657 2064
rect 4721 2000 4729 2064
rect 4409 1999 4729 2000
rect 11340 2064 11660 2065
rect 11340 2000 11348 2064
rect 11412 2000 11428 2064
rect 11492 2000 11508 2064
rect 11572 2000 11588 2064
rect 11652 2000 11660 2064
rect 11340 1999 11660 2000
rect 18270 2064 18590 2065
rect 18270 2000 18278 2064
rect 18342 2000 18358 2064
rect 18422 2000 18438 2064
rect 18502 2000 18518 2064
rect 18582 2000 18590 2064
rect 18270 1999 18590 2000
rect 19241 1994 19307 1997
rect 22520 1994 23000 2024
rect 19241 1992 23000 1994
rect 19241 1936 19246 1992
rect 19302 1936 23000 1992
rect 19241 1934 23000 1936
rect 19241 1931 19307 1934
rect 22520 1904 23000 1934
rect 18597 1450 18663 1453
rect 22520 1450 23000 1480
rect 18597 1448 23000 1450
rect 18597 1392 18602 1448
rect 18658 1392 23000 1448
rect 18597 1390 23000 1392
rect 18597 1387 18663 1390
rect 22520 1360 23000 1390
rect 19241 1042 19307 1045
rect 22520 1042 23000 1072
rect 19241 1040 23000 1042
rect 19241 984 19246 1040
rect 19302 984 23000 1040
rect 19241 982 23000 984
rect 19241 979 19307 982
rect 22520 952 23000 982
rect 18873 498 18939 501
rect 22520 498 23000 528
rect 18873 496 23000 498
rect 18873 440 18878 496
rect 18934 440 23000 496
rect 18873 438 23000 440
rect 18873 435 18939 438
rect 22520 408 23000 438
rect 18965 90 19031 93
rect 22520 90 23000 120
rect 18965 88 23000 90
rect 18965 32 18970 88
rect 19026 32 23000 88
rect 18965 30 23000 32
rect 18965 27 19031 30
rect 22520 0 23000 30
<< via3 >>
rect 4417 20556 4481 20560
rect 4417 20500 4421 20556
rect 4421 20500 4477 20556
rect 4477 20500 4481 20556
rect 4417 20496 4481 20500
rect 4497 20556 4561 20560
rect 4497 20500 4501 20556
rect 4501 20500 4557 20556
rect 4557 20500 4561 20556
rect 4497 20496 4561 20500
rect 4577 20556 4641 20560
rect 4577 20500 4581 20556
rect 4581 20500 4637 20556
rect 4637 20500 4641 20556
rect 4577 20496 4641 20500
rect 4657 20556 4721 20560
rect 4657 20500 4661 20556
rect 4661 20500 4717 20556
rect 4717 20500 4721 20556
rect 4657 20496 4721 20500
rect 11348 20556 11412 20560
rect 11348 20500 11352 20556
rect 11352 20500 11408 20556
rect 11408 20500 11412 20556
rect 11348 20496 11412 20500
rect 11428 20556 11492 20560
rect 11428 20500 11432 20556
rect 11432 20500 11488 20556
rect 11488 20500 11492 20556
rect 11428 20496 11492 20500
rect 11508 20556 11572 20560
rect 11508 20500 11512 20556
rect 11512 20500 11568 20556
rect 11568 20500 11572 20556
rect 11508 20496 11572 20500
rect 11588 20556 11652 20560
rect 11588 20500 11592 20556
rect 11592 20500 11648 20556
rect 11648 20500 11652 20556
rect 11588 20496 11652 20500
rect 18278 20556 18342 20560
rect 18278 20500 18282 20556
rect 18282 20500 18338 20556
rect 18338 20500 18342 20556
rect 18278 20496 18342 20500
rect 18358 20556 18422 20560
rect 18358 20500 18362 20556
rect 18362 20500 18418 20556
rect 18418 20500 18422 20556
rect 18358 20496 18422 20500
rect 18438 20556 18502 20560
rect 18438 20500 18442 20556
rect 18442 20500 18498 20556
rect 18498 20500 18502 20556
rect 18438 20496 18502 20500
rect 18518 20556 18582 20560
rect 18518 20500 18522 20556
rect 18522 20500 18578 20556
rect 18578 20500 18582 20556
rect 18518 20496 18582 20500
rect 7882 20012 7946 20016
rect 7882 19956 7886 20012
rect 7886 19956 7942 20012
rect 7942 19956 7946 20012
rect 7882 19952 7946 19956
rect 7962 20012 8026 20016
rect 7962 19956 7966 20012
rect 7966 19956 8022 20012
rect 8022 19956 8026 20012
rect 7962 19952 8026 19956
rect 8042 20012 8106 20016
rect 8042 19956 8046 20012
rect 8046 19956 8102 20012
rect 8102 19956 8106 20012
rect 8042 19952 8106 19956
rect 8122 20012 8186 20016
rect 8122 19956 8126 20012
rect 8126 19956 8182 20012
rect 8182 19956 8186 20012
rect 8122 19952 8186 19956
rect 14813 20012 14877 20016
rect 14813 19956 14817 20012
rect 14817 19956 14873 20012
rect 14873 19956 14877 20012
rect 14813 19952 14877 19956
rect 14893 20012 14957 20016
rect 14893 19956 14897 20012
rect 14897 19956 14953 20012
rect 14953 19956 14957 20012
rect 14893 19952 14957 19956
rect 14973 20012 15037 20016
rect 14973 19956 14977 20012
rect 14977 19956 15033 20012
rect 15033 19956 15037 20012
rect 14973 19952 15037 19956
rect 15053 20012 15117 20016
rect 15053 19956 15057 20012
rect 15057 19956 15113 20012
rect 15113 19956 15117 20012
rect 15053 19952 15117 19956
rect 4417 19468 4481 19472
rect 4417 19412 4421 19468
rect 4421 19412 4477 19468
rect 4477 19412 4481 19468
rect 4417 19408 4481 19412
rect 4497 19468 4561 19472
rect 4497 19412 4501 19468
rect 4501 19412 4557 19468
rect 4557 19412 4561 19468
rect 4497 19408 4561 19412
rect 4577 19468 4641 19472
rect 4577 19412 4581 19468
rect 4581 19412 4637 19468
rect 4637 19412 4641 19468
rect 4577 19408 4641 19412
rect 4657 19468 4721 19472
rect 4657 19412 4661 19468
rect 4661 19412 4717 19468
rect 4717 19412 4721 19468
rect 4657 19408 4721 19412
rect 11348 19468 11412 19472
rect 11348 19412 11352 19468
rect 11352 19412 11408 19468
rect 11408 19412 11412 19468
rect 11348 19408 11412 19412
rect 11428 19468 11492 19472
rect 11428 19412 11432 19468
rect 11432 19412 11488 19468
rect 11488 19412 11492 19468
rect 11428 19408 11492 19412
rect 11508 19468 11572 19472
rect 11508 19412 11512 19468
rect 11512 19412 11568 19468
rect 11568 19412 11572 19468
rect 11508 19408 11572 19412
rect 11588 19468 11652 19472
rect 11588 19412 11592 19468
rect 11592 19412 11648 19468
rect 11648 19412 11652 19468
rect 11588 19408 11652 19412
rect 18278 19468 18342 19472
rect 18278 19412 18282 19468
rect 18282 19412 18338 19468
rect 18338 19412 18342 19468
rect 18278 19408 18342 19412
rect 18358 19468 18422 19472
rect 18358 19412 18362 19468
rect 18362 19412 18418 19468
rect 18418 19412 18422 19468
rect 18358 19408 18422 19412
rect 18438 19468 18502 19472
rect 18438 19412 18442 19468
rect 18442 19412 18498 19468
rect 18498 19412 18502 19468
rect 18438 19408 18502 19412
rect 18518 19468 18582 19472
rect 18518 19412 18522 19468
rect 18522 19412 18578 19468
rect 18578 19412 18582 19468
rect 18518 19408 18582 19412
rect 7882 18924 7946 18928
rect 7882 18868 7886 18924
rect 7886 18868 7942 18924
rect 7942 18868 7946 18924
rect 7882 18864 7946 18868
rect 7962 18924 8026 18928
rect 7962 18868 7966 18924
rect 7966 18868 8022 18924
rect 8022 18868 8026 18924
rect 7962 18864 8026 18868
rect 8042 18924 8106 18928
rect 8042 18868 8046 18924
rect 8046 18868 8102 18924
rect 8102 18868 8106 18924
rect 8042 18864 8106 18868
rect 8122 18924 8186 18928
rect 8122 18868 8126 18924
rect 8126 18868 8182 18924
rect 8182 18868 8186 18924
rect 8122 18864 8186 18868
rect 14813 18924 14877 18928
rect 14813 18868 14817 18924
rect 14817 18868 14873 18924
rect 14873 18868 14877 18924
rect 14813 18864 14877 18868
rect 14893 18924 14957 18928
rect 14893 18868 14897 18924
rect 14897 18868 14953 18924
rect 14953 18868 14957 18924
rect 14893 18864 14957 18868
rect 14973 18924 15037 18928
rect 14973 18868 14977 18924
rect 14977 18868 15033 18924
rect 15033 18868 15037 18924
rect 14973 18864 15037 18868
rect 15053 18924 15117 18928
rect 15053 18868 15057 18924
rect 15057 18868 15113 18924
rect 15113 18868 15117 18924
rect 15053 18864 15117 18868
rect 18828 18660 18892 18724
rect 4417 18380 4481 18384
rect 4417 18324 4421 18380
rect 4421 18324 4477 18380
rect 4477 18324 4481 18380
rect 4417 18320 4481 18324
rect 4497 18380 4561 18384
rect 4497 18324 4501 18380
rect 4501 18324 4557 18380
rect 4557 18324 4561 18380
rect 4497 18320 4561 18324
rect 4577 18380 4641 18384
rect 4577 18324 4581 18380
rect 4581 18324 4637 18380
rect 4637 18324 4641 18380
rect 4577 18320 4641 18324
rect 4657 18380 4721 18384
rect 4657 18324 4661 18380
rect 4661 18324 4717 18380
rect 4717 18324 4721 18380
rect 4657 18320 4721 18324
rect 11348 18380 11412 18384
rect 11348 18324 11352 18380
rect 11352 18324 11408 18380
rect 11408 18324 11412 18380
rect 11348 18320 11412 18324
rect 11428 18380 11492 18384
rect 11428 18324 11432 18380
rect 11432 18324 11488 18380
rect 11488 18324 11492 18380
rect 11428 18320 11492 18324
rect 11508 18380 11572 18384
rect 11508 18324 11512 18380
rect 11512 18324 11568 18380
rect 11568 18324 11572 18380
rect 11508 18320 11572 18324
rect 11588 18380 11652 18384
rect 11588 18324 11592 18380
rect 11592 18324 11648 18380
rect 11648 18324 11652 18380
rect 11588 18320 11652 18324
rect 18278 18380 18342 18384
rect 18278 18324 18282 18380
rect 18282 18324 18338 18380
rect 18338 18324 18342 18380
rect 18278 18320 18342 18324
rect 18358 18380 18422 18384
rect 18358 18324 18362 18380
rect 18362 18324 18418 18380
rect 18418 18324 18422 18380
rect 18358 18320 18422 18324
rect 18438 18380 18502 18384
rect 18438 18324 18442 18380
rect 18442 18324 18498 18380
rect 18498 18324 18502 18380
rect 18438 18320 18502 18324
rect 18518 18380 18582 18384
rect 18518 18324 18522 18380
rect 18522 18324 18578 18380
rect 18578 18324 18582 18380
rect 18518 18320 18582 18324
rect 7882 17836 7946 17840
rect 7882 17780 7886 17836
rect 7886 17780 7942 17836
rect 7942 17780 7946 17836
rect 7882 17776 7946 17780
rect 7962 17836 8026 17840
rect 7962 17780 7966 17836
rect 7966 17780 8022 17836
rect 8022 17780 8026 17836
rect 7962 17776 8026 17780
rect 8042 17836 8106 17840
rect 8042 17780 8046 17836
rect 8046 17780 8102 17836
rect 8102 17780 8106 17836
rect 8042 17776 8106 17780
rect 8122 17836 8186 17840
rect 8122 17780 8126 17836
rect 8126 17780 8182 17836
rect 8182 17780 8186 17836
rect 8122 17776 8186 17780
rect 14813 17836 14877 17840
rect 14813 17780 14817 17836
rect 14817 17780 14873 17836
rect 14873 17780 14877 17836
rect 14813 17776 14877 17780
rect 14893 17836 14957 17840
rect 14893 17780 14897 17836
rect 14897 17780 14953 17836
rect 14953 17780 14957 17836
rect 14893 17776 14957 17780
rect 14973 17836 15037 17840
rect 14973 17780 14977 17836
rect 14977 17780 15033 17836
rect 15033 17780 15037 17836
rect 14973 17776 15037 17780
rect 15053 17836 15117 17840
rect 15053 17780 15057 17836
rect 15057 17780 15113 17836
rect 15113 17780 15117 17836
rect 15053 17776 15117 17780
rect 4417 17292 4481 17296
rect 4417 17236 4421 17292
rect 4421 17236 4477 17292
rect 4477 17236 4481 17292
rect 4417 17232 4481 17236
rect 4497 17292 4561 17296
rect 4497 17236 4501 17292
rect 4501 17236 4557 17292
rect 4557 17236 4561 17292
rect 4497 17232 4561 17236
rect 4577 17292 4641 17296
rect 4577 17236 4581 17292
rect 4581 17236 4637 17292
rect 4637 17236 4641 17292
rect 4577 17232 4641 17236
rect 4657 17292 4721 17296
rect 4657 17236 4661 17292
rect 4661 17236 4717 17292
rect 4717 17236 4721 17292
rect 4657 17232 4721 17236
rect 11348 17292 11412 17296
rect 11348 17236 11352 17292
rect 11352 17236 11408 17292
rect 11408 17236 11412 17292
rect 11348 17232 11412 17236
rect 11428 17292 11492 17296
rect 11428 17236 11432 17292
rect 11432 17236 11488 17292
rect 11488 17236 11492 17292
rect 11428 17232 11492 17236
rect 11508 17292 11572 17296
rect 11508 17236 11512 17292
rect 11512 17236 11568 17292
rect 11568 17236 11572 17292
rect 11508 17232 11572 17236
rect 11588 17292 11652 17296
rect 11588 17236 11592 17292
rect 11592 17236 11648 17292
rect 11648 17236 11652 17292
rect 11588 17232 11652 17236
rect 18278 17292 18342 17296
rect 18278 17236 18282 17292
rect 18282 17236 18338 17292
rect 18338 17236 18342 17292
rect 18278 17232 18342 17236
rect 18358 17292 18422 17296
rect 18358 17236 18362 17292
rect 18362 17236 18418 17292
rect 18418 17236 18422 17292
rect 18358 17232 18422 17236
rect 18438 17292 18502 17296
rect 18438 17236 18442 17292
rect 18442 17236 18498 17292
rect 18498 17236 18502 17292
rect 18438 17232 18502 17236
rect 18518 17292 18582 17296
rect 18518 17236 18522 17292
rect 18522 17236 18578 17292
rect 18578 17236 18582 17292
rect 18518 17232 18582 17236
rect 18828 16892 18892 16956
rect 7882 16748 7946 16752
rect 7882 16692 7886 16748
rect 7886 16692 7942 16748
rect 7942 16692 7946 16748
rect 7882 16688 7946 16692
rect 7962 16748 8026 16752
rect 7962 16692 7966 16748
rect 7966 16692 8022 16748
rect 8022 16692 8026 16748
rect 7962 16688 8026 16692
rect 8042 16748 8106 16752
rect 8042 16692 8046 16748
rect 8046 16692 8102 16748
rect 8102 16692 8106 16748
rect 8042 16688 8106 16692
rect 8122 16748 8186 16752
rect 8122 16692 8126 16748
rect 8126 16692 8182 16748
rect 8182 16692 8186 16748
rect 8122 16688 8186 16692
rect 14813 16748 14877 16752
rect 14813 16692 14817 16748
rect 14817 16692 14873 16748
rect 14873 16692 14877 16748
rect 14813 16688 14877 16692
rect 14893 16748 14957 16752
rect 14893 16692 14897 16748
rect 14897 16692 14953 16748
rect 14953 16692 14957 16748
rect 14893 16688 14957 16692
rect 14973 16748 15037 16752
rect 14973 16692 14977 16748
rect 14977 16692 15033 16748
rect 15033 16692 15037 16748
rect 14973 16688 15037 16692
rect 15053 16748 15117 16752
rect 15053 16692 15057 16748
rect 15057 16692 15113 16748
rect 15113 16692 15117 16748
rect 15053 16688 15117 16692
rect 4417 16204 4481 16208
rect 4417 16148 4421 16204
rect 4421 16148 4477 16204
rect 4477 16148 4481 16204
rect 4417 16144 4481 16148
rect 4497 16204 4561 16208
rect 4497 16148 4501 16204
rect 4501 16148 4557 16204
rect 4557 16148 4561 16204
rect 4497 16144 4561 16148
rect 4577 16204 4641 16208
rect 4577 16148 4581 16204
rect 4581 16148 4637 16204
rect 4637 16148 4641 16204
rect 4577 16144 4641 16148
rect 4657 16204 4721 16208
rect 4657 16148 4661 16204
rect 4661 16148 4717 16204
rect 4717 16148 4721 16204
rect 4657 16144 4721 16148
rect 11348 16204 11412 16208
rect 11348 16148 11352 16204
rect 11352 16148 11408 16204
rect 11408 16148 11412 16204
rect 11348 16144 11412 16148
rect 11428 16204 11492 16208
rect 11428 16148 11432 16204
rect 11432 16148 11488 16204
rect 11488 16148 11492 16204
rect 11428 16144 11492 16148
rect 11508 16204 11572 16208
rect 11508 16148 11512 16204
rect 11512 16148 11568 16204
rect 11568 16148 11572 16204
rect 11508 16144 11572 16148
rect 11588 16204 11652 16208
rect 11588 16148 11592 16204
rect 11592 16148 11648 16204
rect 11648 16148 11652 16204
rect 11588 16144 11652 16148
rect 18278 16204 18342 16208
rect 18278 16148 18282 16204
rect 18282 16148 18338 16204
rect 18338 16148 18342 16204
rect 18278 16144 18342 16148
rect 18358 16204 18422 16208
rect 18358 16148 18362 16204
rect 18362 16148 18418 16204
rect 18418 16148 18422 16204
rect 18358 16144 18422 16148
rect 18438 16204 18502 16208
rect 18438 16148 18442 16204
rect 18442 16148 18498 16204
rect 18498 16148 18502 16204
rect 18438 16144 18502 16148
rect 18518 16204 18582 16208
rect 18518 16148 18522 16204
rect 18522 16148 18578 16204
rect 18578 16148 18582 16204
rect 18518 16144 18582 16148
rect 7882 15660 7946 15664
rect 7882 15604 7886 15660
rect 7886 15604 7942 15660
rect 7942 15604 7946 15660
rect 7882 15600 7946 15604
rect 7962 15660 8026 15664
rect 7962 15604 7966 15660
rect 7966 15604 8022 15660
rect 8022 15604 8026 15660
rect 7962 15600 8026 15604
rect 8042 15660 8106 15664
rect 8042 15604 8046 15660
rect 8046 15604 8102 15660
rect 8102 15604 8106 15660
rect 8042 15600 8106 15604
rect 8122 15660 8186 15664
rect 8122 15604 8126 15660
rect 8126 15604 8182 15660
rect 8182 15604 8186 15660
rect 8122 15600 8186 15604
rect 14813 15660 14877 15664
rect 14813 15604 14817 15660
rect 14817 15604 14873 15660
rect 14873 15604 14877 15660
rect 14813 15600 14877 15604
rect 14893 15660 14957 15664
rect 14893 15604 14897 15660
rect 14897 15604 14953 15660
rect 14953 15604 14957 15660
rect 14893 15600 14957 15604
rect 14973 15660 15037 15664
rect 14973 15604 14977 15660
rect 14977 15604 15033 15660
rect 15033 15604 15037 15660
rect 14973 15600 15037 15604
rect 15053 15660 15117 15664
rect 15053 15604 15057 15660
rect 15057 15604 15113 15660
rect 15113 15604 15117 15660
rect 15053 15600 15117 15604
rect 4417 15116 4481 15120
rect 4417 15060 4421 15116
rect 4421 15060 4477 15116
rect 4477 15060 4481 15116
rect 4417 15056 4481 15060
rect 4497 15116 4561 15120
rect 4497 15060 4501 15116
rect 4501 15060 4557 15116
rect 4557 15060 4561 15116
rect 4497 15056 4561 15060
rect 4577 15116 4641 15120
rect 4577 15060 4581 15116
rect 4581 15060 4637 15116
rect 4637 15060 4641 15116
rect 4577 15056 4641 15060
rect 4657 15116 4721 15120
rect 4657 15060 4661 15116
rect 4661 15060 4717 15116
rect 4717 15060 4721 15116
rect 4657 15056 4721 15060
rect 11348 15116 11412 15120
rect 11348 15060 11352 15116
rect 11352 15060 11408 15116
rect 11408 15060 11412 15116
rect 11348 15056 11412 15060
rect 11428 15116 11492 15120
rect 11428 15060 11432 15116
rect 11432 15060 11488 15116
rect 11488 15060 11492 15116
rect 11428 15056 11492 15060
rect 11508 15116 11572 15120
rect 11508 15060 11512 15116
rect 11512 15060 11568 15116
rect 11568 15060 11572 15116
rect 11508 15056 11572 15060
rect 11588 15116 11652 15120
rect 11588 15060 11592 15116
rect 11592 15060 11648 15116
rect 11648 15060 11652 15116
rect 11588 15056 11652 15060
rect 18278 15116 18342 15120
rect 18278 15060 18282 15116
rect 18282 15060 18338 15116
rect 18338 15060 18342 15116
rect 18278 15056 18342 15060
rect 18358 15116 18422 15120
rect 18358 15060 18362 15116
rect 18362 15060 18418 15116
rect 18418 15060 18422 15116
rect 18358 15056 18422 15060
rect 18438 15116 18502 15120
rect 18438 15060 18442 15116
rect 18442 15060 18498 15116
rect 18498 15060 18502 15116
rect 18438 15056 18502 15060
rect 18518 15116 18582 15120
rect 18518 15060 18522 15116
rect 18522 15060 18578 15116
rect 18578 15060 18582 15116
rect 18518 15056 18582 15060
rect 7882 14572 7946 14576
rect 7882 14516 7886 14572
rect 7886 14516 7942 14572
rect 7942 14516 7946 14572
rect 7882 14512 7946 14516
rect 7962 14572 8026 14576
rect 7962 14516 7966 14572
rect 7966 14516 8022 14572
rect 8022 14516 8026 14572
rect 7962 14512 8026 14516
rect 8042 14572 8106 14576
rect 8042 14516 8046 14572
rect 8046 14516 8102 14572
rect 8102 14516 8106 14572
rect 8042 14512 8106 14516
rect 8122 14572 8186 14576
rect 8122 14516 8126 14572
rect 8126 14516 8182 14572
rect 8182 14516 8186 14572
rect 8122 14512 8186 14516
rect 14813 14572 14877 14576
rect 14813 14516 14817 14572
rect 14817 14516 14873 14572
rect 14873 14516 14877 14572
rect 14813 14512 14877 14516
rect 14893 14572 14957 14576
rect 14893 14516 14897 14572
rect 14897 14516 14953 14572
rect 14953 14516 14957 14572
rect 14893 14512 14957 14516
rect 14973 14572 15037 14576
rect 14973 14516 14977 14572
rect 14977 14516 15033 14572
rect 15033 14516 15037 14572
rect 14973 14512 15037 14516
rect 15053 14572 15117 14576
rect 15053 14516 15057 14572
rect 15057 14516 15113 14572
rect 15113 14516 15117 14572
rect 15053 14512 15117 14516
rect 4417 14028 4481 14032
rect 4417 13972 4421 14028
rect 4421 13972 4477 14028
rect 4477 13972 4481 14028
rect 4417 13968 4481 13972
rect 4497 14028 4561 14032
rect 4497 13972 4501 14028
rect 4501 13972 4557 14028
rect 4557 13972 4561 14028
rect 4497 13968 4561 13972
rect 4577 14028 4641 14032
rect 4577 13972 4581 14028
rect 4581 13972 4637 14028
rect 4637 13972 4641 14028
rect 4577 13968 4641 13972
rect 4657 14028 4721 14032
rect 4657 13972 4661 14028
rect 4661 13972 4717 14028
rect 4717 13972 4721 14028
rect 4657 13968 4721 13972
rect 11348 14028 11412 14032
rect 11348 13972 11352 14028
rect 11352 13972 11408 14028
rect 11408 13972 11412 14028
rect 11348 13968 11412 13972
rect 11428 14028 11492 14032
rect 11428 13972 11432 14028
rect 11432 13972 11488 14028
rect 11488 13972 11492 14028
rect 11428 13968 11492 13972
rect 11508 14028 11572 14032
rect 11508 13972 11512 14028
rect 11512 13972 11568 14028
rect 11568 13972 11572 14028
rect 11508 13968 11572 13972
rect 11588 14028 11652 14032
rect 11588 13972 11592 14028
rect 11592 13972 11648 14028
rect 11648 13972 11652 14028
rect 11588 13968 11652 13972
rect 18278 14028 18342 14032
rect 18278 13972 18282 14028
rect 18282 13972 18338 14028
rect 18338 13972 18342 14028
rect 18278 13968 18342 13972
rect 18358 14028 18422 14032
rect 18358 13972 18362 14028
rect 18362 13972 18418 14028
rect 18418 13972 18422 14028
rect 18358 13968 18422 13972
rect 18438 14028 18502 14032
rect 18438 13972 18442 14028
rect 18442 13972 18498 14028
rect 18498 13972 18502 14028
rect 18438 13968 18502 13972
rect 18518 14028 18582 14032
rect 18518 13972 18522 14028
rect 18522 13972 18578 14028
rect 18578 13972 18582 14028
rect 18518 13968 18582 13972
rect 7882 13484 7946 13488
rect 7882 13428 7886 13484
rect 7886 13428 7942 13484
rect 7942 13428 7946 13484
rect 7882 13424 7946 13428
rect 7962 13484 8026 13488
rect 7962 13428 7966 13484
rect 7966 13428 8022 13484
rect 8022 13428 8026 13484
rect 7962 13424 8026 13428
rect 8042 13484 8106 13488
rect 8042 13428 8046 13484
rect 8046 13428 8102 13484
rect 8102 13428 8106 13484
rect 8042 13424 8106 13428
rect 8122 13484 8186 13488
rect 8122 13428 8126 13484
rect 8126 13428 8182 13484
rect 8182 13428 8186 13484
rect 8122 13424 8186 13428
rect 14813 13484 14877 13488
rect 14813 13428 14817 13484
rect 14817 13428 14873 13484
rect 14873 13428 14877 13484
rect 14813 13424 14877 13428
rect 14893 13484 14957 13488
rect 14893 13428 14897 13484
rect 14897 13428 14953 13484
rect 14953 13428 14957 13484
rect 14893 13424 14957 13428
rect 14973 13484 15037 13488
rect 14973 13428 14977 13484
rect 14977 13428 15033 13484
rect 15033 13428 15037 13484
rect 14973 13424 15037 13428
rect 15053 13484 15117 13488
rect 15053 13428 15057 13484
rect 15057 13428 15113 13484
rect 15113 13428 15117 13484
rect 15053 13424 15117 13428
rect 4417 12940 4481 12944
rect 4417 12884 4421 12940
rect 4421 12884 4477 12940
rect 4477 12884 4481 12940
rect 4417 12880 4481 12884
rect 4497 12940 4561 12944
rect 4497 12884 4501 12940
rect 4501 12884 4557 12940
rect 4557 12884 4561 12940
rect 4497 12880 4561 12884
rect 4577 12940 4641 12944
rect 4577 12884 4581 12940
rect 4581 12884 4637 12940
rect 4637 12884 4641 12940
rect 4577 12880 4641 12884
rect 4657 12940 4721 12944
rect 4657 12884 4661 12940
rect 4661 12884 4717 12940
rect 4717 12884 4721 12940
rect 4657 12880 4721 12884
rect 11348 12940 11412 12944
rect 11348 12884 11352 12940
rect 11352 12884 11408 12940
rect 11408 12884 11412 12940
rect 11348 12880 11412 12884
rect 11428 12940 11492 12944
rect 11428 12884 11432 12940
rect 11432 12884 11488 12940
rect 11488 12884 11492 12940
rect 11428 12880 11492 12884
rect 11508 12940 11572 12944
rect 11508 12884 11512 12940
rect 11512 12884 11568 12940
rect 11568 12884 11572 12940
rect 11508 12880 11572 12884
rect 11588 12940 11652 12944
rect 11588 12884 11592 12940
rect 11592 12884 11648 12940
rect 11648 12884 11652 12940
rect 11588 12880 11652 12884
rect 18278 12940 18342 12944
rect 18278 12884 18282 12940
rect 18282 12884 18338 12940
rect 18338 12884 18342 12940
rect 18278 12880 18342 12884
rect 18358 12940 18422 12944
rect 18358 12884 18362 12940
rect 18362 12884 18418 12940
rect 18418 12884 18422 12940
rect 18358 12880 18422 12884
rect 18438 12940 18502 12944
rect 18438 12884 18442 12940
rect 18442 12884 18498 12940
rect 18498 12884 18502 12940
rect 18438 12880 18502 12884
rect 18518 12940 18582 12944
rect 18518 12884 18522 12940
rect 18522 12884 18578 12940
rect 18578 12884 18582 12940
rect 18518 12880 18582 12884
rect 7882 12396 7946 12400
rect 7882 12340 7886 12396
rect 7886 12340 7942 12396
rect 7942 12340 7946 12396
rect 7882 12336 7946 12340
rect 7962 12396 8026 12400
rect 7962 12340 7966 12396
rect 7966 12340 8022 12396
rect 8022 12340 8026 12396
rect 7962 12336 8026 12340
rect 8042 12396 8106 12400
rect 8042 12340 8046 12396
rect 8046 12340 8102 12396
rect 8102 12340 8106 12396
rect 8042 12336 8106 12340
rect 8122 12396 8186 12400
rect 8122 12340 8126 12396
rect 8126 12340 8182 12396
rect 8182 12340 8186 12396
rect 8122 12336 8186 12340
rect 14813 12396 14877 12400
rect 14813 12340 14817 12396
rect 14817 12340 14873 12396
rect 14873 12340 14877 12396
rect 14813 12336 14877 12340
rect 14893 12396 14957 12400
rect 14893 12340 14897 12396
rect 14897 12340 14953 12396
rect 14953 12340 14957 12396
rect 14893 12336 14957 12340
rect 14973 12396 15037 12400
rect 14973 12340 14977 12396
rect 14977 12340 15033 12396
rect 15033 12340 15037 12396
rect 14973 12336 15037 12340
rect 15053 12396 15117 12400
rect 15053 12340 15057 12396
rect 15057 12340 15113 12396
rect 15113 12340 15117 12396
rect 15053 12336 15117 12340
rect 4417 11852 4481 11856
rect 4417 11796 4421 11852
rect 4421 11796 4477 11852
rect 4477 11796 4481 11852
rect 4417 11792 4481 11796
rect 4497 11852 4561 11856
rect 4497 11796 4501 11852
rect 4501 11796 4557 11852
rect 4557 11796 4561 11852
rect 4497 11792 4561 11796
rect 4577 11852 4641 11856
rect 4577 11796 4581 11852
rect 4581 11796 4637 11852
rect 4637 11796 4641 11852
rect 4577 11792 4641 11796
rect 4657 11852 4721 11856
rect 4657 11796 4661 11852
rect 4661 11796 4717 11852
rect 4717 11796 4721 11852
rect 4657 11792 4721 11796
rect 11348 11852 11412 11856
rect 11348 11796 11352 11852
rect 11352 11796 11408 11852
rect 11408 11796 11412 11852
rect 11348 11792 11412 11796
rect 11428 11852 11492 11856
rect 11428 11796 11432 11852
rect 11432 11796 11488 11852
rect 11488 11796 11492 11852
rect 11428 11792 11492 11796
rect 11508 11852 11572 11856
rect 11508 11796 11512 11852
rect 11512 11796 11568 11852
rect 11568 11796 11572 11852
rect 11508 11792 11572 11796
rect 11588 11852 11652 11856
rect 11588 11796 11592 11852
rect 11592 11796 11648 11852
rect 11648 11796 11652 11852
rect 11588 11792 11652 11796
rect 18278 11852 18342 11856
rect 18278 11796 18282 11852
rect 18282 11796 18338 11852
rect 18338 11796 18342 11852
rect 18278 11792 18342 11796
rect 18358 11852 18422 11856
rect 18358 11796 18362 11852
rect 18362 11796 18418 11852
rect 18418 11796 18422 11852
rect 18358 11792 18422 11796
rect 18438 11852 18502 11856
rect 18438 11796 18442 11852
rect 18442 11796 18498 11852
rect 18498 11796 18502 11852
rect 18438 11792 18502 11796
rect 18518 11852 18582 11856
rect 18518 11796 18522 11852
rect 18522 11796 18578 11852
rect 18578 11796 18582 11852
rect 18518 11792 18582 11796
rect 7882 11308 7946 11312
rect 7882 11252 7886 11308
rect 7886 11252 7942 11308
rect 7942 11252 7946 11308
rect 7882 11248 7946 11252
rect 7962 11308 8026 11312
rect 7962 11252 7966 11308
rect 7966 11252 8022 11308
rect 8022 11252 8026 11308
rect 7962 11248 8026 11252
rect 8042 11308 8106 11312
rect 8042 11252 8046 11308
rect 8046 11252 8102 11308
rect 8102 11252 8106 11308
rect 8042 11248 8106 11252
rect 8122 11308 8186 11312
rect 8122 11252 8126 11308
rect 8126 11252 8182 11308
rect 8182 11252 8186 11308
rect 8122 11248 8186 11252
rect 14813 11308 14877 11312
rect 14813 11252 14817 11308
rect 14817 11252 14873 11308
rect 14873 11252 14877 11308
rect 14813 11248 14877 11252
rect 14893 11308 14957 11312
rect 14893 11252 14897 11308
rect 14897 11252 14953 11308
rect 14953 11252 14957 11308
rect 14893 11248 14957 11252
rect 14973 11308 15037 11312
rect 14973 11252 14977 11308
rect 14977 11252 15033 11308
rect 15033 11252 15037 11308
rect 14973 11248 15037 11252
rect 15053 11308 15117 11312
rect 15053 11252 15057 11308
rect 15057 11252 15113 11308
rect 15113 11252 15117 11308
rect 15053 11248 15117 11252
rect 4417 10764 4481 10768
rect 4417 10708 4421 10764
rect 4421 10708 4477 10764
rect 4477 10708 4481 10764
rect 4417 10704 4481 10708
rect 4497 10764 4561 10768
rect 4497 10708 4501 10764
rect 4501 10708 4557 10764
rect 4557 10708 4561 10764
rect 4497 10704 4561 10708
rect 4577 10764 4641 10768
rect 4577 10708 4581 10764
rect 4581 10708 4637 10764
rect 4637 10708 4641 10764
rect 4577 10704 4641 10708
rect 4657 10764 4721 10768
rect 4657 10708 4661 10764
rect 4661 10708 4717 10764
rect 4717 10708 4721 10764
rect 4657 10704 4721 10708
rect 11348 10764 11412 10768
rect 11348 10708 11352 10764
rect 11352 10708 11408 10764
rect 11408 10708 11412 10764
rect 11348 10704 11412 10708
rect 11428 10764 11492 10768
rect 11428 10708 11432 10764
rect 11432 10708 11488 10764
rect 11488 10708 11492 10764
rect 11428 10704 11492 10708
rect 11508 10764 11572 10768
rect 11508 10708 11512 10764
rect 11512 10708 11568 10764
rect 11568 10708 11572 10764
rect 11508 10704 11572 10708
rect 11588 10764 11652 10768
rect 11588 10708 11592 10764
rect 11592 10708 11648 10764
rect 11648 10708 11652 10764
rect 11588 10704 11652 10708
rect 18278 10764 18342 10768
rect 18278 10708 18282 10764
rect 18282 10708 18338 10764
rect 18338 10708 18342 10764
rect 18278 10704 18342 10708
rect 18358 10764 18422 10768
rect 18358 10708 18362 10764
rect 18362 10708 18418 10764
rect 18418 10708 18422 10764
rect 18358 10704 18422 10708
rect 18438 10764 18502 10768
rect 18438 10708 18442 10764
rect 18442 10708 18498 10764
rect 18498 10708 18502 10764
rect 18438 10704 18502 10708
rect 18518 10764 18582 10768
rect 18518 10708 18522 10764
rect 18522 10708 18578 10764
rect 18578 10708 18582 10764
rect 18518 10704 18582 10708
rect 7882 10220 7946 10224
rect 7882 10164 7886 10220
rect 7886 10164 7942 10220
rect 7942 10164 7946 10220
rect 7882 10160 7946 10164
rect 7962 10220 8026 10224
rect 7962 10164 7966 10220
rect 7966 10164 8022 10220
rect 8022 10164 8026 10220
rect 7962 10160 8026 10164
rect 8042 10220 8106 10224
rect 8042 10164 8046 10220
rect 8046 10164 8102 10220
rect 8102 10164 8106 10220
rect 8042 10160 8106 10164
rect 8122 10220 8186 10224
rect 8122 10164 8126 10220
rect 8126 10164 8182 10220
rect 8182 10164 8186 10220
rect 8122 10160 8186 10164
rect 14813 10220 14877 10224
rect 14813 10164 14817 10220
rect 14817 10164 14873 10220
rect 14873 10164 14877 10220
rect 14813 10160 14877 10164
rect 14893 10220 14957 10224
rect 14893 10164 14897 10220
rect 14897 10164 14953 10220
rect 14953 10164 14957 10220
rect 14893 10160 14957 10164
rect 14973 10220 15037 10224
rect 14973 10164 14977 10220
rect 14977 10164 15033 10220
rect 15033 10164 15037 10220
rect 14973 10160 15037 10164
rect 15053 10220 15117 10224
rect 15053 10164 15057 10220
rect 15057 10164 15113 10220
rect 15113 10164 15117 10220
rect 15053 10160 15117 10164
rect 4417 9676 4481 9680
rect 4417 9620 4421 9676
rect 4421 9620 4477 9676
rect 4477 9620 4481 9676
rect 4417 9616 4481 9620
rect 4497 9676 4561 9680
rect 4497 9620 4501 9676
rect 4501 9620 4557 9676
rect 4557 9620 4561 9676
rect 4497 9616 4561 9620
rect 4577 9676 4641 9680
rect 4577 9620 4581 9676
rect 4581 9620 4637 9676
rect 4637 9620 4641 9676
rect 4577 9616 4641 9620
rect 4657 9676 4721 9680
rect 4657 9620 4661 9676
rect 4661 9620 4717 9676
rect 4717 9620 4721 9676
rect 4657 9616 4721 9620
rect 11348 9676 11412 9680
rect 11348 9620 11352 9676
rect 11352 9620 11408 9676
rect 11408 9620 11412 9676
rect 11348 9616 11412 9620
rect 11428 9676 11492 9680
rect 11428 9620 11432 9676
rect 11432 9620 11488 9676
rect 11488 9620 11492 9676
rect 11428 9616 11492 9620
rect 11508 9676 11572 9680
rect 11508 9620 11512 9676
rect 11512 9620 11568 9676
rect 11568 9620 11572 9676
rect 11508 9616 11572 9620
rect 11588 9676 11652 9680
rect 11588 9620 11592 9676
rect 11592 9620 11648 9676
rect 11648 9620 11652 9676
rect 11588 9616 11652 9620
rect 18278 9676 18342 9680
rect 18278 9620 18282 9676
rect 18282 9620 18338 9676
rect 18338 9620 18342 9676
rect 18278 9616 18342 9620
rect 18358 9676 18422 9680
rect 18358 9620 18362 9676
rect 18362 9620 18418 9676
rect 18418 9620 18422 9676
rect 18358 9616 18422 9620
rect 18438 9676 18502 9680
rect 18438 9620 18442 9676
rect 18442 9620 18498 9676
rect 18498 9620 18502 9676
rect 18438 9616 18502 9620
rect 18518 9676 18582 9680
rect 18518 9620 18522 9676
rect 18522 9620 18578 9676
rect 18578 9620 18582 9676
rect 18518 9616 18582 9620
rect 7882 9132 7946 9136
rect 7882 9076 7886 9132
rect 7886 9076 7942 9132
rect 7942 9076 7946 9132
rect 7882 9072 7946 9076
rect 7962 9132 8026 9136
rect 7962 9076 7966 9132
rect 7966 9076 8022 9132
rect 8022 9076 8026 9132
rect 7962 9072 8026 9076
rect 8042 9132 8106 9136
rect 8042 9076 8046 9132
rect 8046 9076 8102 9132
rect 8102 9076 8106 9132
rect 8042 9072 8106 9076
rect 8122 9132 8186 9136
rect 8122 9076 8126 9132
rect 8126 9076 8182 9132
rect 8182 9076 8186 9132
rect 8122 9072 8186 9076
rect 14813 9132 14877 9136
rect 14813 9076 14817 9132
rect 14817 9076 14873 9132
rect 14873 9076 14877 9132
rect 14813 9072 14877 9076
rect 14893 9132 14957 9136
rect 14893 9076 14897 9132
rect 14897 9076 14953 9132
rect 14953 9076 14957 9132
rect 14893 9072 14957 9076
rect 14973 9132 15037 9136
rect 14973 9076 14977 9132
rect 14977 9076 15033 9132
rect 15033 9076 15037 9132
rect 14973 9072 15037 9076
rect 15053 9132 15117 9136
rect 15053 9076 15057 9132
rect 15057 9076 15113 9132
rect 15113 9076 15117 9132
rect 15053 9072 15117 9076
rect 4417 8588 4481 8592
rect 4417 8532 4421 8588
rect 4421 8532 4477 8588
rect 4477 8532 4481 8588
rect 4417 8528 4481 8532
rect 4497 8588 4561 8592
rect 4497 8532 4501 8588
rect 4501 8532 4557 8588
rect 4557 8532 4561 8588
rect 4497 8528 4561 8532
rect 4577 8588 4641 8592
rect 4577 8532 4581 8588
rect 4581 8532 4637 8588
rect 4637 8532 4641 8588
rect 4577 8528 4641 8532
rect 4657 8588 4721 8592
rect 4657 8532 4661 8588
rect 4661 8532 4717 8588
rect 4717 8532 4721 8588
rect 4657 8528 4721 8532
rect 11348 8588 11412 8592
rect 11348 8532 11352 8588
rect 11352 8532 11408 8588
rect 11408 8532 11412 8588
rect 11348 8528 11412 8532
rect 11428 8588 11492 8592
rect 11428 8532 11432 8588
rect 11432 8532 11488 8588
rect 11488 8532 11492 8588
rect 11428 8528 11492 8532
rect 11508 8588 11572 8592
rect 11508 8532 11512 8588
rect 11512 8532 11568 8588
rect 11568 8532 11572 8588
rect 11508 8528 11572 8532
rect 11588 8588 11652 8592
rect 11588 8532 11592 8588
rect 11592 8532 11648 8588
rect 11648 8532 11652 8588
rect 11588 8528 11652 8532
rect 18278 8588 18342 8592
rect 18278 8532 18282 8588
rect 18282 8532 18338 8588
rect 18338 8532 18342 8588
rect 18278 8528 18342 8532
rect 18358 8588 18422 8592
rect 18358 8532 18362 8588
rect 18362 8532 18418 8588
rect 18418 8532 18422 8588
rect 18358 8528 18422 8532
rect 18438 8588 18502 8592
rect 18438 8532 18442 8588
rect 18442 8532 18498 8588
rect 18498 8532 18502 8588
rect 18438 8528 18502 8532
rect 18518 8588 18582 8592
rect 18518 8532 18522 8588
rect 18522 8532 18578 8588
rect 18578 8532 18582 8588
rect 18518 8528 18582 8532
rect 7882 8044 7946 8048
rect 7882 7988 7886 8044
rect 7886 7988 7942 8044
rect 7942 7988 7946 8044
rect 7882 7984 7946 7988
rect 7962 8044 8026 8048
rect 7962 7988 7966 8044
rect 7966 7988 8022 8044
rect 8022 7988 8026 8044
rect 7962 7984 8026 7988
rect 8042 8044 8106 8048
rect 8042 7988 8046 8044
rect 8046 7988 8102 8044
rect 8102 7988 8106 8044
rect 8042 7984 8106 7988
rect 8122 8044 8186 8048
rect 8122 7988 8126 8044
rect 8126 7988 8182 8044
rect 8182 7988 8186 8044
rect 8122 7984 8186 7988
rect 14813 8044 14877 8048
rect 14813 7988 14817 8044
rect 14817 7988 14873 8044
rect 14873 7988 14877 8044
rect 14813 7984 14877 7988
rect 14893 8044 14957 8048
rect 14893 7988 14897 8044
rect 14897 7988 14953 8044
rect 14953 7988 14957 8044
rect 14893 7984 14957 7988
rect 14973 8044 15037 8048
rect 14973 7988 14977 8044
rect 14977 7988 15033 8044
rect 15033 7988 15037 8044
rect 14973 7984 15037 7988
rect 15053 8044 15117 8048
rect 15053 7988 15057 8044
rect 15057 7988 15113 8044
rect 15113 7988 15117 8044
rect 15053 7984 15117 7988
rect 4417 7500 4481 7504
rect 4417 7444 4421 7500
rect 4421 7444 4477 7500
rect 4477 7444 4481 7500
rect 4417 7440 4481 7444
rect 4497 7500 4561 7504
rect 4497 7444 4501 7500
rect 4501 7444 4557 7500
rect 4557 7444 4561 7500
rect 4497 7440 4561 7444
rect 4577 7500 4641 7504
rect 4577 7444 4581 7500
rect 4581 7444 4637 7500
rect 4637 7444 4641 7500
rect 4577 7440 4641 7444
rect 4657 7500 4721 7504
rect 4657 7444 4661 7500
rect 4661 7444 4717 7500
rect 4717 7444 4721 7500
rect 4657 7440 4721 7444
rect 11348 7500 11412 7504
rect 11348 7444 11352 7500
rect 11352 7444 11408 7500
rect 11408 7444 11412 7500
rect 11348 7440 11412 7444
rect 11428 7500 11492 7504
rect 11428 7444 11432 7500
rect 11432 7444 11488 7500
rect 11488 7444 11492 7500
rect 11428 7440 11492 7444
rect 11508 7500 11572 7504
rect 11508 7444 11512 7500
rect 11512 7444 11568 7500
rect 11568 7444 11572 7500
rect 11508 7440 11572 7444
rect 11588 7500 11652 7504
rect 11588 7444 11592 7500
rect 11592 7444 11648 7500
rect 11648 7444 11652 7500
rect 11588 7440 11652 7444
rect 18278 7500 18342 7504
rect 18278 7444 18282 7500
rect 18282 7444 18338 7500
rect 18338 7444 18342 7500
rect 18278 7440 18342 7444
rect 18358 7500 18422 7504
rect 18358 7444 18362 7500
rect 18362 7444 18418 7500
rect 18418 7444 18422 7500
rect 18358 7440 18422 7444
rect 18438 7500 18502 7504
rect 18438 7444 18442 7500
rect 18442 7444 18498 7500
rect 18498 7444 18502 7500
rect 18438 7440 18502 7444
rect 18518 7500 18582 7504
rect 18518 7444 18522 7500
rect 18522 7444 18578 7500
rect 18578 7444 18582 7500
rect 18518 7440 18582 7444
rect 7882 6956 7946 6960
rect 7882 6900 7886 6956
rect 7886 6900 7942 6956
rect 7942 6900 7946 6956
rect 7882 6896 7946 6900
rect 7962 6956 8026 6960
rect 7962 6900 7966 6956
rect 7966 6900 8022 6956
rect 8022 6900 8026 6956
rect 7962 6896 8026 6900
rect 8042 6956 8106 6960
rect 8042 6900 8046 6956
rect 8046 6900 8102 6956
rect 8102 6900 8106 6956
rect 8042 6896 8106 6900
rect 8122 6956 8186 6960
rect 8122 6900 8126 6956
rect 8126 6900 8182 6956
rect 8182 6900 8186 6956
rect 8122 6896 8186 6900
rect 14813 6956 14877 6960
rect 14813 6900 14817 6956
rect 14817 6900 14873 6956
rect 14873 6900 14877 6956
rect 14813 6896 14877 6900
rect 14893 6956 14957 6960
rect 14893 6900 14897 6956
rect 14897 6900 14953 6956
rect 14953 6900 14957 6956
rect 14893 6896 14957 6900
rect 14973 6956 15037 6960
rect 14973 6900 14977 6956
rect 14977 6900 15033 6956
rect 15033 6900 15037 6956
rect 14973 6896 15037 6900
rect 15053 6956 15117 6960
rect 15053 6900 15057 6956
rect 15057 6900 15113 6956
rect 15113 6900 15117 6956
rect 15053 6896 15117 6900
rect 4417 6412 4481 6416
rect 4417 6356 4421 6412
rect 4421 6356 4477 6412
rect 4477 6356 4481 6412
rect 4417 6352 4481 6356
rect 4497 6412 4561 6416
rect 4497 6356 4501 6412
rect 4501 6356 4557 6412
rect 4557 6356 4561 6412
rect 4497 6352 4561 6356
rect 4577 6412 4641 6416
rect 4577 6356 4581 6412
rect 4581 6356 4637 6412
rect 4637 6356 4641 6412
rect 4577 6352 4641 6356
rect 4657 6412 4721 6416
rect 4657 6356 4661 6412
rect 4661 6356 4717 6412
rect 4717 6356 4721 6412
rect 4657 6352 4721 6356
rect 11348 6412 11412 6416
rect 11348 6356 11352 6412
rect 11352 6356 11408 6412
rect 11408 6356 11412 6412
rect 11348 6352 11412 6356
rect 11428 6412 11492 6416
rect 11428 6356 11432 6412
rect 11432 6356 11488 6412
rect 11488 6356 11492 6412
rect 11428 6352 11492 6356
rect 11508 6412 11572 6416
rect 11508 6356 11512 6412
rect 11512 6356 11568 6412
rect 11568 6356 11572 6412
rect 11508 6352 11572 6356
rect 11588 6412 11652 6416
rect 11588 6356 11592 6412
rect 11592 6356 11648 6412
rect 11648 6356 11652 6412
rect 11588 6352 11652 6356
rect 18278 6412 18342 6416
rect 18278 6356 18282 6412
rect 18282 6356 18338 6412
rect 18338 6356 18342 6412
rect 18278 6352 18342 6356
rect 18358 6412 18422 6416
rect 18358 6356 18362 6412
rect 18362 6356 18418 6412
rect 18418 6356 18422 6412
rect 18358 6352 18422 6356
rect 18438 6412 18502 6416
rect 18438 6356 18442 6412
rect 18442 6356 18498 6412
rect 18498 6356 18502 6412
rect 18438 6352 18502 6356
rect 18518 6412 18582 6416
rect 18518 6356 18522 6412
rect 18522 6356 18578 6412
rect 18578 6356 18582 6412
rect 18518 6352 18582 6356
rect 7882 5868 7946 5872
rect 7882 5812 7886 5868
rect 7886 5812 7942 5868
rect 7942 5812 7946 5868
rect 7882 5808 7946 5812
rect 7962 5868 8026 5872
rect 7962 5812 7966 5868
rect 7966 5812 8022 5868
rect 8022 5812 8026 5868
rect 7962 5808 8026 5812
rect 8042 5868 8106 5872
rect 8042 5812 8046 5868
rect 8046 5812 8102 5868
rect 8102 5812 8106 5868
rect 8042 5808 8106 5812
rect 8122 5868 8186 5872
rect 8122 5812 8126 5868
rect 8126 5812 8182 5868
rect 8182 5812 8186 5868
rect 8122 5808 8186 5812
rect 14813 5868 14877 5872
rect 14813 5812 14817 5868
rect 14817 5812 14873 5868
rect 14873 5812 14877 5868
rect 14813 5808 14877 5812
rect 14893 5868 14957 5872
rect 14893 5812 14897 5868
rect 14897 5812 14953 5868
rect 14953 5812 14957 5868
rect 14893 5808 14957 5812
rect 14973 5868 15037 5872
rect 14973 5812 14977 5868
rect 14977 5812 15033 5868
rect 15033 5812 15037 5868
rect 14973 5808 15037 5812
rect 15053 5868 15117 5872
rect 15053 5812 15057 5868
rect 15057 5812 15113 5868
rect 15113 5812 15117 5868
rect 15053 5808 15117 5812
rect 4417 5324 4481 5328
rect 4417 5268 4421 5324
rect 4421 5268 4477 5324
rect 4477 5268 4481 5324
rect 4417 5264 4481 5268
rect 4497 5324 4561 5328
rect 4497 5268 4501 5324
rect 4501 5268 4557 5324
rect 4557 5268 4561 5324
rect 4497 5264 4561 5268
rect 4577 5324 4641 5328
rect 4577 5268 4581 5324
rect 4581 5268 4637 5324
rect 4637 5268 4641 5324
rect 4577 5264 4641 5268
rect 4657 5324 4721 5328
rect 4657 5268 4661 5324
rect 4661 5268 4717 5324
rect 4717 5268 4721 5324
rect 4657 5264 4721 5268
rect 11348 5324 11412 5328
rect 11348 5268 11352 5324
rect 11352 5268 11408 5324
rect 11408 5268 11412 5324
rect 11348 5264 11412 5268
rect 11428 5324 11492 5328
rect 11428 5268 11432 5324
rect 11432 5268 11488 5324
rect 11488 5268 11492 5324
rect 11428 5264 11492 5268
rect 11508 5324 11572 5328
rect 11508 5268 11512 5324
rect 11512 5268 11568 5324
rect 11568 5268 11572 5324
rect 11508 5264 11572 5268
rect 11588 5324 11652 5328
rect 11588 5268 11592 5324
rect 11592 5268 11648 5324
rect 11648 5268 11652 5324
rect 11588 5264 11652 5268
rect 18278 5324 18342 5328
rect 18278 5268 18282 5324
rect 18282 5268 18338 5324
rect 18338 5268 18342 5324
rect 18278 5264 18342 5268
rect 18358 5324 18422 5328
rect 18358 5268 18362 5324
rect 18362 5268 18418 5324
rect 18418 5268 18422 5324
rect 18358 5264 18422 5268
rect 18438 5324 18502 5328
rect 18438 5268 18442 5324
rect 18442 5268 18498 5324
rect 18498 5268 18502 5324
rect 18438 5264 18502 5268
rect 18518 5324 18582 5328
rect 18518 5268 18522 5324
rect 18522 5268 18578 5324
rect 18578 5268 18582 5324
rect 18518 5264 18582 5268
rect 7882 4780 7946 4784
rect 7882 4724 7886 4780
rect 7886 4724 7942 4780
rect 7942 4724 7946 4780
rect 7882 4720 7946 4724
rect 7962 4780 8026 4784
rect 7962 4724 7966 4780
rect 7966 4724 8022 4780
rect 8022 4724 8026 4780
rect 7962 4720 8026 4724
rect 8042 4780 8106 4784
rect 8042 4724 8046 4780
rect 8046 4724 8102 4780
rect 8102 4724 8106 4780
rect 8042 4720 8106 4724
rect 8122 4780 8186 4784
rect 8122 4724 8126 4780
rect 8126 4724 8182 4780
rect 8182 4724 8186 4780
rect 8122 4720 8186 4724
rect 14813 4780 14877 4784
rect 14813 4724 14817 4780
rect 14817 4724 14873 4780
rect 14873 4724 14877 4780
rect 14813 4720 14877 4724
rect 14893 4780 14957 4784
rect 14893 4724 14897 4780
rect 14897 4724 14953 4780
rect 14953 4724 14957 4780
rect 14893 4720 14957 4724
rect 14973 4780 15037 4784
rect 14973 4724 14977 4780
rect 14977 4724 15033 4780
rect 15033 4724 15037 4780
rect 14973 4720 15037 4724
rect 15053 4780 15117 4784
rect 15053 4724 15057 4780
rect 15057 4724 15113 4780
rect 15113 4724 15117 4780
rect 15053 4720 15117 4724
rect 4417 4236 4481 4240
rect 4417 4180 4421 4236
rect 4421 4180 4477 4236
rect 4477 4180 4481 4236
rect 4417 4176 4481 4180
rect 4497 4236 4561 4240
rect 4497 4180 4501 4236
rect 4501 4180 4557 4236
rect 4557 4180 4561 4236
rect 4497 4176 4561 4180
rect 4577 4236 4641 4240
rect 4577 4180 4581 4236
rect 4581 4180 4637 4236
rect 4637 4180 4641 4236
rect 4577 4176 4641 4180
rect 4657 4236 4721 4240
rect 4657 4180 4661 4236
rect 4661 4180 4717 4236
rect 4717 4180 4721 4236
rect 4657 4176 4721 4180
rect 11348 4236 11412 4240
rect 11348 4180 11352 4236
rect 11352 4180 11408 4236
rect 11408 4180 11412 4236
rect 11348 4176 11412 4180
rect 11428 4236 11492 4240
rect 11428 4180 11432 4236
rect 11432 4180 11488 4236
rect 11488 4180 11492 4236
rect 11428 4176 11492 4180
rect 11508 4236 11572 4240
rect 11508 4180 11512 4236
rect 11512 4180 11568 4236
rect 11568 4180 11572 4236
rect 11508 4176 11572 4180
rect 11588 4236 11652 4240
rect 11588 4180 11592 4236
rect 11592 4180 11648 4236
rect 11648 4180 11652 4236
rect 11588 4176 11652 4180
rect 18278 4236 18342 4240
rect 18278 4180 18282 4236
rect 18282 4180 18338 4236
rect 18338 4180 18342 4236
rect 18278 4176 18342 4180
rect 18358 4236 18422 4240
rect 18358 4180 18362 4236
rect 18362 4180 18418 4236
rect 18418 4180 18422 4236
rect 18358 4176 18422 4180
rect 18438 4236 18502 4240
rect 18438 4180 18442 4236
rect 18442 4180 18498 4236
rect 18498 4180 18502 4236
rect 18438 4176 18502 4180
rect 18518 4236 18582 4240
rect 18518 4180 18522 4236
rect 18522 4180 18578 4236
rect 18578 4180 18582 4236
rect 18518 4176 18582 4180
rect 7882 3692 7946 3696
rect 7882 3636 7886 3692
rect 7886 3636 7942 3692
rect 7942 3636 7946 3692
rect 7882 3632 7946 3636
rect 7962 3692 8026 3696
rect 7962 3636 7966 3692
rect 7966 3636 8022 3692
rect 8022 3636 8026 3692
rect 7962 3632 8026 3636
rect 8042 3692 8106 3696
rect 8042 3636 8046 3692
rect 8046 3636 8102 3692
rect 8102 3636 8106 3692
rect 8042 3632 8106 3636
rect 8122 3692 8186 3696
rect 8122 3636 8126 3692
rect 8126 3636 8182 3692
rect 8182 3636 8186 3692
rect 8122 3632 8186 3636
rect 14813 3692 14877 3696
rect 14813 3636 14817 3692
rect 14817 3636 14873 3692
rect 14873 3636 14877 3692
rect 14813 3632 14877 3636
rect 14893 3692 14957 3696
rect 14893 3636 14897 3692
rect 14897 3636 14953 3692
rect 14953 3636 14957 3692
rect 14893 3632 14957 3636
rect 14973 3692 15037 3696
rect 14973 3636 14977 3692
rect 14977 3636 15033 3692
rect 15033 3636 15037 3692
rect 14973 3632 15037 3636
rect 15053 3692 15117 3696
rect 15053 3636 15057 3692
rect 15057 3636 15113 3692
rect 15113 3636 15117 3692
rect 15053 3632 15117 3636
rect 4417 3148 4481 3152
rect 4417 3092 4421 3148
rect 4421 3092 4477 3148
rect 4477 3092 4481 3148
rect 4417 3088 4481 3092
rect 4497 3148 4561 3152
rect 4497 3092 4501 3148
rect 4501 3092 4557 3148
rect 4557 3092 4561 3148
rect 4497 3088 4561 3092
rect 4577 3148 4641 3152
rect 4577 3092 4581 3148
rect 4581 3092 4637 3148
rect 4637 3092 4641 3148
rect 4577 3088 4641 3092
rect 4657 3148 4721 3152
rect 4657 3092 4661 3148
rect 4661 3092 4717 3148
rect 4717 3092 4721 3148
rect 4657 3088 4721 3092
rect 11348 3148 11412 3152
rect 11348 3092 11352 3148
rect 11352 3092 11408 3148
rect 11408 3092 11412 3148
rect 11348 3088 11412 3092
rect 11428 3148 11492 3152
rect 11428 3092 11432 3148
rect 11432 3092 11488 3148
rect 11488 3092 11492 3148
rect 11428 3088 11492 3092
rect 11508 3148 11572 3152
rect 11508 3092 11512 3148
rect 11512 3092 11568 3148
rect 11568 3092 11572 3148
rect 11508 3088 11572 3092
rect 11588 3148 11652 3152
rect 11588 3092 11592 3148
rect 11592 3092 11648 3148
rect 11648 3092 11652 3148
rect 11588 3088 11652 3092
rect 18278 3148 18342 3152
rect 18278 3092 18282 3148
rect 18282 3092 18338 3148
rect 18338 3092 18342 3148
rect 18278 3088 18342 3092
rect 18358 3148 18422 3152
rect 18358 3092 18362 3148
rect 18362 3092 18418 3148
rect 18418 3092 18422 3148
rect 18358 3088 18422 3092
rect 18438 3148 18502 3152
rect 18438 3092 18442 3148
rect 18442 3092 18498 3148
rect 18498 3092 18502 3148
rect 18438 3088 18502 3092
rect 18518 3148 18582 3152
rect 18518 3092 18522 3148
rect 18522 3092 18578 3148
rect 18578 3092 18582 3148
rect 18518 3088 18582 3092
rect 7882 2604 7946 2608
rect 7882 2548 7886 2604
rect 7886 2548 7942 2604
rect 7942 2548 7946 2604
rect 7882 2544 7946 2548
rect 7962 2604 8026 2608
rect 7962 2548 7966 2604
rect 7966 2548 8022 2604
rect 8022 2548 8026 2604
rect 7962 2544 8026 2548
rect 8042 2604 8106 2608
rect 8042 2548 8046 2604
rect 8046 2548 8102 2604
rect 8102 2548 8106 2604
rect 8042 2544 8106 2548
rect 8122 2604 8186 2608
rect 8122 2548 8126 2604
rect 8126 2548 8182 2604
rect 8182 2548 8186 2604
rect 8122 2544 8186 2548
rect 14813 2604 14877 2608
rect 14813 2548 14817 2604
rect 14817 2548 14873 2604
rect 14873 2548 14877 2604
rect 14813 2544 14877 2548
rect 14893 2604 14957 2608
rect 14893 2548 14897 2604
rect 14897 2548 14953 2604
rect 14953 2548 14957 2604
rect 14893 2544 14957 2548
rect 14973 2604 15037 2608
rect 14973 2548 14977 2604
rect 14977 2548 15033 2604
rect 15033 2548 15037 2604
rect 14973 2544 15037 2548
rect 15053 2604 15117 2608
rect 15053 2548 15057 2604
rect 15057 2548 15113 2604
rect 15113 2548 15117 2604
rect 15053 2544 15117 2548
rect 4417 2060 4481 2064
rect 4417 2004 4421 2060
rect 4421 2004 4477 2060
rect 4477 2004 4481 2060
rect 4417 2000 4481 2004
rect 4497 2060 4561 2064
rect 4497 2004 4501 2060
rect 4501 2004 4557 2060
rect 4557 2004 4561 2060
rect 4497 2000 4561 2004
rect 4577 2060 4641 2064
rect 4577 2004 4581 2060
rect 4581 2004 4637 2060
rect 4637 2004 4641 2060
rect 4577 2000 4641 2004
rect 4657 2060 4721 2064
rect 4657 2004 4661 2060
rect 4661 2004 4717 2060
rect 4717 2004 4721 2060
rect 4657 2000 4721 2004
rect 11348 2060 11412 2064
rect 11348 2004 11352 2060
rect 11352 2004 11408 2060
rect 11408 2004 11412 2060
rect 11348 2000 11412 2004
rect 11428 2060 11492 2064
rect 11428 2004 11432 2060
rect 11432 2004 11488 2060
rect 11488 2004 11492 2060
rect 11428 2000 11492 2004
rect 11508 2060 11572 2064
rect 11508 2004 11512 2060
rect 11512 2004 11568 2060
rect 11568 2004 11572 2060
rect 11508 2000 11572 2004
rect 11588 2060 11652 2064
rect 11588 2004 11592 2060
rect 11592 2004 11648 2060
rect 11648 2004 11652 2060
rect 11588 2000 11652 2004
rect 18278 2060 18342 2064
rect 18278 2004 18282 2060
rect 18282 2004 18338 2060
rect 18338 2004 18342 2060
rect 18278 2000 18342 2004
rect 18358 2060 18422 2064
rect 18358 2004 18362 2060
rect 18362 2004 18418 2060
rect 18418 2004 18422 2060
rect 18358 2000 18422 2004
rect 18438 2060 18502 2064
rect 18438 2004 18442 2060
rect 18442 2004 18498 2060
rect 18498 2004 18502 2060
rect 18438 2000 18502 2004
rect 18518 2060 18582 2064
rect 18518 2004 18522 2060
rect 18522 2004 18578 2060
rect 18578 2004 18582 2060
rect 18518 2000 18582 2004
<< metal4 >>
rect 4409 20560 4729 20576
rect 4409 20496 4417 20560
rect 4481 20496 4497 20560
rect 4561 20496 4577 20560
rect 4641 20496 4657 20560
rect 4721 20496 4729 20560
rect 4409 19472 4729 20496
rect 4409 19408 4417 19472
rect 4481 19408 4497 19472
rect 4561 19408 4577 19472
rect 4641 19408 4657 19472
rect 4721 19408 4729 19472
rect 4409 18384 4729 19408
rect 4409 18320 4417 18384
rect 4481 18320 4497 18384
rect 4561 18320 4577 18384
rect 4641 18320 4657 18384
rect 4721 18320 4729 18384
rect 4409 17296 4729 18320
rect 4409 17232 4417 17296
rect 4481 17232 4497 17296
rect 4561 17232 4577 17296
rect 4641 17232 4657 17296
rect 4721 17232 4729 17296
rect 4409 16208 4729 17232
rect 4409 16144 4417 16208
rect 4481 16144 4497 16208
rect 4561 16144 4577 16208
rect 4641 16144 4657 16208
rect 4721 16144 4729 16208
rect 4409 15120 4729 16144
rect 4409 15056 4417 15120
rect 4481 15056 4497 15120
rect 4561 15056 4577 15120
rect 4641 15056 4657 15120
rect 4721 15056 4729 15120
rect 4409 14032 4729 15056
rect 4409 13968 4417 14032
rect 4481 13968 4497 14032
rect 4561 13968 4577 14032
rect 4641 13968 4657 14032
rect 4721 13968 4729 14032
rect 4409 12944 4729 13968
rect 4409 12880 4417 12944
rect 4481 12880 4497 12944
rect 4561 12880 4577 12944
rect 4641 12880 4657 12944
rect 4721 12880 4729 12944
rect 4409 11856 4729 12880
rect 4409 11792 4417 11856
rect 4481 11792 4497 11856
rect 4561 11792 4577 11856
rect 4641 11792 4657 11856
rect 4721 11792 4729 11856
rect 4409 10768 4729 11792
rect 4409 10704 4417 10768
rect 4481 10704 4497 10768
rect 4561 10704 4577 10768
rect 4641 10704 4657 10768
rect 4721 10704 4729 10768
rect 4409 9680 4729 10704
rect 4409 9616 4417 9680
rect 4481 9616 4497 9680
rect 4561 9616 4577 9680
rect 4641 9616 4657 9680
rect 4721 9616 4729 9680
rect 4409 8592 4729 9616
rect 4409 8528 4417 8592
rect 4481 8528 4497 8592
rect 4561 8528 4577 8592
rect 4641 8528 4657 8592
rect 4721 8528 4729 8592
rect 4409 7504 4729 8528
rect 4409 7440 4417 7504
rect 4481 7440 4497 7504
rect 4561 7440 4577 7504
rect 4641 7440 4657 7504
rect 4721 7440 4729 7504
rect 4409 6416 4729 7440
rect 4409 6352 4417 6416
rect 4481 6352 4497 6416
rect 4561 6352 4577 6416
rect 4641 6352 4657 6416
rect 4721 6352 4729 6416
rect 4409 5328 4729 6352
rect 4409 5264 4417 5328
rect 4481 5264 4497 5328
rect 4561 5264 4577 5328
rect 4641 5264 4657 5328
rect 4721 5264 4729 5328
rect 4409 4240 4729 5264
rect 4409 4176 4417 4240
rect 4481 4176 4497 4240
rect 4561 4176 4577 4240
rect 4641 4176 4657 4240
rect 4721 4176 4729 4240
rect 4409 3152 4729 4176
rect 4409 3088 4417 3152
rect 4481 3088 4497 3152
rect 4561 3088 4577 3152
rect 4641 3088 4657 3152
rect 4721 3088 4729 3152
rect 4409 2064 4729 3088
rect 4409 2000 4417 2064
rect 4481 2000 4497 2064
rect 4561 2000 4577 2064
rect 4641 2000 4657 2064
rect 4721 2000 4729 2064
rect 4409 1984 4729 2000
rect 7874 20016 8195 20576
rect 7874 19952 7882 20016
rect 7946 19952 7962 20016
rect 8026 19952 8042 20016
rect 8106 19952 8122 20016
rect 8186 19952 8195 20016
rect 7874 18928 8195 19952
rect 7874 18864 7882 18928
rect 7946 18864 7962 18928
rect 8026 18864 8042 18928
rect 8106 18864 8122 18928
rect 8186 18864 8195 18928
rect 7874 17840 8195 18864
rect 7874 17776 7882 17840
rect 7946 17776 7962 17840
rect 8026 17776 8042 17840
rect 8106 17776 8122 17840
rect 8186 17776 8195 17840
rect 7874 16752 8195 17776
rect 7874 16688 7882 16752
rect 7946 16688 7962 16752
rect 8026 16688 8042 16752
rect 8106 16688 8122 16752
rect 8186 16688 8195 16752
rect 7874 15664 8195 16688
rect 7874 15600 7882 15664
rect 7946 15600 7962 15664
rect 8026 15600 8042 15664
rect 8106 15600 8122 15664
rect 8186 15600 8195 15664
rect 7874 14576 8195 15600
rect 7874 14512 7882 14576
rect 7946 14512 7962 14576
rect 8026 14512 8042 14576
rect 8106 14512 8122 14576
rect 8186 14512 8195 14576
rect 7874 13488 8195 14512
rect 7874 13424 7882 13488
rect 7946 13424 7962 13488
rect 8026 13424 8042 13488
rect 8106 13424 8122 13488
rect 8186 13424 8195 13488
rect 7874 12400 8195 13424
rect 7874 12336 7882 12400
rect 7946 12336 7962 12400
rect 8026 12336 8042 12400
rect 8106 12336 8122 12400
rect 8186 12336 8195 12400
rect 7874 11312 8195 12336
rect 7874 11248 7882 11312
rect 7946 11248 7962 11312
rect 8026 11248 8042 11312
rect 8106 11248 8122 11312
rect 8186 11248 8195 11312
rect 7874 10224 8195 11248
rect 7874 10160 7882 10224
rect 7946 10160 7962 10224
rect 8026 10160 8042 10224
rect 8106 10160 8122 10224
rect 8186 10160 8195 10224
rect 7874 9136 8195 10160
rect 7874 9072 7882 9136
rect 7946 9072 7962 9136
rect 8026 9072 8042 9136
rect 8106 9072 8122 9136
rect 8186 9072 8195 9136
rect 7874 8048 8195 9072
rect 7874 7984 7882 8048
rect 7946 7984 7962 8048
rect 8026 7984 8042 8048
rect 8106 7984 8122 8048
rect 8186 7984 8195 8048
rect 7874 6960 8195 7984
rect 7874 6896 7882 6960
rect 7946 6896 7962 6960
rect 8026 6896 8042 6960
rect 8106 6896 8122 6960
rect 8186 6896 8195 6960
rect 7874 5872 8195 6896
rect 7874 5808 7882 5872
rect 7946 5808 7962 5872
rect 8026 5808 8042 5872
rect 8106 5808 8122 5872
rect 8186 5808 8195 5872
rect 7874 4784 8195 5808
rect 7874 4720 7882 4784
rect 7946 4720 7962 4784
rect 8026 4720 8042 4784
rect 8106 4720 8122 4784
rect 8186 4720 8195 4784
rect 7874 3696 8195 4720
rect 7874 3632 7882 3696
rect 7946 3632 7962 3696
rect 8026 3632 8042 3696
rect 8106 3632 8122 3696
rect 8186 3632 8195 3696
rect 7874 2608 8195 3632
rect 7874 2544 7882 2608
rect 7946 2544 7962 2608
rect 8026 2544 8042 2608
rect 8106 2544 8122 2608
rect 8186 2544 8195 2608
rect 7874 1984 8195 2544
rect 11340 20560 11660 20576
rect 11340 20496 11348 20560
rect 11412 20496 11428 20560
rect 11492 20496 11508 20560
rect 11572 20496 11588 20560
rect 11652 20496 11660 20560
rect 11340 19472 11660 20496
rect 11340 19408 11348 19472
rect 11412 19408 11428 19472
rect 11492 19408 11508 19472
rect 11572 19408 11588 19472
rect 11652 19408 11660 19472
rect 11340 18384 11660 19408
rect 11340 18320 11348 18384
rect 11412 18320 11428 18384
rect 11492 18320 11508 18384
rect 11572 18320 11588 18384
rect 11652 18320 11660 18384
rect 11340 17296 11660 18320
rect 11340 17232 11348 17296
rect 11412 17232 11428 17296
rect 11492 17232 11508 17296
rect 11572 17232 11588 17296
rect 11652 17232 11660 17296
rect 11340 16208 11660 17232
rect 11340 16144 11348 16208
rect 11412 16144 11428 16208
rect 11492 16144 11508 16208
rect 11572 16144 11588 16208
rect 11652 16144 11660 16208
rect 11340 15120 11660 16144
rect 11340 15056 11348 15120
rect 11412 15056 11428 15120
rect 11492 15056 11508 15120
rect 11572 15056 11588 15120
rect 11652 15056 11660 15120
rect 11340 14032 11660 15056
rect 11340 13968 11348 14032
rect 11412 13968 11428 14032
rect 11492 13968 11508 14032
rect 11572 13968 11588 14032
rect 11652 13968 11660 14032
rect 11340 12944 11660 13968
rect 11340 12880 11348 12944
rect 11412 12880 11428 12944
rect 11492 12880 11508 12944
rect 11572 12880 11588 12944
rect 11652 12880 11660 12944
rect 11340 11856 11660 12880
rect 11340 11792 11348 11856
rect 11412 11792 11428 11856
rect 11492 11792 11508 11856
rect 11572 11792 11588 11856
rect 11652 11792 11660 11856
rect 11340 10768 11660 11792
rect 11340 10704 11348 10768
rect 11412 10704 11428 10768
rect 11492 10704 11508 10768
rect 11572 10704 11588 10768
rect 11652 10704 11660 10768
rect 11340 9680 11660 10704
rect 11340 9616 11348 9680
rect 11412 9616 11428 9680
rect 11492 9616 11508 9680
rect 11572 9616 11588 9680
rect 11652 9616 11660 9680
rect 11340 8592 11660 9616
rect 11340 8528 11348 8592
rect 11412 8528 11428 8592
rect 11492 8528 11508 8592
rect 11572 8528 11588 8592
rect 11652 8528 11660 8592
rect 11340 7504 11660 8528
rect 11340 7440 11348 7504
rect 11412 7440 11428 7504
rect 11492 7440 11508 7504
rect 11572 7440 11588 7504
rect 11652 7440 11660 7504
rect 11340 6416 11660 7440
rect 11340 6352 11348 6416
rect 11412 6352 11428 6416
rect 11492 6352 11508 6416
rect 11572 6352 11588 6416
rect 11652 6352 11660 6416
rect 11340 5328 11660 6352
rect 11340 5264 11348 5328
rect 11412 5264 11428 5328
rect 11492 5264 11508 5328
rect 11572 5264 11588 5328
rect 11652 5264 11660 5328
rect 11340 4240 11660 5264
rect 11340 4176 11348 4240
rect 11412 4176 11428 4240
rect 11492 4176 11508 4240
rect 11572 4176 11588 4240
rect 11652 4176 11660 4240
rect 11340 3152 11660 4176
rect 11340 3088 11348 3152
rect 11412 3088 11428 3152
rect 11492 3088 11508 3152
rect 11572 3088 11588 3152
rect 11652 3088 11660 3152
rect 11340 2064 11660 3088
rect 11340 2000 11348 2064
rect 11412 2000 11428 2064
rect 11492 2000 11508 2064
rect 11572 2000 11588 2064
rect 11652 2000 11660 2064
rect 11340 1984 11660 2000
rect 14805 20016 15125 20576
rect 14805 19952 14813 20016
rect 14877 19952 14893 20016
rect 14957 19952 14973 20016
rect 15037 19952 15053 20016
rect 15117 19952 15125 20016
rect 14805 18928 15125 19952
rect 14805 18864 14813 18928
rect 14877 18864 14893 18928
rect 14957 18864 14973 18928
rect 15037 18864 15053 18928
rect 15117 18864 15125 18928
rect 14805 17840 15125 18864
rect 14805 17776 14813 17840
rect 14877 17776 14893 17840
rect 14957 17776 14973 17840
rect 15037 17776 15053 17840
rect 15117 17776 15125 17840
rect 14805 16752 15125 17776
rect 14805 16688 14813 16752
rect 14877 16688 14893 16752
rect 14957 16688 14973 16752
rect 15037 16688 15053 16752
rect 15117 16688 15125 16752
rect 14805 15664 15125 16688
rect 14805 15600 14813 15664
rect 14877 15600 14893 15664
rect 14957 15600 14973 15664
rect 15037 15600 15053 15664
rect 15117 15600 15125 15664
rect 14805 14576 15125 15600
rect 14805 14512 14813 14576
rect 14877 14512 14893 14576
rect 14957 14512 14973 14576
rect 15037 14512 15053 14576
rect 15117 14512 15125 14576
rect 14805 13488 15125 14512
rect 14805 13424 14813 13488
rect 14877 13424 14893 13488
rect 14957 13424 14973 13488
rect 15037 13424 15053 13488
rect 15117 13424 15125 13488
rect 14805 12400 15125 13424
rect 14805 12336 14813 12400
rect 14877 12336 14893 12400
rect 14957 12336 14973 12400
rect 15037 12336 15053 12400
rect 15117 12336 15125 12400
rect 14805 11312 15125 12336
rect 14805 11248 14813 11312
rect 14877 11248 14893 11312
rect 14957 11248 14973 11312
rect 15037 11248 15053 11312
rect 15117 11248 15125 11312
rect 14805 10224 15125 11248
rect 14805 10160 14813 10224
rect 14877 10160 14893 10224
rect 14957 10160 14973 10224
rect 15037 10160 15053 10224
rect 15117 10160 15125 10224
rect 14805 9136 15125 10160
rect 14805 9072 14813 9136
rect 14877 9072 14893 9136
rect 14957 9072 14973 9136
rect 15037 9072 15053 9136
rect 15117 9072 15125 9136
rect 14805 8048 15125 9072
rect 14805 7984 14813 8048
rect 14877 7984 14893 8048
rect 14957 7984 14973 8048
rect 15037 7984 15053 8048
rect 15117 7984 15125 8048
rect 14805 6960 15125 7984
rect 14805 6896 14813 6960
rect 14877 6896 14893 6960
rect 14957 6896 14973 6960
rect 15037 6896 15053 6960
rect 15117 6896 15125 6960
rect 14805 5872 15125 6896
rect 14805 5808 14813 5872
rect 14877 5808 14893 5872
rect 14957 5808 14973 5872
rect 15037 5808 15053 5872
rect 15117 5808 15125 5872
rect 14805 4784 15125 5808
rect 14805 4720 14813 4784
rect 14877 4720 14893 4784
rect 14957 4720 14973 4784
rect 15037 4720 15053 4784
rect 15117 4720 15125 4784
rect 14805 3696 15125 4720
rect 14805 3632 14813 3696
rect 14877 3632 14893 3696
rect 14957 3632 14973 3696
rect 15037 3632 15053 3696
rect 15117 3632 15125 3696
rect 14805 2608 15125 3632
rect 14805 2544 14813 2608
rect 14877 2544 14893 2608
rect 14957 2544 14973 2608
rect 15037 2544 15053 2608
rect 15117 2544 15125 2608
rect 14805 1984 15125 2544
rect 18270 20560 18590 20576
rect 18270 20496 18278 20560
rect 18342 20496 18358 20560
rect 18422 20496 18438 20560
rect 18502 20496 18518 20560
rect 18582 20496 18590 20560
rect 18270 19472 18590 20496
rect 18270 19408 18278 19472
rect 18342 19408 18358 19472
rect 18422 19408 18438 19472
rect 18502 19408 18518 19472
rect 18582 19408 18590 19472
rect 18270 18384 18590 19408
rect 18827 18724 18893 18725
rect 18827 18660 18828 18724
rect 18892 18660 18893 18724
rect 18827 18659 18893 18660
rect 18270 18320 18278 18384
rect 18342 18320 18358 18384
rect 18422 18320 18438 18384
rect 18502 18320 18518 18384
rect 18582 18320 18590 18384
rect 18270 17296 18590 18320
rect 18270 17232 18278 17296
rect 18342 17232 18358 17296
rect 18422 17232 18438 17296
rect 18502 17232 18518 17296
rect 18582 17232 18590 17296
rect 18270 16208 18590 17232
rect 18830 16957 18890 18659
rect 18827 16956 18893 16957
rect 18827 16892 18828 16956
rect 18892 16892 18893 16956
rect 18827 16891 18893 16892
rect 18270 16144 18278 16208
rect 18342 16144 18358 16208
rect 18422 16144 18438 16208
rect 18502 16144 18518 16208
rect 18582 16144 18590 16208
rect 18270 15120 18590 16144
rect 18270 15056 18278 15120
rect 18342 15056 18358 15120
rect 18422 15056 18438 15120
rect 18502 15056 18518 15120
rect 18582 15056 18590 15120
rect 18270 14032 18590 15056
rect 18270 13968 18278 14032
rect 18342 13968 18358 14032
rect 18422 13968 18438 14032
rect 18502 13968 18518 14032
rect 18582 13968 18590 14032
rect 18270 12944 18590 13968
rect 18270 12880 18278 12944
rect 18342 12880 18358 12944
rect 18422 12880 18438 12944
rect 18502 12880 18518 12944
rect 18582 12880 18590 12944
rect 18270 11856 18590 12880
rect 18270 11792 18278 11856
rect 18342 11792 18358 11856
rect 18422 11792 18438 11856
rect 18502 11792 18518 11856
rect 18582 11792 18590 11856
rect 18270 10768 18590 11792
rect 18270 10704 18278 10768
rect 18342 10704 18358 10768
rect 18422 10704 18438 10768
rect 18502 10704 18518 10768
rect 18582 10704 18590 10768
rect 18270 9680 18590 10704
rect 18270 9616 18278 9680
rect 18342 9616 18358 9680
rect 18422 9616 18438 9680
rect 18502 9616 18518 9680
rect 18582 9616 18590 9680
rect 18270 8592 18590 9616
rect 18270 8528 18278 8592
rect 18342 8528 18358 8592
rect 18422 8528 18438 8592
rect 18502 8528 18518 8592
rect 18582 8528 18590 8592
rect 18270 7504 18590 8528
rect 18270 7440 18278 7504
rect 18342 7440 18358 7504
rect 18422 7440 18438 7504
rect 18502 7440 18518 7504
rect 18582 7440 18590 7504
rect 18270 6416 18590 7440
rect 18270 6352 18278 6416
rect 18342 6352 18358 6416
rect 18422 6352 18438 6416
rect 18502 6352 18518 6416
rect 18582 6352 18590 6416
rect 18270 5328 18590 6352
rect 18270 5264 18278 5328
rect 18342 5264 18358 5328
rect 18422 5264 18438 5328
rect 18502 5264 18518 5328
rect 18582 5264 18590 5328
rect 18270 4240 18590 5264
rect 18270 4176 18278 4240
rect 18342 4176 18358 4240
rect 18422 4176 18438 4240
rect 18502 4176 18518 4240
rect 18582 4176 18590 4240
rect 18270 3152 18590 4176
rect 18270 3088 18278 3152
rect 18342 3088 18358 3152
rect 18422 3088 18438 3152
rect 18502 3088 18518 3152
rect 18582 3088 18590 3152
rect 18270 2064 18590 3088
rect 18270 2000 18278 2064
rect 18342 2000 18358 2064
rect 18422 2000 18438 2064
rect 18502 2000 18518 2064
rect 18582 2000 18590 2064
rect 18270 1984 18590 2000
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 3956 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_32
timestamp 1604681595
transform 1 0 4048 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1604681595
transform 1 0 6808 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1604681595
transform 1 0 5152 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_56
timestamp 1604681595
transform 1 0 6256 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_68
timestamp 1604681595
transform 1 0 7360 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_80
timestamp 1604681595
transform 1 0 8464 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1604681595
transform 1 0 9660 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 9568 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1604681595
transform 1 0 9108 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1604681595
transform 1 0 9660 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1604681595
transform 1 0 12512 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604681595
transform 1 0 10856 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1604681595
transform 1 0 11960 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_105
timestamp 1604681595
transform 1 0 10764 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_117
timestamp 1604681595
transform 1 0 11868 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1604681595
transform 1 0 13708 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_129
timestamp 1604681595
transform 1 0 12972 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_141
timestamp 1604681595
transform 1 0 14076 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1604681595
transform 1 0 15364 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 15180 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1604681595
transform 1 0 14812 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_154
timestamp 1604681595
transform 1 0 15272 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_166
timestamp 1604681595
transform 1 0 16376 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 18216 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604681595
transform 1 0 16560 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604681595
transform 1 0 17664 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_178
timestamp 1604681595
transform 1 0 17480 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604681595
transform 1 0 19412 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_190
timestamp 1604681595
transform 1 0 18584 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_202
timestamp 1604681595
transform 1 0 19688 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 21896 0 -1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 21896 0 1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 21068 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 20792 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604681595
transform 1 0 20516 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 21528 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_215 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 20884 0 1 2576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_39
timestamp 1604681595
transform 1 0 4692 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 6716 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_51
timestamp 1604681595
transform 1 0 5796 0 -1 3664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6532 0 -1 3664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_62
timestamp 1604681595
transform 1 0 6808 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_74
timestamp 1604681595
transform 1 0 7912 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_86
timestamp 1604681595
transform 1 0 9016 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_98
timestamp 1604681595
transform 1 0 10120 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 12328 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_110
timestamp 1604681595
transform 1 0 11224 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1604681595
transform 1 0 12420 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_135
timestamp 1604681595
transform 1 0 13524 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_147
timestamp 1604681595
transform 1 0 14628 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_159
timestamp 1604681595
transform 1 0 15732 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 17940 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_171
timestamp 1604681595
transform 1 0 16836 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_184
timestamp 1604681595
transform 1 0 18032 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_196
timestamp 1604681595
transform 1 0 19136 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_208
timestamp 1604681595
transform 1 0 20240 0 -1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _60_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 20516 0 -1 3664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 21896 0 -1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 3956 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1604681595
transform 1 0 4048 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1604681595
transform 1 0 5152 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_56
timestamp 1604681595
transform 1 0 6256 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_68
timestamp 1604681595
transform 1 0 7360 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_80
timestamp 1604681595
transform 1 0 8464 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 9568 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1604681595
transform 1 0 9660 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_105
timestamp 1604681595
transform 1 0 10764 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_117
timestamp 1604681595
transform 1 0 11868 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_129
timestamp 1604681595
transform 1 0 12972 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_141
timestamp 1604681595
transform 1 0 14076 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 15180 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_154
timestamp 1604681595
transform 1 0 15272 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_166
timestamp 1604681595
transform 1 0 16376 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_178
timestamp 1604681595
transform 1 0 17480 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_190
timestamp 1604681595
transform 1 0 18584 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_202
timestamp 1604681595
transform 1 0 19688 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 21896 0 1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 20792 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_215
timestamp 1604681595
transform 1 0 20884 0 1 3664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_39
timestamp 1604681595
transform 1 0 4692 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 6716 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_51
timestamp 1604681595
transform 1 0 5796 0 -1 4752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1604681595
transform 1 0 6532 0 -1 4752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_62
timestamp 1604681595
transform 1 0 6808 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_74
timestamp 1604681595
transform 1 0 7912 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_86
timestamp 1604681595
transform 1 0 9016 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_98
timestamp 1604681595
transform 1 0 10120 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 12328 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_110
timestamp 1604681595
transform 1 0 11224 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_123
timestamp 1604681595
transform 1 0 12420 0 -1 4752
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 12972 0 -1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_133
timestamp 1604681595
transform 1 0 13340 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_157
timestamp 1604681595
transform 1 0 15548 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 17940 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_169
timestamp 1604681595
transform 1 0 16652 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_181
timestamp 1604681595
transform 1 0 17756 0 -1 4752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_184
timestamp 1604681595
transform 1 0 18032 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_196
timestamp 1604681595
transform 1 0 19136 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_208
timestamp 1604681595
transform 1 0 20240 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 21896 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_220
timestamp 1604681595
transform 1 0 21344 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 3956 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_32
timestamp 1604681595
transform 1 0 4048 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1604681595
transform 1 0 5152 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_56
timestamp 1604681595
transform 1 0 6256 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_68
timestamp 1604681595
transform 1 0 7360 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_80
timestamp 1604681595
transform 1 0 8464 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 9568 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1604681595
transform 1 0 9660 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_105
timestamp 1604681595
transform 1 0 10764 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_117
timestamp 1604681595
transform 1 0 11868 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_129
timestamp 1604681595
transform 1 0 12972 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_141
timestamp 1604681595
transform 1 0 14076 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 15180 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_154
timestamp 1604681595
transform 1 0 15272 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_166
timestamp 1604681595
transform 1 0 16376 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_178
timestamp 1604681595
transform 1 0 17480 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_190
timestamp 1604681595
transform 1 0 18584 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_202
timestamp 1604681595
transform 1 0 19688 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 21896 0 1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 20792 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_215
timestamp 1604681595
transform 1 0 20884 0 1 4752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 3956 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_39
timestamp 1604681595
transform 1 0 4692 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_32
timestamp 1604681595
transform 1 0 4048 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 6716 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_51
timestamp 1604681595
transform 1 0 5796 0 -1 5840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_59
timestamp 1604681595
transform 1 0 6532 0 -1 5840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_62
timestamp 1604681595
transform 1 0 6808 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1604681595
transform 1 0 5152 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_56
timestamp 1604681595
transform 1 0 6256 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_74
timestamp 1604681595
transform 1 0 7912 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_68
timestamp 1604681595
transform 1 0 7360 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1604681595
transform 1 0 8464 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 9568 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_86
timestamp 1604681595
transform 1 0 9016 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_98
timestamp 1604681595
transform 1 0 10120 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1604681595
transform 1 0 9660 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 12328 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_110
timestamp 1604681595
transform 1 0 11224 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1604681595
transform 1 0 12420 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_105
timestamp 1604681595
transform 1 0 10764 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_117
timestamp 1604681595
transform 1 0 11868 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_135
timestamp 1604681595
transform 1 0 13524 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_129
timestamp 1604681595
transform 1 0 12972 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_141
timestamp 1604681595
transform 1 0 14076 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 15180 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_147
timestamp 1604681595
transform 1 0 14628 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_159
timestamp 1604681595
transform 1 0 15732 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_154
timestamp 1604681595
transform 1 0 15272 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_166
timestamp 1604681595
transform 1 0 16376 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 17940 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_171
timestamp 1604681595
transform 1 0 16836 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1604681595
transform 1 0 18032 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_178
timestamp 1604681595
transform 1 0 17480 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1604681595
transform 1 0 19136 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_208
timestamp 1604681595
transform 1 0 20240 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_190
timestamp 1604681595
transform 1 0 18584 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_202
timestamp 1604681595
transform 1 0 19688 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 20516 0 -1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 21896 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 21896 0 1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 20792 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_215
timestamp 1604681595
transform 1 0 20884 0 1 5840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_39
timestamp 1604681595
transform 1 0 4692 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 6716 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_51
timestamp 1604681595
transform 1 0 5796 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_59
timestamp 1604681595
transform 1 0 6532 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_62
timestamp 1604681595
transform 1 0 6808 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7912 0 -1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_90
timestamp 1604681595
transform 1 0 9384 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_102
timestamp 1604681595
transform 1 0 10488 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10764 0 -1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 12328 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_114
timestamp 1604681595
transform 1 0 11592 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1604681595
transform 1 0 12420 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_135
timestamp 1604681595
transform 1 0 13524 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_157
timestamp 1604681595
transform 1 0 15548 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 17940 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_169
timestamp 1604681595
transform 1 0 16652 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_181
timestamp 1604681595
transform 1 0 17756 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_184
timestamp 1604681595
transform 1 0 18032 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 19412 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_196
timestamp 1604681595
transform 1 0 19136 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_203
timestamp 1604681595
transform 1 0 19780 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 20516 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 21896 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 3956 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_32
timestamp 1604681595
transform 1 0 4048 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_44
timestamp 1604681595
transform 1 0 5152 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_56
timestamp 1604681595
transform 1 0 6256 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_68
timestamp 1604681595
transform 1 0 7360 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_80
timestamp 1604681595
transform 1 0 8464 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 9568 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1604681595
transform 1 0 9660 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12788 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_126
timestamp 1604681595
transform 1 0 12696 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_143
timestamp 1604681595
transform 1 0 14260 0 1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 15180 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_151
timestamp 1604681595
transform 1 0 14996 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_154
timestamp 1604681595
transform 1 0 15272 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_166
timestamp 1604681595
transform 1 0 16376 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16468 0 1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_176
timestamp 1604681595
transform 1 0 17296 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_188
timestamp 1604681595
transform 1 0 18400 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_200
timestamp 1604681595
transform 1 0 19504 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 21896 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 20792 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_212
timestamp 1604681595
transform 1 0 20608 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_215
timestamp 1604681595
transform 1 0 20884 0 1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1604681595
transform 1 0 4692 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 6716 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_51
timestamp 1604681595
transform 1 0 5796 0 -1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1604681595
transform 1 0 6532 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_62
timestamp 1604681595
transform 1 0 6808 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_74
timestamp 1604681595
transform 1 0 7912 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9752 0 -1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_86
timestamp 1604681595
transform 1 0 9016 0 -1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 12328 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_110
timestamp 1604681595
transform 1 0 11224 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_123
timestamp 1604681595
transform 1 0 12420 0 -1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _25_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13248 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14260 0 -1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_131
timestamp 1604681595
transform 1 0 13156 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_135
timestamp 1604681595
transform 1 0 13524 0 -1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_159
timestamp 1604681595
transform 1 0 15732 0 -1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 16468 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 17940 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_170
timestamp 1604681595
transform 1 0 16744 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_182
timestamp 1604681595
transform 1 0 17848 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_184
timestamp 1604681595
transform 1 0 18032 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 19412 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_196
timestamp 1604681595
transform 1 0 19136 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_203
timestamp 1604681595
transform 1 0 19780 0 -1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 20516 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 21896 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 3956 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_32
timestamp 1604681595
transform 1 0 4048 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_44
timestamp 1604681595
transform 1 0 5152 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_56
timestamp 1604681595
transform 1 0 6256 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_68
timestamp 1604681595
transform 1 0 7360 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_80
timestamp 1604681595
transform 1 0 8464 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1604681595
transform 1 0 10304 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 9568 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_93
timestamp 1604681595
transform 1 0 9660 0 1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_99
timestamp 1604681595
transform 1 0 10212 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_103
timestamp 1604681595
transform 1 0 10580 0 1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11316 0 1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13524 0 1 8016
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_127
timestamp 1604681595
transform 1 0 12788 0 1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_144
timestamp 1604681595
transform 1 0 14352 0 1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15548 0 1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 15180 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_152
timestamp 1604681595
transform 1 0 15088 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_154
timestamp 1604681595
transform 1 0 15272 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_173
timestamp 1604681595
transform 1 0 17020 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_185
timestamp 1604681595
transform 1 0 18124 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_197
timestamp 1604681595
transform 1 0 19228 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 21896 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 20792 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_209
timestamp 1604681595
transform 1 0 20332 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_213
timestamp 1604681595
transform 1 0 20700 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_215
timestamp 1604681595
transform 1 0 20884 0 1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_39
timestamp 1604681595
transform 1 0 4692 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 6716 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_51
timestamp 1604681595
transform 1 0 5796 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1604681595
transform 1 0 6532 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_62
timestamp 1604681595
transform 1 0 6808 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_74
timestamp 1604681595
transform 1 0 7912 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_86
timestamp 1604681595
transform 1 0 9016 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_98
timestamp 1604681595
transform 1 0 10120 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 11040 0 -1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 12328 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_106
timestamp 1604681595
transform 1 0 10856 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_114
timestamp 1604681595
transform 1 0 11592 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_123
timestamp 1604681595
transform 1 0 12420 0 -1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13064 0 -1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_129
timestamp 1604681595
transform 1 0 12972 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_136
timestamp 1604681595
transform 1 0 13616 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 14720 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15916 0 -1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_152
timestamp 1604681595
transform 1 0 15088 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_160
timestamp 1604681595
transform 1 0 15824 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 18032 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 17940 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_170
timestamp 1604681595
transform 1 0 16744 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_182
timestamp 1604681595
transform 1 0 17848 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_187
timestamp 1604681595
transform 1 0 18308 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 19412 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_203
timestamp 1604681595
transform 1 0 19780 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 20516 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 21896 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 3956 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_32
timestamp 1604681595
transform 1 0 4048 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_39
timestamp 1604681595
transform 1 0 4692 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_44
timestamp 1604681595
transform 1 0 5152 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_56
timestamp 1604681595
transform 1 0 6256 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_51
timestamp 1604681595
transform 1 0 5796 0 -1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_59
timestamp 1604681595
transform 1 0 6532 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_62
timestamp 1604681595
transform 1 0 6808 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_68
timestamp 1604681595
transform 1 0 7360 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_80
timestamp 1604681595
transform 1 0 8464 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_74
timestamp 1604681595
transform 1 0 7912 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 9568 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1604681595
transform 1 0 9660 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_86
timestamp 1604681595
transform 1 0 9016 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_98
timestamp 1604681595
transform 1 0 10120 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 11500 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_105
timestamp 1604681595
transform 1 0 10764 0 1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_117
timestamp 1604681595
transform 1 0 11868 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_110
timestamp 1604681595
transform 1 0 11224 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_123
timestamp 1604681595
transform 1 0 12420 0 -1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 13064 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12972 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_13_129
timestamp 1604681595
transform 1 0 12972 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_134
timestamp 1604681595
transform 1 0 13432 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 15180 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_146
timestamp 1604681595
transform 1 0 14536 0 1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_152
timestamp 1604681595
transform 1 0 15088 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1604681595
transform 1 0 15824 0 1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_153
timestamp 1604681595
transform 1 0 15180 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_163
timestamp 1604681595
transform 1 0 16100 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16560 0 1 9104
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 -1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_175
timestamp 1604681595
transform 1 0 17204 0 -1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 19688 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_196
timestamp 1604681595
transform 1 0 19136 0 1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_206
timestamp 1604681595
transform 1 0 20056 0 1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_193
timestamp 1604681595
transform 1 0 18860 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_205
timestamp 1604681595
transform 1 0 19964 0 -1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 20516 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 21896 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 21896 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 20792 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1604681595
transform 1 0 20884 0 1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 3956 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1604681595
transform 1 0 3588 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_32
timestamp 1604681595
transform 1 0 4048 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1604681595
transform 1 0 5152 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_56
timestamp 1604681595
transform 1 0 6256 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_68
timestamp 1604681595
transform 1 0 7360 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_80
timestamp 1604681595
transform 1 0 8464 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 9568 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10396 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_93
timestamp 1604681595
transform 1 0 9660 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_104
timestamp 1604681595
transform 1 0 10672 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11868 0 1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_116
timestamp 1604681595
transform 1 0 11776 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604681595
transform 1 0 14168 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_133
timestamp 1604681595
transform 1 0 13340 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_141
timestamp 1604681595
transform 1 0 14076 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_145
timestamp 1604681595
transform 1 0 14444 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 15180 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_163
timestamp 1604681595
transform 1 0 16100 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17296 0 1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 19688 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_192
timestamp 1604681595
transform 1 0 18768 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1604681595
transform 1 0 19504 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_206
timestamp 1604681595
transform 1 0 20056 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 21896 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 20792 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_215
timestamp 1604681595
transform 1 0 20884 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604681595
transform 1 0 2484 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_39
timestamp 1604681595
transform 1 0 4692 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 6716 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_51
timestamp 1604681595
transform 1 0 5796 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1604681595
transform 1 0 6532 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_62
timestamp 1604681595
transform 1 0 6808 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_74
timestamp 1604681595
transform 1 0 7912 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_86
timestamp 1604681595
transform 1 0 9016 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_98
timestamp 1604681595
transform 1 0 10120 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12512 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 12328 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_110
timestamp 1604681595
transform 1 0 11224 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_123
timestamp 1604681595
transform 1 0 12420 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 14352 0 -1 11280
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 14076 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_133
timestamp 1604681595
transform 1 0 13340 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_160
timestamp 1604681595
transform 1 0 15824 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 16836 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 17940 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_168
timestamp 1604681595
transform 1 0 16560 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_175
timestamp 1604681595
transform 1 0 17204 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_193
timestamp 1604681595
transform 1 0 18860 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_205
timestamp 1604681595
transform 1 0 19964 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 20332 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 21896 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_213
timestamp 1604681595
transform 1 0 20700 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1604681595
transform 1 0 21436 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1604681595
transform 1 0 2484 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 3956 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1604681595
transform 1 0 3588 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_32
timestamp 1604681595
transform 1 0 4048 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_44
timestamp 1604681595
transform 1 0 5152 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_56
timestamp 1604681595
transform 1 0 6256 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_68
timestamp 1604681595
transform 1 0 7360 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_80
timestamp 1604681595
transform 1 0 8464 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 9568 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1604681595
transform 1 0 9660 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 12328 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_105
timestamp 1604681595
transform 1 0 10764 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1604681595
transform 1 0 11868 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1604681595
transform 1 0 12236 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_125
timestamp 1604681595
transform 1 0 12604 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1604681595
transform 1 0 13616 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_133
timestamp 1604681595
transform 1 0 13340 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_139
timestamp 1604681595
transform 1 0 13892 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 15180 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_151
timestamp 1604681595
transform 1 0 14996 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_163
timestamp 1604681595
transform 1 0 16100 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 16836 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17848 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_174
timestamp 1604681595
transform 1 0 17112 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_188
timestamp 1604681595
transform 1 0 18400 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_206
timestamp 1604681595
transform 1 0 20056 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 21896 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 20792 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_215
timestamp 1604681595
transform 1 0 20884 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604681595
transform 1 0 2484 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_39
timestamp 1604681595
transform 1 0 4692 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 6716 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_51
timestamp 1604681595
transform 1 0 5796 0 -1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_59
timestamp 1604681595
transform 1 0 6532 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_62
timestamp 1604681595
transform 1 0 6808 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1604681595
transform 1 0 7268 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8648 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_66
timestamp 1604681595
transform 1 0 7176 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_70
timestamp 1604681595
transform 1 0 7544 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_98
timestamp 1604681595
transform 1 0 10120 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12604 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 12328 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_110
timestamp 1604681595
transform 1 0 11224 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_123
timestamp 1604681595
transform 1 0 12420 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 14352 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_134
timestamp 1604681595
transform 1 0 13432 0 -1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_142
timestamp 1604681595
transform 1 0 14168 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15456 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_148
timestamp 1604681595
transform 1 0 14720 0 -1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 18308 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 17940 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_172
timestamp 1604681595
transform 1 0 16928 0 -1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_180
timestamp 1604681595
transform 1 0 17664 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_184
timestamp 1604681595
transform 1 0 18032 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 19412 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_191
timestamp 1604681595
transform 1 0 18676 0 -1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_203
timestamp 1604681595
transform 1 0 19780 0 -1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 20516 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 21896 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604681595
transform 1 0 2484 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 3956 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp 1604681595
transform 1 0 3588 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_32
timestamp 1604681595
transform 1 0 4048 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_39
timestamp 1604681595
transform 1 0 4692 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5980 0 1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 6716 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_44
timestamp 1604681595
transform 1 0 5152 0 1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_52
timestamp 1604681595
transform 1 0 5888 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_51
timestamp 1604681595
transform 1 0 5796 0 -1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_59
timestamp 1604681595
transform 1 0 6532 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_62
timestamp 1604681595
transform 1 0 6808 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6992 0 -1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1604681595
transform 1 0 7452 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_81
timestamp 1604681595
transform 1 0 8556 0 1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_73
timestamp 1604681595
transform 1 0 7820 0 -1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1604681595
transform 1 0 8556 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10120 0 -1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8832 0 -1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 9568 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_89
timestamp 1604681595
transform 1 0 9292 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1604681595
transform 1 0 9660 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_90
timestamp 1604681595
transform 1 0 9384 0 -1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11224 0 1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 -1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 12328 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_105
timestamp 1604681595
transform 1 0 10764 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_109
timestamp 1604681595
transform 1 0 11132 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_114
timestamp 1604681595
transform 1 0 11592 0 -1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13432 0 1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14352 0 -1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_126
timestamp 1604681595
transform 1 0 12696 0 1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_143
timestamp 1604681595
transform 1 0 14260 0 1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_132
timestamp 1604681595
transform 1 0 13248 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 15548 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16284 0 -1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 15180 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 16100 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_151
timestamp 1604681595
transform 1 0 14996 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_154
timestamp 1604681595
transform 1 0 15272 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_161
timestamp 1604681595
transform 1 0 15916 0 1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_150
timestamp 1604681595
transform 1 0 14904 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_162
timestamp 1604681595
transform 1 0 16008 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16652 0 1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 17940 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_185
timestamp 1604681595
transform 1 0 18124 0 1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_174
timestamp 1604681595
transform 1 0 17112 0 -1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_182
timestamp 1604681595
transform 1 0 17848 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_184
timestamp 1604681595
transform 1 0 18032 0 -1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18584 0 -1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18860 0 1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20148 0 -1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_202
timestamp 1604681595
transform 1 0 19688 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_199
timestamp 1604681595
transform 1 0 19412 0 -1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 21896 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 21896 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 20792 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_215
timestamp 1604681595
transform 1 0 20884 0 1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_213
timestamp 1604681595
transform 1 0 20700 0 -1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1604681595
transform 1 0 21436 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604681595
transform 1 0 2484 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 3956 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1604681595
transform 1 0 3588 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_32
timestamp 1604681595
transform 1 0 4048 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_44
timestamp 1604681595
transform 1 0 5152 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_56
timestamp 1604681595
transform 1 0 6256 0 1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6900 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_72
timestamp 1604681595
transform 1 0 7728 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10212 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 9568 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_84
timestamp 1604681595
transform 1 0 8832 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_93
timestamp 1604681595
transform 1 0 9660 0 1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 11776 0 1 13456
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_21_108
timestamp 1604681595
transform 1 0 11040 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_145
timestamp 1604681595
transform 1 0 14444 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15824 0 1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 15180 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_154
timestamp 1604681595
transform 1 0 15272 0 1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_166
timestamp 1604681595
transform 1 0 16376 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 17112 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18216 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_178
timestamp 1604681595
transform 1 0 17480 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 19780 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_195
timestamp 1604681595
transform 1 0 19044 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_206
timestamp 1604681595
transform 1 0 20056 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 21896 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 20792 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_215
timestamp 1604681595
transform 1 0 20884 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_39
timestamp 1604681595
transform 1 0 4692 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 6716 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_51
timestamp 1604681595
transform 1 0 5796 0 -1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_59
timestamp 1604681595
transform 1 0 6532 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_78
timestamp 1604681595
transform 1 0 8280 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9936 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_22_90
timestamp 1604681595
transform 1 0 9384 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 12328 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_112
timestamp 1604681595
transform 1 0 11408 0 -1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_120
timestamp 1604681595
transform 1 0 12144 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_139
timestamp 1604681595
transform 1 0 13892 0 -1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1604681595
transform 1 0 14720 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15732 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_147
timestamp 1604681595
transform 1 0 14628 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_151
timestamp 1604681595
transform 1 0 14996 0 -1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18032 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 17940 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_175
timestamp 1604681595
transform 1 0 17204 0 -1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_200
timestamp 1604681595
transform 1 0 19504 0 -1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_208
timestamp 1604681595
transform 1 0 20240 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 20516 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 21896 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_32
timestamp 1604681595
transform 1 0 4048 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_44
timestamp 1604681595
transform 1 0 5152 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_56
timestamp 1604681595
transform 1 0 6256 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7360 0 1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_84
timestamp 1604681595
transform 1 0 8832 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_102
timestamp 1604681595
transform 1 0 10488 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11224 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_119
timestamp 1604681595
transform 1 0 12052 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12788 0 1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_143
timestamp 1604681595
transform 1 0 14260 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_151
timestamp 1604681595
transform 1 0 14996 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_163
timestamp 1604681595
transform 1 0 16100 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 17296 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_175
timestamp 1604681595
transform 1 0 17204 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_180
timestamp 1604681595
transform 1 0 17664 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 18400 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_192
timestamp 1604681595
transform 1 0 18768 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_206
timestamp 1604681595
transform 1 0 20056 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 21896 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_215
timestamp 1604681595
transform 1 0 20884 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_39
timestamp 1604681595
transform 1 0 4692 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 -1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 6716 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_51
timestamp 1604681595
transform 1 0 5796 0 -1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_59
timestamp 1604681595
transform 1 0 6532 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8372 0 -1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_71
timestamp 1604681595
transform 1 0 7636 0 -1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 10580 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_95
timestamp 1604681595
transform 1 0 9844 0 -1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 12328 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 11592 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_106
timestamp 1604681595
transform 1 0 10856 0 -1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_117
timestamp 1604681595
transform 1 0 11868 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_121
timestamp 1604681595
transform 1 0 12236 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1604681595
transform 1 0 12420 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13892 0 -1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1604681595
transform 1 0 13524 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 15824 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_148
timestamp 1604681595
transform 1 0 14720 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_163
timestamp 1604681595
transform 1 0 16100 0 -1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 16836 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18216 0 -1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 17940 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_175
timestamp 1604681595
transform 1 0 17204 0 -1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_184
timestamp 1604681595
transform 1 0 18032 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19964 0 -1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_195
timestamp 1604681595
transform 1 0 19044 0 -1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_203
timestamp 1604681595
transform 1 0 19780 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 21896 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_211
timestamp 1604681595
transform 1 0 20516 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 3956 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_32
timestamp 1604681595
transform 1 0 4048 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5704 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_25_44
timestamp 1604681595
transform 1 0 5152 0 1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_66
timestamp 1604681595
transform 1 0 7176 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_78
timestamp 1604681595
transform 1 0 8280 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10120 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 9568 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_90
timestamp 1604681595
transform 1 0 9384 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_93
timestamp 1604681595
transform 1 0 9660 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_97
timestamp 1604681595
transform 1 0 10028 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_107
timestamp 1604681595
transform 1 0 10948 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_119
timestamp 1604681595
transform 1 0 12052 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12788 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_136
timestamp 1604681595
transform 1 0 13616 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15548 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 15180 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_148
timestamp 1604681595
transform 1 0 14720 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_152
timestamp 1604681595
transform 1 0 15088 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_154
timestamp 1604681595
transform 1 0 15272 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_166
timestamp 1604681595
transform 1 0 16376 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17296 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_174
timestamp 1604681595
transform 1 0 17112 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_192
timestamp 1604681595
transform 1 0 18768 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_206
timestamp 1604681595
transform 1 0 20056 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 21896 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 20792 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_215
timestamp 1604681595
transform 1 0 20884 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 3956 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_39
timestamp 1604681595
transform 1 0 4692 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1604681595
transform 1 0 4048 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6256 0 1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 6716 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_51
timestamp 1604681595
transform 1 0 5796 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_59
timestamp 1604681595
transform 1 0 6532 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_62
timestamp 1604681595
transform 1 0 6808 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1604681595
transform 1 0 5152 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1604681595
transform 1 0 7360 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_71
timestamp 1604681595
transform 1 0 7636 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1604681595
transform 1 0 8740 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_72
timestamp 1604681595
transform 1 0 7728 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9108 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10488 0 1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 9568 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 8832 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_103
timestamp 1604681595
transform 1 0 10580 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_84
timestamp 1604681595
transform 1 0 8832 0 1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_93
timestamp 1604681595
transform 1 0 9660 0 1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_101
timestamp 1604681595
transform 1 0 10396 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604681595
transform 1 0 11316 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 12328 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_114
timestamp 1604681595
transform 1 0 11592 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_118
timestamp 1604681595
transform 1 0 11960 0 1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12972 0 1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 12696 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_139
timestamp 1604681595
transform 1 0 13892 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_145
timestamp 1604681595
transform 1 0 14444 0 1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 14628 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15732 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 15180 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_151
timestamp 1604681595
transform 1 0 14996 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 17940 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_175
timestamp 1604681595
transform 1 0 17204 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_170
timestamp 1604681595
transform 1 0 16744 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_182
timestamp 1604681595
transform 1 0 17848 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 18400 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19872 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_193
timestamp 1604681595
transform 1 0 18860 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_201
timestamp 1604681595
transform 1 0 19596 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_192
timestamp 1604681595
transform 1 0 18768 0 1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_206
timestamp 1604681595
transform 1 0 20056 0 1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 21896 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 21896 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 20792 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_210
timestamp 1604681595
transform 1 0 20424 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_222
timestamp 1604681595
transform 1 0 21528 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_215
timestamp 1604681595
transform 1 0 20884 0 1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_39
timestamp 1604681595
transform 1 0 4692 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 6716 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_51
timestamp 1604681595
transform 1 0 5796 0 -1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_59
timestamp 1604681595
transform 1 0 6532 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_62
timestamp 1604681595
transform 1 0 6808 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_72
timestamp 1604681595
transform 1 0 7728 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9200 0 -1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1604681595
transform 1 0 10028 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 11316 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 -1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 12328 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_109
timestamp 1604681595
transform 1 0 11132 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_114
timestamp 1604681595
transform 1 0 11592 0 -1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_132
timestamp 1604681595
transform 1 0 13248 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_144
timestamp 1604681595
transform 1 0 14352 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14536 0 -1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_155
timestamp 1604681595
transform 1 0 15364 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 16836 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18124 0 -1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 17940 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_167
timestamp 1604681595
transform 1 0 16468 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_175
timestamp 1604681595
transform 1 0 17204 0 -1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_184
timestamp 1604681595
transform 1 0 18032 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19872 0 -1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_194
timestamp 1604681595
transform 1 0 18952 0 -1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 21896 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_210
timestamp 1604681595
transform 1 0 20424 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_222
timestamp 1604681595
transform 1 0 21528 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 3956 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1604681595
transform 1 0 4048 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5520 0 1 17808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_44
timestamp 1604681595
transform 1 0 5152 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7728 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_64
timestamp 1604681595
transform 1 0 6992 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_81
timestamp 1604681595
transform 1 0 8556 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1604681595
transform 1 0 9844 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 9568 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_89
timestamp 1604681595
transform 1 0 9292 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_93
timestamp 1604681595
transform 1 0 9660 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1604681595
transform 1 0 10856 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 11868 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_109
timestamp 1604681595
transform 1 0 11132 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_121
timestamp 1604681595
transform 1 0 12236 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 12972 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 14076 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_133
timestamp 1604681595
transform 1 0 13340 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_145
timestamp 1604681595
transform 1 0 14444 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 16100 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 15180 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_154
timestamp 1604681595
transform 1 0 15272 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_162
timestamp 1604681595
transform 1 0 16008 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17204 0 1 17808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_29_167
timestamp 1604681595
transform 1 0 16468 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 19688 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_191
timestamp 1604681595
transform 1 0 18676 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_199
timestamp 1604681595
transform 1 0 19412 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_206
timestamp 1604681595
transform 1 0 20056 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 21896 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 20792 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_215
timestamp 1604681595
transform 1 0 20884 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_39
timestamp 1604681595
transform 1 0 4692 0 -1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 6716 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_51
timestamp 1604681595
transform 1 0 5796 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_59
timestamp 1604681595
transform 1 0 6532 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_62
timestamp 1604681595
transform 1 0 6808 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6992 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8556 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_73
timestamp 1604681595
transform 1 0 7820 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10120 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_90
timestamp 1604681595
transform 1 0 9384 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 12328 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_107
timestamp 1604681595
transform 1 0 10948 0 -1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_119
timestamp 1604681595
transform 1 0 12052 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_132
timestamp 1604681595
transform 1 0 13248 0 -1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_144
timestamp 1604681595
transform 1 0 14352 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604681595
transform 1 0 14628 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15732 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_151
timestamp 1604681595
transform 1 0 14996 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 17940 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_175
timestamp 1604681595
transform 1 0 17204 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19872 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_193
timestamp 1604681595
transform 1 0 18860 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_201
timestamp 1604681595
transform 1 0 19596 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 21896 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_210
timestamp 1604681595
transform 1 0 20424 0 -1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_222
timestamp 1604681595
transform 1 0 21528 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 3956 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_32
timestamp 1604681595
transform 1 0 4048 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1604681595
transform 1 0 6348 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_44
timestamp 1604681595
transform 1 0 5152 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_56
timestamp 1604681595
transform 1 0 6256 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_60
timestamp 1604681595
transform 1 0 6624 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7360 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 9568 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_84
timestamp 1604681595
transform 1 0 8832 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11868 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_109
timestamp 1604681595
transform 1 0 11132 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 14076 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_133
timestamp 1604681595
transform 1 0 13340 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_145
timestamp 1604681595
transform 1 0 14444 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 15180 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 17756 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_170
timestamp 1604681595
transform 1 0 16744 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_178
timestamp 1604681595
transform 1 0 17480 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_185
timestamp 1604681595
transform 1 0 18124 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18860 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_199
timestamp 1604681595
transform 1 0 19412 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 21896 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 20792 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_211
timestamp 1604681595
transform 1 0 20516 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_215
timestamp 1604681595
transform 1 0 20884 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_39
timestamp 1604681595
transform 1 0 4692 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6808 0 -1 19984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_51
timestamp 1604681595
transform 1 0 5796 0 -1 19984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_59
timestamp 1604681595
transform 1 0 6532 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_78
timestamp 1604681595
transform 1 0 8280 0 -1 19984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9108 0 -1 19984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_32_86
timestamp 1604681595
transform 1 0 9016 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_103
timestamp 1604681595
transform 1 0 10580 0 -1 19984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1604681595
transform 1 0 11316 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_114
timestamp 1604681595
transform 1 0 11592 0 -1 19984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_123
timestamp 1604681595
transform 1 0 12420 0 -1 19984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13340 0 -1 19984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_131
timestamp 1604681595
transform 1 0 13156 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15548 0 -1 19984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_149
timestamp 1604681595
transform 1 0 14812 0 -1 19984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1604681595
transform 1 0 16376 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_178
timestamp 1604681595
transform 1 0 17480 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_182
timestamp 1604681595
transform 1 0 17848 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19780 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1604681595
transform 1 0 18584 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_202
timestamp 1604681595
transform 1 0 19688 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 21896 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1604681595
transform 1 0 20332 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1604681595
transform 1 0 21436 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 3956 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_32
timestamp 1604681595
transform 1 0 4048 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 6808 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_44
timestamp 1604681595
transform 1 0 5152 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_56
timestamp 1604681595
transform 1 0 6256 0 1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7176 0 1 19984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_33_63
timestamp 1604681595
transform 1 0 6900 0 1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_75
timestamp 1604681595
transform 1 0 8004 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1604681595
transform 1 0 10396 0 1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9660 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_87
timestamp 1604681595
transform 1 0 9108 0 1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_94
timestamp 1604681595
transform 1 0 9752 0 1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_100
timestamp 1604681595
transform 1 0 10304 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_104
timestamp 1604681595
transform 1 0 10672 0 1 19984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 11408 0 1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12512 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_116
timestamp 1604681595
transform 1 0 11776 0 1 19984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_125
timestamp 1604681595
transform 1 0 12604 0 1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12972 0 1 19984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_33_138
timestamp 1604681595
transform 1 0 13800 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16008 0 1 19984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 15364 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_150
timestamp 1604681595
transform 1 0 14904 0 1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_154
timestamp 1604681595
transform 1 0 15272 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_156
timestamp 1604681595
transform 1 0 15456 0 1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18308 0 1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 18216 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_171
timestamp 1604681595
transform 1 0 16836 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_183
timestamp 1604681595
transform 1 0 17940 0 1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 19964 0 1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1604681595
transform 1 0 18860 0 1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 21896 0 1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 21068 0 1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_209
timestamp 1604681595
transform 1 0 20332 0 1 19984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1604681595
transform 1 0 21160 0 1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1604681595
transform 1 0 21528 0 1 19984
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 5576 480 5696 6 ccff_head
port 0 nsew default input
rlabel metal3 s 0 17000 480 17120 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 22520 2856 23000 2976 6 chanx_right_in[0]
port 2 nsew default input
rlabel metal3 s 22520 7752 23000 7872 6 chanx_right_in[10]
port 3 nsew default input
rlabel metal3 s 22520 8296 23000 8416 6 chanx_right_in[11]
port 4 nsew default input
rlabel metal3 s 22520 8704 23000 8824 6 chanx_right_in[12]
port 5 nsew default input
rlabel metal3 s 22520 9248 23000 9368 6 chanx_right_in[13]
port 6 nsew default input
rlabel metal3 s 22520 9656 23000 9776 6 chanx_right_in[14]
port 7 nsew default input
rlabel metal3 s 22520 10200 23000 10320 6 chanx_right_in[15]
port 8 nsew default input
rlabel metal3 s 22520 10744 23000 10864 6 chanx_right_in[16]
port 9 nsew default input
rlabel metal3 s 22520 11152 23000 11272 6 chanx_right_in[17]
port 10 nsew default input
rlabel metal3 s 22520 11696 23000 11816 6 chanx_right_in[18]
port 11 nsew default input
rlabel metal3 s 22520 12104 23000 12224 6 chanx_right_in[19]
port 12 nsew default input
rlabel metal3 s 22520 3400 23000 3520 6 chanx_right_in[1]
port 13 nsew default input
rlabel metal3 s 22520 3808 23000 3928 6 chanx_right_in[2]
port 14 nsew default input
rlabel metal3 s 22520 4352 23000 4472 6 chanx_right_in[3]
port 15 nsew default input
rlabel metal3 s 22520 4760 23000 4880 6 chanx_right_in[4]
port 16 nsew default input
rlabel metal3 s 22520 5304 23000 5424 6 chanx_right_in[5]
port 17 nsew default input
rlabel metal3 s 22520 5848 23000 5968 6 chanx_right_in[6]
port 18 nsew default input
rlabel metal3 s 22520 6256 23000 6376 6 chanx_right_in[7]
port 19 nsew default input
rlabel metal3 s 22520 6800 23000 6920 6 chanx_right_in[8]
port 20 nsew default input
rlabel metal3 s 22520 7208 23000 7328 6 chanx_right_in[9]
port 21 nsew default input
rlabel metal3 s 22520 12648 23000 12768 6 chanx_right_out[0]
port 22 nsew default tristate
rlabel metal3 s 22520 17544 23000 17664 6 chanx_right_out[10]
port 23 nsew default tristate
rlabel metal3 s 22520 18088 23000 18208 6 chanx_right_out[11]
port 24 nsew default tristate
rlabel metal3 s 22520 18496 23000 18616 6 chanx_right_out[12]
port 25 nsew default tristate
rlabel metal3 s 22520 19040 23000 19160 6 chanx_right_out[13]
port 26 nsew default tristate
rlabel metal3 s 22520 19448 23000 19568 6 chanx_right_out[14]
port 27 nsew default tristate
rlabel metal3 s 22520 19992 23000 20112 6 chanx_right_out[15]
port 28 nsew default tristate
rlabel metal3 s 22520 20536 23000 20656 6 chanx_right_out[16]
port 29 nsew default tristate
rlabel metal3 s 22520 20944 23000 21064 6 chanx_right_out[17]
port 30 nsew default tristate
rlabel metal3 s 22520 21488 23000 21608 6 chanx_right_out[18]
port 31 nsew default tristate
rlabel metal3 s 22520 21896 23000 22016 6 chanx_right_out[19]
port 32 nsew default tristate
rlabel metal3 s 22520 13192 23000 13312 6 chanx_right_out[1]
port 33 nsew default tristate
rlabel metal3 s 22520 13600 23000 13720 6 chanx_right_out[2]
port 34 nsew default tristate
rlabel metal3 s 22520 14144 23000 14264 6 chanx_right_out[3]
port 35 nsew default tristate
rlabel metal3 s 22520 14552 23000 14672 6 chanx_right_out[4]
port 36 nsew default tristate
rlabel metal3 s 22520 15096 23000 15216 6 chanx_right_out[5]
port 37 nsew default tristate
rlabel metal3 s 22520 15640 23000 15760 6 chanx_right_out[6]
port 38 nsew default tristate
rlabel metal3 s 22520 16048 23000 16168 6 chanx_right_out[7]
port 39 nsew default tristate
rlabel metal3 s 22520 16592 23000 16712 6 chanx_right_out[8]
port 40 nsew default tristate
rlabel metal3 s 22520 17000 23000 17120 6 chanx_right_out[9]
port 41 nsew default tristate
rlabel metal2 s 846 22376 902 22856 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 6458 22376 6514 22856 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 7010 22376 7066 22856 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 7562 22376 7618 22856 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 8114 22376 8170 22856 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 8666 22376 8722 22856 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 9218 22376 9274 22856 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 9770 22376 9826 22856 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 10322 22376 10378 22856 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 10874 22376 10930 22856 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 11426 22376 11482 22856 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 1398 22376 1454 22856 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 1950 22376 2006 22856 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 2502 22376 2558 22856 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 3054 22376 3110 22856 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 3606 22376 3662 22856 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 4158 22376 4214 22856 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 4710 22376 4766 22856 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 5262 22376 5318 22856 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 5814 22376 5870 22856 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 12070 22376 12126 22856 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 17682 22376 17738 22856 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 18234 22376 18290 22856 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 18786 22376 18842 22856 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 19338 22376 19394 22856 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 19890 22376 19946 22856 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 20442 22376 20498 22856 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 20994 22376 21050 22856 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 21546 22376 21602 22856 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 22098 22376 22154 22856 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 22650 22376 22706 22856 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 12622 22376 12678 22856 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 13174 22376 13230 22856 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 13726 22376 13782 22856 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 14278 22376 14334 22856 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 14830 22376 14886 22856 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 15382 22376 15438 22856 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 15934 22376 15990 22856 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 16486 22376 16542 22856 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 17038 22376 17094 22856 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 22520 22440 23000 22560 6 prog_clk
port 82 nsew default input
rlabel metal3 s 22520 2312 23000 2432 6 right_bottom_grid_pin_11_
port 83 nsew default input
rlabel metal3 s 22520 0 23000 120 6 right_bottom_grid_pin_1_
port 84 nsew default input
rlabel metal3 s 22520 408 23000 528 6 right_bottom_grid_pin_3_
port 85 nsew default input
rlabel metal3 s 22520 952 23000 1072 6 right_bottom_grid_pin_5_
port 86 nsew default input
rlabel metal3 s 22520 1360 23000 1480 6 right_bottom_grid_pin_7_
port 87 nsew default input
rlabel metal3 s 22520 1904 23000 2024 6 right_bottom_grid_pin_9_
port 88 nsew default input
rlabel metal2 s 294 22376 350 22856 6 top_left_grid_pin_1_
port 89 nsew default input
rlabel metal4 s 4409 1984 4729 20576 6 VPWR
port 90 nsew default input
rlabel metal4 s 7875 1984 8195 20576 6 VGND
port 91 nsew default input
<< properties >>
string FIXED_BBOX 0 0 23000 22856
<< end >>
