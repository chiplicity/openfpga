* NGSPICE file created from grid_clb.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfxtp_1 abstract view
.subckt sky130_fd_sc_hd__sdfxtp_1 D Q SCD SCE CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt grid_clb SC_IN_BOT SC_IN_TOP SC_OUT_BOT SC_OUT_TOP Test_en bottom_width_0_height_0__pin_50_
+ bottom_width_0_height_0__pin_51_ ccff_head ccff_tail clk left_width_0_height_0__pin_52_
+ prog_clk right_width_0_height_0__pin_16_ right_width_0_height_0__pin_17_ right_width_0_height_0__pin_18_
+ right_width_0_height_0__pin_19_ right_width_0_height_0__pin_20_ right_width_0_height_0__pin_21_
+ right_width_0_height_0__pin_22_ right_width_0_height_0__pin_23_ right_width_0_height_0__pin_24_
+ right_width_0_height_0__pin_25_ right_width_0_height_0__pin_26_ right_width_0_height_0__pin_27_
+ right_width_0_height_0__pin_28_ right_width_0_height_0__pin_29_ right_width_0_height_0__pin_30_
+ right_width_0_height_0__pin_31_ right_width_0_height_0__pin_42_lower right_width_0_height_0__pin_42_upper
+ right_width_0_height_0__pin_43_lower right_width_0_height_0__pin_43_upper right_width_0_height_0__pin_44_lower
+ right_width_0_height_0__pin_44_upper right_width_0_height_0__pin_45_lower right_width_0_height_0__pin_45_upper
+ right_width_0_height_0__pin_46_lower right_width_0_height_0__pin_46_upper right_width_0_height_0__pin_47_lower
+ right_width_0_height_0__pin_47_upper right_width_0_height_0__pin_48_lower right_width_0_height_0__pin_48_upper
+ right_width_0_height_0__pin_49_lower right_width_0_height_0__pin_49_upper top_width_0_height_0__pin_0_
+ top_width_0_height_0__pin_10_ top_width_0_height_0__pin_11_ top_width_0_height_0__pin_12_
+ top_width_0_height_0__pin_13_ top_width_0_height_0__pin_14_ top_width_0_height_0__pin_15_
+ top_width_0_height_0__pin_1_ top_width_0_height_0__pin_2_ top_width_0_height_0__pin_32_
+ top_width_0_height_0__pin_33_ top_width_0_height_0__pin_34_lower top_width_0_height_0__pin_34_upper
+ top_width_0_height_0__pin_35_lower top_width_0_height_0__pin_35_upper top_width_0_height_0__pin_36_lower
+ top_width_0_height_0__pin_36_upper top_width_0_height_0__pin_37_lower top_width_0_height_0__pin_37_upper
+ top_width_0_height_0__pin_38_lower top_width_0_height_0__pin_38_upper top_width_0_height_0__pin_39_lower
+ top_width_0_height_0__pin_39_upper top_width_0_height_0__pin_3_ top_width_0_height_0__pin_40_lower
+ top_width_0_height_0__pin_40_upper top_width_0_height_0__pin_41_lower top_width_0_height_0__pin_41_upper
+ top_width_0_height_0__pin_4_ top_width_0_height_0__pin_5_ top_width_0_height_0__pin_6_
+ top_width_0_height_0__pin_7_ top_width_0_height_0__pin_8_ top_width_0_height_0__pin_9_
+ VPWR VGND
X_83_ top_width_0_height_0__pin_41_lower top_width_0_height_0__pin_41_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _49_/HI ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_48_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_66_ SC_OUT_BOT SC_OUT_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ top_width_0_height_0__pin_1_ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_49_ _49_/HI _49_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xclkbuf_3_4_0_prog_clk clkbuf_2_2_0_prog_clk/X clkbuf_4_9_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ccff_head ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ right_width_0_height_0__pin_22_ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_82_ top_width_0_height_0__pin_40_lower top_width_0_height_0__pin_40_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_65_ SC_IN_BOT SC_IN_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ top_width_0_height_0__pin_0_ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xclkbuf_4_6_0_prog_clk clkbuf_4_7_0_prog_clk/A clkbuf_4_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ SC_OUT_BOT ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_48_ _48_/HI _48_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_81_ top_width_0_height_0__pin_39_lower top_width_0_height_0__pin_39_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ right_width_0_height_0__pin_21_ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_64_ _64_/HI bottom_width_0_height_0__pin_51_ VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_47_ _47_/HI _47_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_1_0_prog_clk clkbuf_1_0_0_prog_clk/X clkbuf_3_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_80_ top_width_0_height_0__pin_38_lower top_width_0_height_0__pin_38_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ right_width_0_height_0__pin_20_ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_63_ _63_/HI _63_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
X_46_ _46_/HI _46_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_3_3_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_4_7_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _32_/HI ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ top_width_0_height_0__pin_41_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_62_ _62_/HI _62_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_5_0_prog_clk clkbuf_4_5_0_prog_clk/A clkbuf_4_5_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_45_ _45_/HI _45_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ Test_en clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _61_/HI ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ top_width_0_height_0__pin_38_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_61_ _61_/HI _61_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_5_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_44_ _44_/HI _44_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _39_/HI ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XFILLER_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ top_width_0_height_0__pin_3_ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_60_ _60_/HI _60_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0_0_prog_clk clkbuf_1_0_0_prog_clk/X clkbuf_2_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_43_ _43_/HI _43_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_4_5_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ Test_en clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ top_width_0_height_0__pin_10_ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_42_ _42_/HI _42_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_4_0_prog_clk clkbuf_4_5_0_prog_clk/A clkbuf_4_4_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ right_width_0_height_0__pin_23_ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _51_/HI ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_21_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ top_width_0_height_0__pin_9_ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _50_/HI ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ccff_tail ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_17_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_41_ _41_/HI _41_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ right_width_0_height_0__pin_30_ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ top_width_0_height_0__pin_8_ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ Test_en clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_40_ _40_/HI _40_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ right_width_0_height_0__pin_29_ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _36_/HI ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_43_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_prog_clk clkbuf_2_0_0_prog_clk/X clkbuf_4_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ right_width_0_height_0__pin_28_ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_3_0_prog_clk clkbuf_4_3_0_prog_clk/A clkbuf_4_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _33_/HI ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ top_width_0_height_0__pin_40_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _46_/HI ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ SC_OUT_BOT ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XFILLER_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_0_0_prog_clk clkbuf_2_0_0_prog_clk/X clkbuf_4_1_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _63_/HI ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_79_ top_width_0_height_0__pin_37_lower top_width_0_height_0__pin_37_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ top_width_0_height_0__pin_11_ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_2_0_prog_clk clkbuf_4_3_0_prog_clk/A clkbuf_4_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_78_ top_width_0_height_0__pin_36_lower top_width_0_height_0__pin_36_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
Xclkbuf_4_15_0_prog_clk clkbuf_3_7_0_prog_clk/X clkbuf_4_15_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ right_width_0_height_0__pin_18_ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _42_/HI ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_77_ top_width_0_height_0__pin_35_lower top_width_0_height_0__pin_35_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ccff_tail clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ right_width_0_height_0__pin_31_ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_21_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ right_width_0_height_0__pin_17_ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _40_/HI ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_45_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_76_ top_width_0_height_0__pin_34_lower top_width_0_height_0__pin_34_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_59_ _59_/HI _59_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ right_width_0_height_0__pin_16_ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _37_/HI ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_42_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_1_0_prog_clk clkbuf_4_1_0_prog_clk/A clkbuf_4_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
X_75_ right_width_0_height_0__pin_49_lower right_width_0_height_0__pin_49_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_58_ _58_/HI _58_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_16_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_4_14_0_prog_clk clkbuf_3_7_0_prog_clk/X clkbuf_4_14_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ Test_en clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_74_ right_width_0_height_0__pin_48_lower right_width_0_height_0__pin_48_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_clk clkbuf_0_clk/X clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_57_ _57_/HI _57_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _38_/HI ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _43_/HI ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_73_ right_width_0_height_0__pin_47_lower right_width_0_height_0__pin_47_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_56_ _56_/HI _56_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_39_ _39_/HI _39_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_clk clkbuf_0_clk/X clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_72_ right_width_0_height_0__pin_46_lower right_width_0_height_0__pin_46_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ Test_en clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_55_ _55_/HI _55_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_0_0_prog_clk clkbuf_4_1_0_prog_clk/A clkbuf_4_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _52_/HI ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ top_width_0_height_0__pin_35_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_38_ _38_/HI _38_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_22_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ top_width_0_height_0__pin_6_ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_13_0_prog_clk clkbuf_3_6_0_prog_clk/X clkbuf_4_13_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__clkbuf_1
X_71_ right_width_0_height_0__pin_45_lower right_width_0_height_0__pin_45_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _55_/HI ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_54_ _54_/HI _54_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ right_width_0_height_0__pin_19_ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_37_ _37_/HI _37_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ top_width_0_height_0__pin_5_ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _44_/HI ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_47_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_70_ right_width_0_height_0__pin_44_lower right_width_0_height_0__pin_44_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_53_ _53_/HI _53_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _34_/HI ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ right_width_0_height_0__pin_26_ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_36_ _36_/HI _36_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ top_width_0_height_0__pin_4_ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _41_/HI ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_44_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_52_ _52_/HI _52_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ right_width_0_height_0__pin_25_ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_35_ _35_/HI _35_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_30_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xclkbuf_4_12_0_prog_clk clkbuf_3_6_0_prog_clk/X clkbuf_4_12_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_51_ _51_/HI _51_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ right_width_0_height_0__pin_24_ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_34_ _34_/HI _34_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_50_ _50_/HI _50_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
X_33_ _33_/HI _33_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _62_/HI ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_3_7_0_prog_clk clkbuf_3_7_0_prog_clk/A clkbuf_3_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_32_ _32_/HI _32_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _56_/HI ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ top_width_0_height_0__pin_37_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_9_0_prog_clk clkbuf_4_9_0_prog_clk/A clkbuf_4_9_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _35_/HI ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_14_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ top_width_0_height_0__pin_7_ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_11_0_prog_clk clkbuf_3_5_0_prog_clk/X clkbuf_4_11_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _53_/HI ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ top_width_0_height_0__pin_34_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _48_/HI ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_49_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ top_width_0_height_0__pin_14_ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ Test_en clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ right_width_0_height_0__pin_27_ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_15_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _45_/HI ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_46_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_6_0_prog_clk clkbuf_3_7_0_prog_clk/A clkbuf_3_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ top_width_0_height_0__pin_13_ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _58_/HI ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_prog_clk clkbuf_4_9_0_prog_clk/A clkbuf_4_8_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ top_width_0_height_0__pin_12_ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_10_0_prog_clk clkbuf_3_5_0_prog_clk/X clkbuf_4_10_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_0 _34_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ Test_en clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_22_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_3_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_3_7_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_1 _34_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_prog_clk clkbuf_2_2_0_prog_clk/X clkbuf_3_5_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_69_ right_width_0_height_0__pin_43_lower right_width_0_height_0__pin_43_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _47_/HI ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _60_/HI ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ top_width_0_height_0__pin_39_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_2 _50_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_4_7_0_prog_clk clkbuf_4_7_0_prog_clk/A clkbuf_4_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _54_/HI ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ SC_IN_BOT Test_en clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_68_ right_width_0_height_0__pin_42_lower right_width_0_height_0__pin_42_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _57_/HI ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ top_width_0_height_0__pin_36_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_3 _50_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_1_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ top_width_0_height_0__pin_2_ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ top_width_0_height_0__pin_32_ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_67_ SC_OUT_BOT bottom_width_0_height_0__pin_50_ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_28_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_28_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_2_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_2_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _59_/HI ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ top_width_0_height_0__pin_15_ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
.ends

