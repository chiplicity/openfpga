* NGSPICE file created from grid_clb.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfxtp_1 abstract view
.subckt sky130_fd_sc_hd__sdfxtp_1 D Q SCD SCE CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

.subckt grid_clb SC_IN_BOT SC_IN_TOP SC_OUT_BOT SC_OUT_TOP Test_en bottom_width_0_height_0__pin_50_
+ bottom_width_0_height_0__pin_51_ ccff_head ccff_tail clk left_width_0_height_0__pin_52_
+ prog_clk right_width_0_height_0__pin_16_ right_width_0_height_0__pin_17_ right_width_0_height_0__pin_18_
+ right_width_0_height_0__pin_19_ right_width_0_height_0__pin_20_ right_width_0_height_0__pin_21_
+ right_width_0_height_0__pin_22_ right_width_0_height_0__pin_23_ right_width_0_height_0__pin_24_
+ right_width_0_height_0__pin_25_ right_width_0_height_0__pin_26_ right_width_0_height_0__pin_27_
+ right_width_0_height_0__pin_28_ right_width_0_height_0__pin_29_ right_width_0_height_0__pin_30_
+ right_width_0_height_0__pin_31_ right_width_0_height_0__pin_42_lower right_width_0_height_0__pin_42_upper
+ right_width_0_height_0__pin_43_lower right_width_0_height_0__pin_43_upper right_width_0_height_0__pin_44_lower
+ right_width_0_height_0__pin_44_upper right_width_0_height_0__pin_45_lower right_width_0_height_0__pin_45_upper
+ right_width_0_height_0__pin_46_lower right_width_0_height_0__pin_46_upper right_width_0_height_0__pin_47_lower
+ right_width_0_height_0__pin_47_upper right_width_0_height_0__pin_48_lower right_width_0_height_0__pin_48_upper
+ right_width_0_height_0__pin_49_lower right_width_0_height_0__pin_49_upper top_width_0_height_0__pin_0_
+ top_width_0_height_0__pin_10_ top_width_0_height_0__pin_11_ top_width_0_height_0__pin_12_
+ top_width_0_height_0__pin_13_ top_width_0_height_0__pin_14_ top_width_0_height_0__pin_15_
+ top_width_0_height_0__pin_1_ top_width_0_height_0__pin_2_ top_width_0_height_0__pin_32_
+ top_width_0_height_0__pin_33_ top_width_0_height_0__pin_34_lower top_width_0_height_0__pin_34_upper
+ top_width_0_height_0__pin_35_lower top_width_0_height_0__pin_35_upper top_width_0_height_0__pin_36_lower
+ top_width_0_height_0__pin_36_upper top_width_0_height_0__pin_37_lower top_width_0_height_0__pin_37_upper
+ top_width_0_height_0__pin_38_lower top_width_0_height_0__pin_38_upper top_width_0_height_0__pin_39_lower
+ top_width_0_height_0__pin_39_upper top_width_0_height_0__pin_3_ top_width_0_height_0__pin_40_lower
+ top_width_0_height_0__pin_40_upper top_width_0_height_0__pin_41_lower top_width_0_height_0__pin_41_upper
+ top_width_0_height_0__pin_4_ top_width_0_height_0__pin_5_ top_width_0_height_0__pin_6_
+ top_width_0_height_0__pin_7_ top_width_0_height_0__pin_8_ top_width_0_height_0__pin_9_
+ VPWR VGND
XFILLER_27_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_83_ top_width_0_height_0__pin_41_lower top_width_0_height_0__pin_41_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _49_/HI ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_48_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_50_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_66_ SC_OUT_BOT bottom_width_0_height_0__pin_50_ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ top_width_0_height_0__pin_1_ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_15_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1_0_prog_clk_A clkbuf_2_1_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_49_ _49_/HI _49_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xclkbuf_3_4_0_prog_clk clkbuf_2_2_0_prog_clk/X clkbuf_4_9_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ccff_head ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _45_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ right_width_0_height_0__pin_22_ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_82_ top_width_0_height_0__pin_40_lower top_width_0_height_0__pin_40_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_prog_clk clkbuf_4_7_0_prog_clk/A clkbuf_4_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_52_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ top_width_0_height_0__pin_0_ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_65_ SC_OUT_BOT SC_OUT_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ SC_OUT_BOT ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_48_ _48_/HI _48_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_60_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_81_ top_width_0_height_0__pin_39_lower top_width_0_height_0__pin_39_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ right_width_0_height_0__pin_21_ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_44_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_50_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_42_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _37_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_64_ SC_IN_BOT SC_IN_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_64_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_47_ _47_/HI _47_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_1_0_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_62_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_1_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_80_ top_width_0_height_0__pin_38_lower top_width_0_height_0__pin_38_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ right_width_0_height_0__pin_20_ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_51_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_50_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_63_ _63_/HI _63_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_32_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_4_0_prog_clk_A clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XFILLER_37_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_46_ _46_/HI _46_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _61_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_50_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_3_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_4_7_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _32_/HI ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ top_width_0_height_0__pin_41_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_4_9_0_prog_clk_A clkbuf_4_9_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_62_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_53_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ right_width_0_height_0__pin_27_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_50_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_62_ _62_/HI _62_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_45_ _45_/HI _45_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_prog_clk clkbuf_3_2_0_prog_clk/X clkbuf_4_5_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_28_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
+ ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _53_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_clk_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ Test_en clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _61_/HI ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ top_width_0_height_0__pin_38_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_53_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_61_ _61_/HI _61_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_44_ _44_/HI _44_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_64_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _39_/HI ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_3_0_prog_clk_A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ right_width_0_height_0__pin_29_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XFILLER_3_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ top_width_0_height_0__pin_3_ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_13_0_prog_clk_A clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_26_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_0_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_3_1_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_60_ _60_/HI _60_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ right_width_0_height_0__pin_24_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _43_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_43_ _43_/HI _43_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ top_width_0_height_0__pin_15_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_42_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_2_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ Test_en clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_35_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ top_width_0_height_0__pin_10_ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_41_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_49_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_49_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_42_ _42_/HI _42_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ right_width_0_height_0__pin_22_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_2_0_prog_clk_A clkbuf_2_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_4_0_prog_clk clkbuf_3_2_0_prog_clk/X clkbuf_4_4_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ right_width_0_height_0__pin_23_ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XFILLER_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _51_/HI ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_47_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_23_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ right_width_0_height_0__pin_17_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ top_width_0_height_0__pin_9_ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _50_/HI ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ccff_tail ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_41_ _41_/HI _41_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__64__A SC_IN_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_42_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ top_width_0_height_0__pin_12_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ right_width_0_height_0__pin_30_ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ top_width_0_height_0__pin_3_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__72__A right_width_0_height_0__pin_46_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ top_width_0_height_0__pin_32_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_58_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ top_width_0_height_0__pin_8_ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_48_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ Test_en clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_40_ _40_/HI _40_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_1__f_clk_A clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__80__A top_width_0_height_0__pin_38_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_42_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__75__A right_width_0_height_0__pin_49_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ right_width_0_height_0__pin_29_ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_0_0_prog_clk_A clkbuf_4_1_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_1_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ top_width_0_height_0__pin_10_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _36_/HI ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_43_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__83__A top_width_0_height_0__pin_41_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_3_1_0_prog_clk clkbuf_3_1_0_prog_clk/A clkbuf_4_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__78__A top_width_0_height_0__pin_36_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5_0_prog_clk_A clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ top_width_0_height_0__pin_5_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _35_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ right_width_0_height_0__pin_28_ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_38_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_3_0_prog_clk clkbuf_4_3_0_prog_clk/A clkbuf_4_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _33_/HI ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ top_width_0_height_0__pin_40_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ top_width_0_height_0__pin_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_43_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _48_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_42_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _50_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _46_/HI ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_53_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ SC_OUT_BOT ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XFILLER_6_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_54_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_46_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_18_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _40_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_3_4_0_prog_clk_A clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _42_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_53_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_14_0_prog_clk_A clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_prog_clk clkbuf_3_1_0_prog_clk/A clkbuf_4_1_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_50_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_42_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _63_/HI ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_79_ top_width_0_height_0__pin_37_lower top_width_0_height_0__pin_37_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ top_width_0_height_0__pin_11_ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _32_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_2_0_prog_clk clkbuf_4_3_0_prog_clk/A clkbuf_4_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_31_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_54_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _34_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_45_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_78_ top_width_0_height_0__pin_36_lower top_width_0_height_0__pin_36_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_51_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_15_0_prog_clk clkbuf_3_7_0_prog_clk/X clkbuf_4_15_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_46_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3_0_prog_clk_A clkbuf_2_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ right_width_0_height_0__pin_18_ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_28_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _56_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _59_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _42_/HI ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ccff_tail clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_77_ top_width_0_height_0__pin_35_lower top_width_0_height_0__pin_35_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_51_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _58_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ right_width_0_height_0__pin_31_ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_62_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ right_width_0_height_0__pin_17_ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _40_/HI ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_45_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_60_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_60_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_76_ top_width_0_height_0__pin_34_lower top_width_0_height_0__pin_34_upper VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_59_ _59_/HI _59_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ right_width_0_height_0__pin_23_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XFILLER_46_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ right_width_0_height_0__pin_16_ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_1_0_prog_clk_A clkbuf_4_1_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _37_/HI ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_42_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_1_0_prog_clk clkbuf_4_1_0_prog_clk/A clkbuf_4_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_75_ right_width_0_height_0__pin_49_lower right_width_0_height_0__pin_49_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_64_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_58_ _58_/HI _58_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ right_width_0_height_0__pin_30_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_6_0_prog_clk_A clkbuf_4_7_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_14_0_prog_clk clkbuf_3_7_0_prog_clk/X clkbuf_4_14_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _49_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ Test_en clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_63_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ right_width_0_height_0__pin_25_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_74_ right_width_0_height_0__pin_48_lower right_width_0_height_0__pin_48_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_51_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_57_ _57_/HI _57_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ right_width_0_height_0__pin_20_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _38_/HI ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ top_width_0_height_0__pin_11_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _43_/HI ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_0_0_prog_clk_A clkbuf_3_1_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _41_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_73_ right_width_0_height_0__pin_47_lower right_width_0_height_0__pin_47_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_56_ _56_/HI _56_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f_clk clkbuf_0_clk/X clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_52_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_39_ _39_/HI _39_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_10_0_prog_clk_A clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _51_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_1_0__f_clk_A clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_5_0_prog_clk_A clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ right_width_0_height_0__pin_18_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__70__A right_width_0_height_0__pin_44_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ Test_en clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_72_ right_width_0_height_0__pin_46_lower right_width_0_height_0__pin_46_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_51_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_15_0_prog_clk_A clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__65__A SC_OUT_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_55_ _55_/HI _55_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _33_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_0_0_prog_clk clkbuf_4_1_0_prog_clk/A clkbuf_4_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ top_width_0_height_0__pin_13_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_38_ _38_/HI _38_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _52_/HI ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ top_width_0_height_0__pin_35_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ top_width_0_height_0__pin_6_ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__73__A right_width_0_height_0__pin_47_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_62_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__68__A right_width_0_height_0__pin_42_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_13_0_prog_clk clkbuf_3_6_0_prog_clk/X clkbuf_4_13_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ top_width_0_height_0__pin_8_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_71_ right_width_0_height_0__pin_45_lower right_width_0_height_0__pin_45_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_39_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__81__A top_width_0_height_0__pin_39_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _55_/HI ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_49_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ right_width_0_height_0__pin_19_ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XFILLER_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_54_ _54_/HI _54_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_52_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__76__A top_width_0_height_0__pin_34_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _47_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_37_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_37_ _37_/HI _37_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_16_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _57_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ top_width_0_height_0__pin_5_ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _44_/HI ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_47_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__79__A top_width_0_height_0__pin_37_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_70_ right_width_0_height_0__pin_44_lower right_width_0_height_0__pin_44_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_58_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_53_ _53_/HI _53_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_49_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ top_width_0_height_0__pin_6_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _34_/HI ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ right_width_0_height_0__pin_26_ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_36_ _36_/HI _36_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_60_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_43_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ top_width_0_height_0__pin_4_ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ top_width_0_height_0__pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _41_/HI ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_44_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_50_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_52_ _52_/HI _52_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ right_width_0_height_0__pin_25_ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_35_ _35_/HI _35_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_57_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ SC_IN_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_47_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_2_0_prog_clk_A clkbuf_4_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0_prog_clk clkbuf_3_6_0_prog_clk/X clkbuf_4_12_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_35_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_58_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_51_ _51_/HI _51_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_49_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_52_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ right_width_0_height_0__pin_24_ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_34_ _34_/HI _34_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7_0_prog_clk_A clkbuf_4_7_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_38_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_50_ _50_/HI _50_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_55_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_33_ _33_/HI _33_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_58_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_21_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f_clk clkbuf_0_clk/X clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_29_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_53_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _39_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _62_/HI ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_3_7_0_prog_clk clkbuf_3_6_0_prog_clk/A clkbuf_3_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_50_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_prog_clk_A clkbuf_3_1_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_61_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32_ _32_/HI _32_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_52_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_51_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ right_width_0_height_0__pin_31_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _56_/HI ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ top_width_0_height_0__pin_37_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_47_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_38_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_9_0_prog_clk clkbuf_4_9_0_prog_clk/A clkbuf_4_9_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_11_0_prog_clk_A clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_6_0_prog_clk_A clkbuf_3_6_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _35_/HI ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_58_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_38_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_50_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_31_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ top_width_0_height_0__pin_7_ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XFILLER_46_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_prog_clk clkbuf_3_5_0_prog_clk/X clkbuf_4_11_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_60_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_51_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XFILLER_18_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _53_/HI ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ top_width_0_height_0__pin_34_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_35_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _48_/HI ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_49_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_2_0_0_prog_clk_A clkbuf_2_1_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ top_width_0_height_0__pin_14_ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_59_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ right_width_0_height_0__pin_28_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_50_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ Test_en clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
XFILLER_53_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ right_width_0_height_0__pin_19_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ right_width_0_height_0__pin_27_ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _45_/HI ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_46_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_48_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_prog_clk clkbuf_3_6_0_prog_clk/A clkbuf_3_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_60_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ SC_OUT_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _44_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ top_width_0_height_0__pin_13_ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_59_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _58_/HI ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_62_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _46_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_53_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_8_0_prog_clk clkbuf_4_9_0_prog_clk/A clkbuf_4_8_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ right_width_0_height_0__pin_26_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_55_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__CLK
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ clkbuf_4_14_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_45_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_51_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ top_width_0_height_0__pin_12_ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_47_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _63_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_10_0_prog_clk clkbuf_3_5_0_prog_clk/X clkbuf_4_10_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_59_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ right_width_0_height_0__pin_21_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _36_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_47_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_38_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__CLK
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_44_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _38_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ Test_en clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ right_width_0_height_0__pin_16_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_4_3_0_prog_clk_A clkbuf_4_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_51_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__CLK
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ top_width_0_height_0__pin_7_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_3_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_3_6_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_28_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_38_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_53_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_prog_clk_A clkbuf_4_9_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _60_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__CLK
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_40_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__71__A right_width_0_height_0__pin_45_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_49_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__66__A SC_OUT_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _62_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__CLK
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_5_0_prog_clk clkbuf_2_2_0_prog_clk/X clkbuf_3_5_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_33_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ top_width_0_height_0__pin_14_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_69_ right_width_0_height_0__pin_43_lower right_width_0_height_0__pin_43_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _47_/HI ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6__CLK
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__74__A right_width_0_height_0__pin_48_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ _60_/HI ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ top_width_0_height_0__pin_39_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__CLK
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__69__A right_width_0_height_0__pin_43_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ top_width_0_height_0__pin_9_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _52_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_7_0_prog_clk clkbuf_4_7_0_prog_clk/A clkbuf_4_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_54_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ _54_/HI ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_45_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__82__A top_width_0_height_0__pin_40_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_63_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ SC_IN_BOT Test_en clkbuf_1_1__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__77__A top_width_0_height_0__pin_35_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_prog_clk_A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_68_ right_width_0_height_0__pin_42_lower right_width_0_height_0__pin_42_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_49_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14__CLK
+ clkbuf_4_12_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _54_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ top_width_0_height_0__pin_4_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_8_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
+ clkbuf_4_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_53_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ _57_/HI ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ top_width_0_height_0__pin_36_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12_0_prog_clk_A clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_7_0_prog_clk_A clkbuf_3_6_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__CLK
+ clkbuf_4_9_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3__CLK
+ clkbuf_4_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_48_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_1_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
+ clkbuf_1_0__f_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ clkbuf_4_11_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
+ clkbuf_4_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_67_ _67_/A bottom_width_0_height_0__pin_51_ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ top_width_0_height_0__pin_2_ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ top_width_0_height_0__pin_32_ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5__CLK
+ clkbuf_4_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__CLK
+ clkbuf_4_10_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_50_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ clkbuf_4_13_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ clkbuf_4_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_38_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_46_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ clkbuf_4_15_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_40_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_2_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_2_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ top_width_0_height_0__pin_2_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _59_/HI ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7__CLK
+ clkbuf_4_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_7.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _55_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_mode_fle_0.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ clkbuf_4_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_5.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_/D
+ top_width_0_height_0__pin_15_ ltile_clb_mode_0.ltile_clb_mode_fle_3.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XFILLER_36_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_mode_fle_4.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_2.ltile_clb_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_mode_fle_1.ltile_clb_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
+ ltile_clb_mode_0.ltile_clb_mode_fle_6.ltile_clb_physical__fabric_0.ltile_clb__frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

