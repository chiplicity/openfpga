* NGSPICE file created from sb_0__3_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

.subckt sb_0__3_ address[0] address[1] address[2] address[3] address[4] address[5]
+ bottom_left_grid_pin_11_ bottom_left_grid_pin_13_ bottom_left_grid_pin_15_ bottom_left_grid_pin_1_
+ bottom_left_grid_pin_3_ bottom_left_grid_pin_5_ bottom_left_grid_pin_7_ bottom_left_grid_pin_9_
+ bottom_right_grid_pin_11_ chanx_right_in[0] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4]
+ chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_out[0]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ data_in enable right_bottom_grid_pin_12_ right_top_grid_pin_11_ right_top_grid_pin_13_
+ right_top_grid_pin_15_ right_top_grid_pin_1_ right_top_grid_pin_3_ right_top_grid_pin_5_
+ right_top_grid_pin_7_ right_top_grid_pin_9_ vpwr vgnd
XFILLER_39_222 vgnd vpwr scs8hd_decap_12
Xmem_right_track_12.LATCH_1_.latch data_in _097_/A _143_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_166 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_41 vpwr vgnd scs8hd_fill_2
XFILLER_13_111 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_56 vpwr vgnd scs8hd_fill_2
XFILLER_3_12 vpwr vgnd scs8hd_fill_2
XFILLER_3_89 vpwr vgnd scs8hd_fill_2
XFILLER_8_192 vgnd vpwr scs8hd_decap_12
XFILLER_27_269 vgnd vpwr scs8hd_decap_8
XFILLER_6_107 vgnd vpwr scs8hd_fill_1
XFILLER_10_103 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _097_/A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_87 vgnd vpwr scs8hd_decap_4
XFILLER_12_98 vpwr vgnd scs8hd_fill_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_95 vgnd vpwr scs8hd_decap_8
XANTENNA__124__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_151 vgnd vpwr scs8hd_decap_3
XFILLER_24_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_200_ _200_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__209__A _209_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XFILLER_23_42 vpwr vgnd scs8hd_fill_2
X_131_ _162_/A _130_/X _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_121 vpwr vgnd scs8hd_fill_2
XFILLER_9_66 vgnd vpwr scs8hd_fill_1
XANTENNA__119__A _119_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _209_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _104_/Y mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_18_64 vgnd vpwr scs8hd_decap_4
XFILLER_11_220 vgnd vpwr scs8hd_decap_12
XFILLER_7_224 vgnd vpwr scs8hd_decap_12
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
X_114_ _114_/A _114_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _191_/HI _101_/Y mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__121__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_32 vpwr vgnd scs8hd_fill_2
XFILLER_29_74 vgnd vpwr scs8hd_decap_12
XFILLER_28_150 vgnd vpwr scs8hd_decap_3
XFILLER_6_23 vpwr vgnd scs8hd_fill_2
XANTENNA__132__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_fill_1
Xmem_right_track_8.LATCH_1_.latch data_in _093_/A _137_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_219 vgnd vpwr scs8hd_decap_12
XFILLER_1_208 vgnd vpwr scs8hd_decap_4
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _092_/A mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _118_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_274 vgnd vpwr scs8hd_decap_3
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XANTENNA__127__A address[3] vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _096_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_234 vgnd vpwr scs8hd_decap_8
XFILLER_39_201 vgnd vpwr scs8hd_decap_12
XFILLER_22_178 vgnd vpwr scs8hd_decap_12
XFILLER_26_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_20 vgnd vpwr scs8hd_decap_8
XFILLER_13_156 vgnd vpwr scs8hd_decap_12
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_138 vpwr vgnd scs8hd_fill_2
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_37_74 vgnd vpwr scs8hd_decap_6
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
XANTENNA__124__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _104_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB _175_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
XFILLER_23_262 vgnd vpwr scs8hd_decap_12
X_130_ address[3] _142_/B _142_/C _161_/D _130_/X vgnd vpwr scs8hd_or4_4
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA__135__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_9_34 vpwr vgnd scs8hd_fill_2
XFILLER_9_78 vpwr vgnd scs8hd_fill_2
XFILLER_14_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _120_/A vgnd
+ vpwr scs8hd_diode_2
X_113_ _113_/A _113_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_236 vgnd vpwr scs8hd_decap_8
XFILLER_11_232 vgnd vpwr scs8hd_decap_12
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _098_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _100_/A mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_37_162 vgnd vpwr scs8hd_decap_12
XFILLER_37_140 vgnd vpwr scs8hd_decap_3
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_20_66 vpwr vgnd scs8hd_fill_2
XFILLER_29_86 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_46 vgnd vpwr scs8hd_decap_4
XANTENNA__132__B _130_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_151 vgnd vpwr scs8hd_decap_12
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_10 vgnd vpwr scs8hd_decap_12
XFILLER_15_77 vpwr vgnd scs8hd_fill_2
XFILLER_15_99 vgnd vpwr scs8hd_decap_3
XFILLER_31_98 vgnd vpwr scs8hd_decap_12
XFILLER_31_135 vgnd vpwr scs8hd_decap_12
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _106_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__127__B address[2] vgnd vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vgnd vpwr scs8hd_decap_12
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_213 vpwr vgnd scs8hd_fill_2
XFILLER_30_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _087_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_76 vgnd vpwr scs8hd_decap_12
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _205_/A vgnd vpwr scs8hd_inv_1
XFILLER_3_69 vgnd vpwr scs8hd_decap_4
XFILLER_3_47 vpwr vgnd scs8hd_fill_2
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_10_138 vgnd vpwr scs8hd_fill_1
XFILLER_12_56 vpwr vgnd scs8hd_fill_2
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
XANTENNA__140__B _140_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB _146_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_208 vgnd vpwr scs8hd_decap_12
XFILLER_23_274 vgnd vpwr scs8hd_decap_3
XFILLER_23_77 vgnd vpwr scs8hd_decap_6
XFILLER_23_66 vpwr vgnd scs8hd_fill_2
XFILLER_23_99 vpwr vgnd scs8hd_fill_2
XFILLER_2_167 vgnd vpwr scs8hd_decap_4
XFILLER_0_37 vpwr vgnd scs8hd_fill_2
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
X_189_ _189_/HI _189_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__135__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_57 vgnd vpwr scs8hd_fill_1
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_20_255 vpwr vgnd scs8hd_fill_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
X_112_ _112_/A _112_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__146__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XFILLER_37_174 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _089_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_207 vgnd vpwr scs8hd_decap_6
Xmux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _087_/A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_23 vgnd vpwr scs8hd_decap_6
XFILLER_20_45 vgnd vpwr scs8hd_decap_6
XFILLER_20_89 vgnd vpwr scs8hd_fill_1
XFILLER_29_21 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_69 vgnd vpwr scs8hd_decap_6
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_163 vgnd vpwr scs8hd_decap_12
XFILLER_19_196 vgnd vpwr scs8hd_decap_12
XFILLER_40_158 vgnd vpwr scs8hd_decap_12
XFILLER_40_125 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_56 vgnd vpwr scs8hd_decap_3
XFILLER_31_22 vgnd vpwr scs8hd_decap_12
XFILLER_0_221 vpwr vgnd scs8hd_fill_2
XFILLER_16_144 vgnd vpwr scs8hd_decap_8
XFILLER_16_166 vgnd vpwr scs8hd_decap_12
XFILLER_31_147 vgnd vpwr scs8hd_decap_12
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C _142_/C vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _144_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_125 vgnd vpwr scs8hd_decap_4
Xmem_right_track_4.LATCH_1_.latch data_in _089_/A _131_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_26_88 vgnd vpwr scs8hd_decap_4
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _194_/HI _091_/Y mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XANTENNA__138__B _138_/B vgnd vpwr scs8hd_diode_2
XANTENNA__154__A address[0] vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_15_ mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_24 vpwr vgnd scs8hd_fill_2
XFILLER_12_35 vgnd vpwr scs8hd_decap_6
XFILLER_12_79 vpwr vgnd scs8hd_fill_2
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_18_239 vgnd vpwr scs8hd_decap_12
XFILLER_5_187 vpwr vgnd scs8hd_fill_2
XANTENNA__149__A address[3] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _119_/A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_220 vgnd vpwr scs8hd_decap_12
XFILLER_23_253 vpwr vgnd scs8hd_fill_2
XFILLER_23_23 vgnd vpwr scs8hd_decap_4
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_9_14 vgnd vpwr scs8hd_fill_1
X_188_ _188_/HI _188_/LO vgnd vpwr scs8hd_conb_1
XFILLER_29_3 vgnd vpwr scs8hd_decap_3
Xmux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _095_/A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__151__B _151_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_245 vgnd vpwr scs8hd_fill_1
XFILLER_18_45 vgnd vpwr scs8hd_decap_8
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
X_111_ _111_/A _111_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_245 vgnd vpwr scs8hd_decap_12
XANTENNA__146__B _147_/B vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _162_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_33 vgnd vpwr scs8hd_decap_12
XFILLER_20_79 vpwr vgnd scs8hd_fill_2
XFILLER_29_99 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _195_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_7 vgnd vpwr scs8hd_fill_1
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_19_175 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _190_/HI _099_/Y mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_123 vgnd vpwr scs8hd_decap_12
XFILLER_25_112 vpwr vgnd scs8hd_fill_2
XFILLER_25_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_24 vpwr vgnd scs8hd_fill_2
XFILLER_15_35 vpwr vgnd scs8hd_fill_2
XFILLER_31_34 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_244 vgnd vpwr scs8hd_decap_4
XFILLER_16_123 vpwr vgnd scs8hd_fill_2
XFILLER_16_178 vgnd vpwr scs8hd_decap_12
XFILLER_31_159 vgnd vpwr scs8hd_decap_12
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__D _139_/D vgnd vpwr scs8hd_diode_2
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_259 vpwr vgnd scs8hd_fill_2
XFILLER_39_248 vpwr vgnd scs8hd_fill_2
XFILLER_11_3 vgnd vpwr scs8hd_decap_3
XFILLER_22_104 vgnd vpwr scs8hd_decap_6
XFILLER_26_45 vgnd vpwr scs8hd_decap_8
XFILLER_13_115 vgnd vpwr scs8hd_decap_4
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_16 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _090_/A mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__154__B _153_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_163 vpwr vgnd scs8hd_fill_2
XANTENNA__170__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_107 vgnd vpwr scs8hd_fill_1
XFILLER_10_129 vgnd vpwr scs8hd_decap_3
XANTENNA__080__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_37_11 vgnd vpwr scs8hd_decap_12
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__149__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_17_262 vgnd vpwr scs8hd_decap_12
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_232 vgnd vpwr scs8hd_decap_12
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_23_46 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_13_ mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_125 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/HI _187_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_90 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _094_/Y mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_20_202 vgnd vpwr scs8hd_decap_12
XFILLER_18_68 vgnd vpwr scs8hd_fill_1
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XFILLER_11_257 vgnd vpwr scs8hd_decap_12
X_110_ _110_/A _110_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _117_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _095_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__B _163_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_154 vpwr vgnd scs8hd_fill_2
XFILLER_37_132 vpwr vgnd scs8hd_fill_2
XFILLER_1_71 vpwr vgnd scs8hd_fill_2
XFILLER_1_82 vpwr vgnd scs8hd_fill_2
XFILLER_29_45 vgnd vpwr scs8hd_decap_12
XFILLER_28_154 vgnd vpwr scs8hd_decap_12
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XANTENNA__157__B _156_/B vgnd vpwr scs8hd_diode_2
XANTENNA__173__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_25_135 vgnd vpwr scs8hd_decap_12
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _098_/A mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__083__A enable vgnd vpwr scs8hd_diode_2
XFILLER_31_46 vgnd vpwr scs8hd_decap_12
XFILLER_0_212 vgnd vpwr scs8hd_decap_4
XFILLER_24_190 vgnd vpwr scs8hd_decap_12
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_102 vpwr vgnd scs8hd_fill_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _103_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_138 vgnd vpwr scs8hd_decap_12
XFILLER_7_92 vpwr vgnd scs8hd_fill_2
XFILLER_13_149 vgnd vpwr scs8hd_decap_4
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_171 vgnd vpwr scs8hd_decap_12
XANTENNA__170__B _142_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _119_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_23 vgnd vpwr scs8hd_decap_12
XFILLER_26_263 vgnd vpwr scs8hd_decap_12
Xmem_right_track_0.LATCH_1_.latch data_in _086_/A _124_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _097_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ _102_/Y mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_5_134 vpwr vgnd scs8hd_fill_2
XFILLER_5_156 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__149__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_17_274 vgnd vpwr scs8hd_decap_3
XANTENNA__165__B _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vpwr vgnd scs8hd_fill_2
XFILLER_2_104 vgnd vpwr scs8hd_decap_6
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_148 vgnd vpwr scs8hd_decap_4
XFILLER_9_38 vpwr vgnd scs8hd_fill_2
X_186_ _186_/HI _186_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _090_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__176__A _139_/D vgnd vpwr scs8hd_diode_2
XFILLER_18_14 vpwr vgnd scs8hd_fill_2
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
XFILLER_1_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _105_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_10.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_11_ mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_169_ address[0] _169_/B _169_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_7.LATCH_0_.latch data_in _110_/A _163_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_57 vgnd vpwr scs8hd_decap_4
XFILLER_28_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_111 vpwr vgnd scs8hd_fill_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_34_125 vgnd vpwr scs8hd_decap_12
XANTENNA__173__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_25_147 vgnd vpwr scs8hd_decap_12
XFILLER_31_58 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _086_/A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _169_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_180 vgnd vpwr scs8hd_decap_3
XANTENNA__094__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _092_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_132 vpwr vgnd scs8hd_fill_2
XFILLER_16_80 vgnd vpwr scs8hd_fill_1
XANTENNA__170__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_12_16 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.tap_buf4_0_.scs8hd_inv_1 mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _198_/A vgnd vpwr scs8hd_inv_1
XFILLER_37_35 vgnd vpwr scs8hd_decap_12
XANTENNA__089__A _089_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_168 vpwr vgnd scs8hd_fill_2
XANTENNA__149__D _161_/D vgnd vpwr scs8hd_diode_2
XFILLER_17_220 vgnd vpwr scs8hd_decap_12
XFILLER_17_253 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _193_/HI _089_/Y mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_50 vpwr vgnd scs8hd_fill_2
XFILLER_23_245 vgnd vpwr scs8hd_decap_8
XFILLER_9_28 vgnd vpwr scs8hd_decap_4
X_185_ _185_/HI _185_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_6.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_160 vgnd vpwr scs8hd_decap_3
XFILLER_1_193 vpwr vgnd scs8hd_fill_2
XANTENNA__176__B _174_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_215 vgnd vpwr scs8hd_decap_12
XFILLER_20_259 vgnd vpwr scs8hd_decap_12
XFILLER_18_26 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _117_/A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_24_80 vgnd vpwr scs8hd_decap_12
X_168_ _162_/A _169_/B _168_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_3 vgnd vpwr scs8hd_decap_4
X_099_ _099_/A _099_/Y vgnd vpwr scs8hd_inv_8
XFILLER_28_178 vgnd vpwr scs8hd_decap_12
XANTENNA__097__A _097_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_15.LATCH_0_.latch data_in _118_/A _175_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_71 vgnd vpwr scs8hd_decap_4
XFILLER_10_93 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_137 vgnd vpwr scs8hd_decap_12
XFILLER_19_134 vpwr vgnd scs8hd_fill_2
XANTENNA__173__C address[4] vgnd vpwr scs8hd_diode_2
XFILLER_25_159 vgnd vpwr scs8hd_decap_12
XFILLER_15_16 vpwr vgnd scs8hd_fill_2
XFILLER_0_258 vpwr vgnd scs8hd_fill_2
XFILLER_0_225 vgnd vpwr scs8hd_decap_12
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_81 vgnd vpwr scs8hd_fill_1
XFILLER_39_218 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_38_251 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.tap_buf4_0_.scs8hd_inv_1 mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _201_/A vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_15_ mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_59 vgnd vpwr scs8hd_decap_8
Xmux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _189_/HI _097_/Y mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_12
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_12_151 vpwr vgnd scs8hd_fill_2
XANTENNA__170__D _139_/D vgnd vpwr scs8hd_diode_2
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XFILLER_12_28 vgnd vpwr scs8hd_decap_3
XFILLER_37_47 vgnd vpwr scs8hd_decap_12
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_114 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _211_/A vgnd vpwr scs8hd_inv_1
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XFILLER_27_80 vpwr vgnd scs8hd_fill_2
XFILLER_17_232 vgnd vpwr scs8hd_decap_12
XFILLER_4_84 vpwr vgnd scs8hd_fill_2
XFILLER_4_40 vgnd vpwr scs8hd_fill_1
Xmux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _088_/A mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
X_184_ _184_/HI _184_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__176__C _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
X_098_ _098_/A _098_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_231 vgnd vpwr scs8hd_decap_12
X_167_ _161_/A _142_/B _161_/C _161_/D _169_/B vgnd vpwr scs8hd_or4_4
Xmux_right_track_4.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_102 vgnd vpwr scs8hd_decap_12
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _092_/Y mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XFILLER_34_149 vgnd vpwr scs8hd_decap_4
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_92 vgnd vpwr scs8hd_fill_1
XANTENNA__173__D _080_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_105 vpwr vgnd scs8hd_fill_2
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XFILLER_25_116 vgnd vpwr scs8hd_decap_6
XFILLER_15_39 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_3.LATCH_0_.latch data_in _106_/A _157_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_127 vpwr vgnd scs8hd_fill_2
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_2 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _120_/A mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_15_160 vgnd vpwr scs8hd_decap_12
XFILLER_30_141 vgnd vpwr scs8hd_decap_12
XFILLER_7_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _120_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XFILLER_26_16 vpwr vgnd scs8hd_fill_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _098_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_119 vgnd vpwr scs8hd_fill_1
XFILLER_21_196 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _096_/A mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_145 vpwr vgnd scs8hd_fill_2
XFILLER_8_167 vgnd vpwr scs8hd_decap_4
XFILLER_12_163 vgnd vpwr scs8hd_decap_12
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_15.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _106_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_183_ _183_/HI _183_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_80 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _100_/Y mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_20_239 vgnd vpwr scs8hd_decap_6
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
X_097_ _097_/A _097_/Y vgnd vpwr scs8hd_inv_8
X_166_ address[0] _164_/X _166_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_243 vgnd vpwr scs8hd_decap_12
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
XFILLER_37_136 vpwr vgnd scs8hd_fill_2
XFILLER_37_114 vpwr vgnd scs8hd_fill_2
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XFILLER_37_158 vpwr vgnd scs8hd_fill_2
XFILLER_1_75 vpwr vgnd scs8hd_fill_2
XFILLER_1_86 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _100_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_114 vgnd vpwr scs8hd_decap_12
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_3_202 vgnd vpwr scs8hd_decap_12
XFILLER_10_84 vgnd vpwr scs8hd_decap_8
XFILLER_19_71 vpwr vgnd scs8hd_fill_2
XFILLER_34_117 vgnd vpwr scs8hd_decap_6
X_149_ address[3] address[2] _161_/C _161_/D _151_/B vgnd vpwr scs8hd_or4_4
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _207_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
XFILLER_0_216 vgnd vpwr scs8hd_fill_1
Xmux_right_track_2.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_106 vgnd vpwr scs8hd_decap_4
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_50 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_11.LATCH_0_.latch data_in _114_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_172 vgnd vpwr scs8hd_decap_8
XFILLER_7_52 vgnd vpwr scs8hd_decap_3
XFILLER_26_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _108_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_220 vgnd vpwr scs8hd_decap_12
XFILLER_8_102 vgnd vpwr scs8hd_decap_3
XFILLER_16_83 vgnd vpwr scs8hd_decap_6
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _089_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_175 vgnd vpwr scs8hd_decap_12
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_60 vgnd vpwr scs8hd_fill_1
XFILLER_17_245 vgnd vpwr scs8hd_decap_8
XFILLER_40_270 vgnd vpwr scs8hd_decap_4
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_97 vgnd vpwr scs8hd_decap_3
XFILLER_23_29 vpwr vgnd scs8hd_fill_2
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
X_182_ _182_/HI _182_/LO vgnd vpwr scs8hd_conb_1
XFILLER_22_270 vgnd vpwr scs8hd_decap_4
XFILLER_13_95 vgnd vpwr scs8hd_decap_3
XFILLER_1_174 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A _100_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_11_ mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_18 vgnd vpwr scs8hd_decap_8
Xmux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _192_/HI _087_/Y mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_251 vgnd vpwr scs8hd_decap_12
X_165_ _162_/A _164_/X _165_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
X_096_ _096_/A _096_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_255 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.INVTX1_0_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_21 vpwr vgnd scs8hd_fill_2
XFILLER_20_19 vpwr vgnd scs8hd_fill_2
XFILLER_29_17 vpwr vgnd scs8hd_fill_2
XFILLER_28_126 vgnd vpwr scs8hd_decap_12
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XFILLER_3_214 vgnd vpwr scs8hd_decap_12
XFILLER_10_30 vgnd vpwr scs8hd_fill_1
XFILLER_10_52 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _091_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_115 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _115_/A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_148_ address[4] _080_/Y _161_/C vgnd vpwr scs8hd_nand2_4
XFILLER_25_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_151 vpwr vgnd scs8hd_fill_2
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_73 vpwr vgnd scs8hd_fill_2
XFILLER_21_95 vpwr vgnd scs8hd_fill_2
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vgnd vpwr scs8hd_decap_12
XFILLER_7_31 vpwr vgnd scs8hd_fill_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_143 vpwr vgnd scs8hd_fill_2
XFILLER_29_232 vgnd vpwr scs8hd_decap_12
XFILLER_12_121 vpwr vgnd scs8hd_fill_2
XFILLER_12_187 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _176_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__103__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _182_/HI _119_/Y mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _188_/HI _095_/Y mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_54 vgnd vpwr scs8hd_decap_4
XFILLER_4_32 vgnd vpwr scs8hd_decap_6
XFILLER_4_10 vpwr vgnd scs8hd_fill_2
XFILLER_23_19 vpwr vgnd scs8hd_fill_2
XFILLER_14_205 vgnd vpwr scs8hd_decap_8
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
XFILLER_13_30 vpwr vgnd scs8hd_fill_2
X_181_ _181_/HI _181_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_131 vpwr vgnd scs8hd_fill_2
Xmem_right_track_14.LATCH_0_.latch data_in _100_/A _147_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_1_197 vgnd vpwr scs8hd_decap_4
XFILLER_9_220 vgnd vpwr scs8hd_decap_12
XFILLER_11_208 vgnd vpwr scs8hd_decap_12
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ _085_/A mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_095_ _095_/A _095_/Y vgnd vpwr scs8hd_inv_8
XFILLER_24_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_267 vgnd vpwr scs8hd_decap_8
XFILLER_10_263 vgnd vpwr scs8hd_decap_12
X_164_ _161_/A address[2] _161_/C _139_/D _164_/X vgnd vpwr scs8hd_or4_4
XFILLER_27_7 vgnd vpwr scs8hd_fill_1
XANTENNA__111__A _111_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_138 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_11.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_9_ mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_226 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_171 vgnd vpwr scs8hd_decap_12
XFILLER_19_51 vgnd vpwr scs8hd_decap_4
XFILLER_19_95 vgnd vpwr scs8hd_decap_4
XFILLER_19_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__106__A _106_/A vgnd vpwr scs8hd_diode_2
X_147_ address[0] _147_/B _147_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _188_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.INVTX1_0_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _090_/Y mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_15_196 vgnd vpwr scs8hd_decap_12
XFILLER_38_211 vgnd vpwr scs8hd_decap_3
XFILLER_8_115 vpwr vgnd scs8hd_fill_2
XFILLER_12_199 vgnd vpwr scs8hd_decap_12
XFILLER_16_63 vpwr vgnd scs8hd_fill_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XFILLER_7_181 vpwr vgnd scs8hd_fill_2
XFILLER_7_192 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _118_/A mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_84 vpwr vgnd scs8hd_fill_2
XFILLER_27_62 vgnd vpwr scs8hd_decap_3
XFILLER_27_40 vgnd vpwr scs8hd_decap_12
XFILLER_17_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_195 vgnd vpwr scs8hd_decap_12
XFILLER_4_88 vgnd vpwr scs8hd_decap_4
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_239 vgnd vpwr scs8hd_decap_12
X_180_ _180_/HI _180_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _178_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_53 vgnd vpwr scs8hd_decap_3
XANTENNA__109__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_232 vgnd vpwr scs8hd_decap_12
X_094_ _094_/A _094_/Y vgnd vpwr scs8hd_inv_8
X_163_ address[0] _163_/B _163_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
XFILLER_1_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _119_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _097_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _098_/Y mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__212__A _212_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_238 vgnd vpwr scs8hd_decap_6
XFILLER_10_32 vgnd vpwr scs8hd_decap_6
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
XANTENNA__122__A address[1] vgnd vpwr scs8hd_diode_2
X_146_ _162_/A _147_/B _146_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_208 vpwr vgnd scs8hd_fill_2
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_131 vgnd vpwr scs8hd_decap_12
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
XFILLER_7_88 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_3 vgnd vpwr scs8hd_fill_1
X_129_ address[0] _129_/B _129_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _111_/A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _105_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_123 vgnd vpwr scs8hd_decap_3
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
XFILLER_16_20 vgnd vpwr scs8hd_decap_6
Xmem_bottom_track_7.LATCH_1_.latch data_in _109_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_3.INVTX1_0_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_149 vpwr vgnd scs8hd_fill_2
XFILLER_12_134 vgnd vpwr scs8hd_decap_8
XFILLER_12_145 vgnd vpwr scs8hd_decap_4
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
XFILLER_27_52 vgnd vpwr scs8hd_decap_8
XFILLER_40_251 vgnd vpwr scs8hd_decap_4
XFILLER_4_163 vpwr vgnd scs8hd_fill_2
XFILLER_4_152 vgnd vpwr scs8hd_fill_1
XFILLER_4_67 vgnd vpwr scs8hd_decap_6
XFILLER_4_23 vpwr vgnd scs8hd_fill_2
XANTENNA__130__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_31_262 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _099_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_144 vpwr vgnd scs8hd_fill_2
XFILLER_38_84 vgnd vpwr scs8hd_decap_8
XANTENNA__125__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _092_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_192 vpwr vgnd scs8hd_fill_2
XFILLER_39_170 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_162_ _162_/A _163_/B _162_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_20 vgnd vpwr scs8hd_decap_8
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
X_093_ _093_/A _093_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_118 vpwr vgnd scs8hd_fill_2
XFILLER_1_13 vpwr vgnd scs8hd_fill_2
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
Xmem_right_track_10.LATCH_0_.latch data_in _096_/A _141_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _107_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_151 vpwr vgnd scs8hd_fill_2
XFILLER_10_22 vpwr vgnd scs8hd_fill_2
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XFILLER_19_75 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _187_/HI _086_/Y mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_145_ _161_/A _142_/B _142_/C _139_/D _147_/B vgnd vpwr scs8hd_or4_4
XANTENNA__122__B _122_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_143 vgnd vpwr scs8hd_decap_8
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_12
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_54 vgnd vpwr scs8hd_fill_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_132 vpwr vgnd scs8hd_fill_2
XANTENNA__133__A address[3] vgnd vpwr scs8hd_diode_2
X_128_ _162_/A _129_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_3 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _113_/A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XFILLER_12_102 vpwr vgnd scs8hd_fill_2
XFILLER_16_43 vgnd vpwr scs8hd_decap_3
XFILLER_16_76 vgnd vpwr scs8hd_decap_4
XFILLER_8_128 vpwr vgnd scs8hd_fill_2
XFILLER_20_190 vgnd vpwr scs8hd_decap_12
XANTENNA__128__A _162_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_15.LATCH_1_.latch data_in _117_/A _174_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _094_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XFILLER_40_274 vgnd vpwr scs8hd_fill_1
XFILLER_4_175 vgnd vpwr scs8hd_decap_12
XANTENNA__130__B _142_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_274 vgnd vpwr scs8hd_decap_3
XFILLER_13_11 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _181_/HI _117_/Y mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_274 vgnd vpwr scs8hd_fill_1
XFILLER_13_77 vpwr vgnd scs8hd_fill_2
XFILLER_1_178 vgnd vpwr scs8hd_decap_3
XFILLER_1_156 vpwr vgnd scs8hd_fill_2
XFILLER_1_101 vgnd vpwr scs8hd_decap_6
XFILLER_1_123 vpwr vgnd scs8hd_fill_2
Xmem_right_track_6.LATCH_0_.latch data_in _092_/A _135_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__125__B _124_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XANTENNA__141__A address[0] vgnd vpwr scs8hd_diode_2
X_161_ _161_/A address[2] _161_/C _161_/D _163_/B vgnd vpwr scs8hd_or4_4
XFILLER_24_32 vgnd vpwr scs8hd_decap_3
XFILLER_10_211 vgnd vpwr scs8hd_decap_3
X_092_ _092_/A _092_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__136__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_67 vpwr vgnd scs8hd_fill_2
XFILLER_19_21 vgnd vpwr scs8hd_decap_4
XFILLER_19_32 vpwr vgnd scs8hd_fill_2
XFILLER_19_119 vgnd vpwr scs8hd_fill_1
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_213_ _213_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
X_144_ address[0] _144_/B _144_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.tap_buf4_0_.scs8hd_inv_1 mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _203_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_152 vgnd vpwr scs8hd_fill_1
XFILLER_18_163 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_166 vgnd vpwr scs8hd_decap_12
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_22 vpwr vgnd scs8hd_fill_2
XFILLER_21_33 vpwr vgnd scs8hd_fill_2
XFILLER_21_77 vgnd vpwr scs8hd_decap_4
XFILLER_21_99 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_111 vpwr vgnd scs8hd_fill_2
XANTENNA__133__B _142_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_35 vpwr vgnd scs8hd_fill_2
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
X_127_ address[3] address[2] _142_/C _139_/D _129_/B vgnd vpwr scs8hd_or4_4
XFILLER_16_3 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _213_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
XFILLER_21_147 vgnd vpwr scs8hd_decap_12
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_107 vgnd vpwr scs8hd_decap_8
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA__128__B _129_/B vgnd vpwr scs8hd_diode_2
XANTENNA__144__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_7_151 vpwr vgnd scs8hd_fill_2
XFILLER_7_173 vpwr vgnd scs8hd_fill_2
XFILLER_7_184 vgnd vpwr scs8hd_decap_8
Xmux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _088_/Y mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_26_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_76 vpwr vgnd scs8hd_fill_2
XFILLER_27_32 vpwr vgnd scs8hd_fill_2
XFILLER_27_21 vpwr vgnd scs8hd_fill_2
XFILLER_27_10 vpwr vgnd scs8hd_fill_2
XFILLER_4_187 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_3.LATCH_1_.latch data_in _105_/A _156_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__130__C _142_/C vgnd vpwr scs8hd_diode_2
XFILLER_31_253 vpwr vgnd scs8hd_fill_2
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA__139__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_34 vpwr vgnd scs8hd_fill_2
XFILLER_1_113 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _116_/A mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_13_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
XANTENNA__141__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_40_21 vgnd vpwr scs8hd_decap_8
XFILLER_24_44 vgnd vpwr scs8hd_decap_12
X_091_ _091_/A _091_/Y vgnd vpwr scs8hd_inv_8
X_160_ address[0] _159_/B _160_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__136__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__152__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_36_131 vgnd vpwr scs8hd_decap_12
XFILLER_27_120 vpwr vgnd scs8hd_fill_2
XFILLER_19_88 vgnd vpwr scs8hd_decap_4
XFILLER_19_99 vgnd vpwr scs8hd_fill_1
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
X_212_ _212_/A chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
X_143_ _162_/A _144_/B _143_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _120_/Y mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_142 vpwr vgnd scs8hd_fill_2
XFILLER_18_175 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _189_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__147__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_178 vgnd vpwr scs8hd_decap_12
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _096_/Y mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_7_14 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__133__C _142_/C vgnd vpwr scs8hd_diode_2
X_126_ address[1] enable _139_/D vgnd vpwr scs8hd_nand2_4
XFILLER_7_69 vpwr vgnd scs8hd_fill_2
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_21_159 vgnd vpwr scs8hd_decap_12
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_16_89 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _100_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__144__B _144_/B vgnd vpwr scs8hd_diode_2
X_109_ _109_/A _109_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_196 vpwr vgnd scs8hd_fill_2
XANTENNA__160__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
XFILLER_27_88 vpwr vgnd scs8hd_fill_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _109_/A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_144 vpwr vgnd scs8hd_fill_2
XFILLER_4_122 vgnd vpwr scs8hd_decap_3
XANTENNA__130__D _161_/D vgnd vpwr scs8hd_diode_2
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XANTENNA__155__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_16_251 vgnd vpwr scs8hd_decap_12
XANTENNA__139__B address[2] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_11.LATCH_1_.latch data_in _113_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_6 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _183_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _108_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_91 vpwr vgnd scs8hd_fill_2
XFILLER_39_184 vgnd vpwr scs8hd_decap_8
XFILLER_39_162 vgnd vpwr scs8hd_decap_8
XFILLER_24_56 vgnd vpwr scs8hd_decap_4
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
X_090_ _090_/A _090_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_38 vpwr vgnd scs8hd_fill_2
XANTENNA__136__C _142_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__152__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XFILLER_36_143 vgnd vpwr scs8hd_decap_8
XFILLER_36_121 vgnd vpwr scs8hd_fill_1
Xmem_right_track_2.LATCH_0_.latch data_in _088_/A _129_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
X_211_ _211_/A chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
X_142_ _161_/A _142_/B _142_/C _161_/D _144_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _102_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
XANTENNA__147__B _147_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_187 vgnd vpwr scs8hd_decap_12
XANTENNA__163__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_102 vgnd vpwr scs8hd_decap_8
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_46 vpwr vgnd scs8hd_fill_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_30_105 vgnd vpwr scs8hd_decap_12
X_125_ address[0] _124_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_48 vpwr vgnd scs8hd_fill_2
XFILLER_30_7 vpwr vgnd scs8hd_fill_2
XANTENNA__133__D _139_/D vgnd vpwr scs8hd_diode_2
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XANTENNA__158__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_16_35 vpwr vgnd scs8hd_fill_2
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _110_/A vgnd
+ vpwr scs8hd_diode_2
X_108_ _108_/A _108_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__160__B _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _091_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _114_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_208 vgnd vpwr scs8hd_decap_12
XFILLER_4_167 vgnd vpwr scs8hd_decap_4
XFILLER_4_27 vpwr vgnd scs8hd_fill_2
XANTENNA__139__C _142_/C vgnd vpwr scs8hd_diode_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__155__B _142_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
XANTENNA__171__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_58 vgnd vpwr scs8hd_decap_3
XFILLER_1_148 vpwr vgnd scs8hd_fill_2
XANTENNA__081__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _179_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__166__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_8_270 vgnd vpwr scs8hd_decap_4
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_1_17 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _180_/HI _115_/Y mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__136__D _161_/D vgnd vpwr scs8hd_diode_2
XANTENNA__152__C _161_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _112_/A mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XFILLER_10_26 vpwr vgnd scs8hd_fill_2
XFILLER_10_48 vpwr vgnd scs8hd_fill_2
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
X_210_ _210_/A chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
X_141_ address[0] _140_/B _141_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_147 vgnd vpwr scs8hd_decap_12
XFILLER_18_199 vgnd vpwr scs8hd_decap_12
XANTENNA__163__B _163_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_14.LATCH_1_.latch data_in _099_/A _146_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _093_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_60 vpwr vgnd scs8hd_fill_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
XFILLER_15_136 vpwr vgnd scs8hd_fill_2
XFILLER_23_180 vgnd vpwr scs8hd_decap_3
X_124_ _162_/A _124_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
XANTENNA__158__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA__174__A _161_/D vgnd vpwr scs8hd_diode_2
XFILLER_21_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_106 vpwr vgnd scs8hd_fill_2
XFILLER_12_117 vpwr vgnd scs8hd_fill_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XANTENNA__084__A address[0] vgnd vpwr scs8hd_diode_2
X_107_ _107_/A _107_/Y vgnd vpwr scs8hd_inv_8
XFILLER_14_3 vpwr vgnd scs8hd_fill_2
XANTENNA__169__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_19_261 vgnd vpwr scs8hd_decap_12
XFILLER_25_220 vgnd vpwr scs8hd_decap_12
XFILLER_4_113 vgnd vpwr scs8hd_decap_4
XANTENNA__139__D _139_/D vgnd vpwr scs8hd_diode_2
XFILLER_17_90 vgnd vpwr scs8hd_decap_3
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_8
XANTENNA__155__C _161_/C vgnd vpwr scs8hd_diode_2
XANTENNA__171__B _172_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_15 vpwr vgnd scs8hd_fill_2
XFILLER_1_127 vpwr vgnd scs8hd_fill_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ _085_/Y mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_160 vgnd vpwr scs8hd_fill_1
XANTENNA__166__B _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_71 vgnd vpwr scs8hd_decap_4
XFILLER_39_197 vpwr vgnd scs8hd_fill_2
XFILLER_39_175 vpwr vgnd scs8hd_fill_2
XFILLER_24_69 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__092__A _092_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_219 vgnd vpwr scs8hd_decap_12
XFILLER_5_241 vgnd vpwr scs8hd_decap_3
XANTENNA__152__D _139_/D vgnd vpwr scs8hd_diode_2
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XANTENNA__177__A _139_/D vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _114_/A mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_38 vgnd vpwr scs8hd_fill_1
XFILLER_27_101 vpwr vgnd scs8hd_fill_2
XFILLER_19_47 vpwr vgnd scs8hd_fill_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_27_123 vgnd vpwr scs8hd_decap_12
XFILLER_27_112 vgnd vpwr scs8hd_decap_8
XANTENNA__087__A _087_/A vgnd vpwr scs8hd_diode_2
X_140_ _162_/A _140_/B _140_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_159 vgnd vpwr scs8hd_decap_12
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_129 vgnd vpwr scs8hd_decap_12
XFILLER_15_115 vgnd vpwr scs8hd_decap_4
X_123_ address[3] address[2] _142_/C _161_/D _124_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__158__C _161_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_14_181 vgnd vpwr scs8hd_decap_12
XANTENNA__174__B _174_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _118_/Y mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_16_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_162 vpwr vgnd scs8hd_fill_2
XFILLER_11_173 vpwr vgnd scs8hd_fill_2
XFILLER_7_155 vpwr vgnd scs8hd_fill_2
XFILLER_7_177 vpwr vgnd scs8hd_fill_2
X_106_ _106_/A _106_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_184 vgnd vpwr scs8hd_decap_12
XANTENNA__169__B _169_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XFILLER_19_273 vgnd vpwr scs8hd_decap_4
XFILLER_27_36 vpwr vgnd scs8hd_fill_2
XFILLER_27_25 vpwr vgnd scs8hd_fill_2
XFILLER_25_232 vgnd vpwr scs8hd_decap_12
XANTENNA__095__A _095_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__155__D _161_/D vgnd vpwr scs8hd_diode_2
XFILLER_3_191 vpwr vgnd scs8hd_fill_2
XFILLER_13_38 vgnd vpwr scs8hd_decap_4
XFILLER_22_202 vgnd vpwr scs8hd_decap_12
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_1_117 vgnd vpwr scs8hd_decap_3
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
XFILLER_0_172 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_9_ mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _107_/A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_132 vpwr vgnd scs8hd_fill_2
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
XFILLER_6_6 vpwr vgnd scs8hd_fill_2
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
XANTENNA__177__B _174_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_135 vgnd vpwr scs8hd_decap_12
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _099_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_102 vpwr vgnd scs8hd_fill_2
XFILLER_18_146 vgnd vpwr scs8hd_decap_6
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_26_190 vgnd vpwr scs8hd_decap_12
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ _199_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_2_84 vpwr vgnd scs8hd_fill_2
XFILLER_2_73 vpwr vgnd scs8hd_fill_2
XFILLER_2_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _190_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _186_/HI _111_/Y mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__098__A _098_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_18 vpwr vgnd scs8hd_fill_2
XFILLER_15_149 vgnd vpwr scs8hd_decap_8
X_122_ address[1] _122_/B _161_/D vgnd vpwr scs8hd_or2_4
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_9 vgnd vpwr scs8hd_fill_1
XANTENNA__158__D _139_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_193 vgnd vpwr scs8hd_decap_12
XANTENNA__174__C _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_208 vgnd vpwr scs8hd_decap_12
XFILLER_16_16 vpwr vgnd scs8hd_fill_2
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
Xmem_right_track_10.LATCH_1_.latch data_in _095_/A _140_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_152 vgnd vpwr scs8hd_fill_1
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _107_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_123 vpwr vgnd scs8hd_fill_2
XFILLER_7_134 vpwr vgnd scs8hd_fill_2
X_105_ _105_/A _105_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_141 vgnd vpwr scs8hd_decap_6
XFILLER_11_196 vgnd vpwr scs8hd_decap_12
XFILLER_40_258 vgnd vpwr scs8hd_decap_12
XFILLER_4_148 vgnd vpwr scs8hd_decap_4
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_258 vpwr vgnd scs8hd_fill_2
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_247 vpwr vgnd scs8hd_fill_2
XFILLER_22_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _101_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _184_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_251 vgnd vpwr scs8hd_decap_4
XFILLER_39_144 vgnd vpwr scs8hd_decap_3
XFILLER_39_100 vgnd vpwr scs8hd_decap_12
XFILLER_5_95 vgnd vpwr scs8hd_decap_8
XFILLER_24_16 vpwr vgnd scs8hd_fill_2
XFILLER_40_15 vgnd vpwr scs8hd_decap_3
XFILLER_10_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _094_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__177__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_10_18 vpwr vgnd scs8hd_fill_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_147 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_7_ mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_180 vgnd vpwr scs8hd_decap_3
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_2_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _109_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_125 vpwr vgnd scs8hd_fill_2
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_25_81 vgnd vpwr scs8hd_decap_4
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ _198_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _113_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _179_/HI _113_/Y mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_6.LATCH_1_.latch data_in _091_/A _134_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _110_/A mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_121_ address[4] address[5] _142_/C vgnd vpwr scs8hd_or2_4
XFILLER_11_83 vpwr vgnd scs8hd_fill_2
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XFILLER_14_150 vgnd vpwr scs8hd_decap_3
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
XFILLER_16_28 vgnd vpwr scs8hd_decap_3
XFILLER_16_39 vpwr vgnd scs8hd_fill_2
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_113 vgnd vpwr scs8hd_decap_3
XFILLER_7_168 vgnd vpwr scs8hd_decap_3
XFILLER_11_131 vgnd vpwr scs8hd_fill_1
X_104_ _104_/A _104_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_60 vgnd vpwr scs8hd_fill_1
XFILLER_19_220 vgnd vpwr scs8hd_decap_12
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_8_73 vpwr vgnd scs8hd_fill_2
XFILLER_8_84 vpwr vgnd scs8hd_fill_2
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vgnd vpwr scs8hd_decap_12
XFILLER_4_127 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_182 vgnd vpwr scs8hd_fill_1
XFILLER_12_3 vpwr vgnd scs8hd_fill_2
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_9_208 vgnd vpwr scs8hd_decap_12
XFILLER_0_196 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _180_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_274 vgnd vpwr scs8hd_fill_1
XFILLER_39_112 vgnd vpwr scs8hd_fill_1
XFILLER_24_28 vgnd vpwr scs8hd_fill_1
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
XFILLER_36_115 vgnd vpwr scs8hd_decap_6
XFILLER_19_17 vpwr vgnd scs8hd_fill_2
XFILLER_19_28 vpwr vgnd scs8hd_fill_2
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XFILLER_27_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _085_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_14.tap_buf4_0_.scs8hd_inv_1 mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _197_/A vgnd vpwr scs8hd_inv_1
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
X_197_ _197_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_181 vpwr vgnd scs8hd_fill_2
XFILLER_21_18 vpwr vgnd scs8hd_fill_2
XFILLER_21_29 vpwr vgnd scs8hd_fill_2
XFILLER_23_184 vgnd vpwr scs8hd_decap_12
X_120_ _120_/A _120_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_4.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_5_ mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_51 vpwr vgnd scs8hd_fill_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_154 vgnd vpwr scs8hd_decap_12
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
X_103_ _103_/A _103_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_72 vgnd vpwr scs8hd_decap_12
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_14_7 vpwr vgnd scs8hd_fill_2
XFILLER_19_232 vgnd vpwr scs8hd_decap_12
XFILLER_8_52 vgnd vpwr scs8hd_decap_8
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_139 vgnd vpwr scs8hd_decap_3
XFILLER_4_117 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _116_/Y mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_16_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_83 vpwr vgnd scs8hd_fill_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_172 vpwr vgnd scs8hd_fill_2
XFILLER_22_227 vgnd vpwr scs8hd_decap_12
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_31 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_75 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_15.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_39_179 vgnd vpwr scs8hd_decap_4
XFILLER_5_212 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _200_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XFILLER_39_70 vgnd vpwr scs8hd_decap_8
XFILLER_36_105 vgnd vpwr scs8hd_decap_8
XANTENNA__101__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_105 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _105_/A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_6 vpwr vgnd scs8hd_fill_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_138 vpwr vgnd scs8hd_fill_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
X_196_ _196_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _210_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_10 vpwr vgnd scs8hd_fill_2
XFILLER_24_119 vgnd vpwr scs8hd_decap_12
XFILLER_32_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_119 vgnd vpwr scs8hd_fill_1
XFILLER_23_196 vgnd vpwr scs8hd_decap_12
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_179_ _179_/HI _179_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_122 vgnd vpwr scs8hd_decap_8
XFILLER_20_144 vgnd vpwr scs8hd_decap_8
XFILLER_20_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _185_/HI _109_/Y mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_2.LATCH_1_.latch data_in _087_/A _128_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_100 vpwr vgnd scs8hd_fill_2
XFILLER_11_111 vpwr vgnd scs8hd_fill_2
X_102_ _102_/A _102_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_177 vgnd vpwr scs8hd_decap_6
Xmux_right_track_2.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_3_ mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _102_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_40_206 vgnd vpwr scs8hd_decap_8
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_17_62 vpwr vgnd scs8hd_fill_2
XFILLER_17_95 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_239 vgnd vpwr scs8hd_decap_8
XFILLER_0_121 vgnd vpwr scs8hd_fill_1
XFILLER_0_176 vgnd vpwr scs8hd_decap_8
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_43 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_9.LATCH_0_.latch data_in _112_/A _166_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_158 vpwr vgnd scs8hd_fill_2
XFILLER_39_136 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _110_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_29 vpwr vgnd scs8hd_fill_2
XFILLER_14_30 vgnd vpwr scs8hd_fill_1
XFILLER_14_41 vgnd vpwr scs8hd_decap_4
XFILLER_14_52 vpwr vgnd scs8hd_fill_2
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _114_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_13.INVTX1_0_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_106 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vgnd vpwr scs8hd_decap_4
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ _195_/HI _195_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_7 vpwr vgnd scs8hd_fill_2
XFILLER_2_77 vpwr vgnd scs8hd_fill_2
XFILLER_2_44 vgnd vpwr scs8hd_fill_1
XFILLER_1_271 vgnd vpwr scs8hd_decap_6
XANTENNA__112__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vpwr vgnd scs8hd_fill_2
XFILLER_17_161 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _191_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__107__A _107_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_142 vgnd vpwr scs8hd_decap_8
X_178_ _178_/HI _178_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
XFILLER_28_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_178 vgnd vpwr scs8hd_decap_12
X_101_ _101_/A _101_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_105 vpwr vgnd scs8hd_fill_2
XFILLER_7_138 vpwr vgnd scs8hd_fill_2
XFILLER_11_123 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _108_/A mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_245 vpwr vgnd scs8hd_fill_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_10 vpwr vgnd scs8hd_fill_2
XFILLER_8_32 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _112_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__210__A _210_/A vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _093_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _116_/A vgnd
+ vpwr scs8hd_diode_2
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XANTENNA__120__A _120_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_1_ mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_240 vpwr vgnd scs8hd_fill_2
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _206_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _185_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_251 vgnd vpwr scs8hd_decap_12
XANTENNA__115__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_115 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _112_/Y mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _187_/HI vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_17.LATCH_0_.latch data_in _120_/A _177_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_30 vgnd vpwr scs8hd_fill_1
XFILLER_5_203 vgnd vpwr scs8hd_fill_1
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_14_86 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XFILLER_26_151 vpwr vgnd scs8hd_fill_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_85 vgnd vpwr scs8hd_fill_1
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _194_/HI _194_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_56 vpwr vgnd scs8hd_fill_2
XFILLER_2_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_17_173 vgnd vpwr scs8hd_decap_8
XFILLER_17_184 vgnd vpwr scs8hd_decap_12
XFILLER_23_132 vgnd vpwr scs8hd_decap_12
XANTENNA__213__A _213_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_21 vpwr vgnd scs8hd_fill_2
XFILLER_11_65 vpwr vgnd scs8hd_fill_2
XFILLER_11_87 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB _174_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.INVTX1_0_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_121 vpwr vgnd scs8hd_fill_2
X_177_ _139_/D _174_/B address[0] _177_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA__123__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_20_102 vpwr vgnd scs8hd_fill_2
XFILLER_9_180 vgnd vpwr scs8hd_decap_3
XFILLER_28_202 vgnd vpwr scs8hd_decap_12
X_100_ _100_/A _100_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__208__A _208_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_86 vgnd vpwr scs8hd_decap_4
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_77 vpwr vgnd scs8hd_fill_2
XFILLER_8_88 vgnd vpwr scs8hd_decap_4
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_4_109 vpwr vgnd scs8hd_fill_2
XFILLER_17_20 vpwr vgnd scs8hd_fill_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XFILLER_3_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XFILLER_13_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _086_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_263 vgnd vpwr scs8hd_decap_12
XFILLER_0_156 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_74 vgnd vpwr scs8hd_decap_12
XFILLER_8_212 vpwr vgnd scs8hd_fill_2
XFILLER_12_263 vgnd vpwr scs8hd_decap_12
XFILLER_5_78 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _114_/Y mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _181_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__131__A _162_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_65 vpwr vgnd scs8hd_fill_2
XFILLER_39_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_171 vgnd vpwr scs8hd_decap_12
XANTENNA__126__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_5.LATCH_0_.latch data_in _108_/A _160_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XFILLER_25_31 vgnd vpwr scs8hd_fill_1
XFILLER_25_20 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_18_119 vgnd vpwr scs8hd_decap_4
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_193_ _193_/HI _193_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_251 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_35 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_17_196 vgnd vpwr scs8hd_decap_12
XFILLER_23_144 vgnd vpwr scs8hd_decap_12
XFILLER_2_6 vpwr vgnd scs8hd_fill_2
XFILLER_11_55 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _103_/A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_176_ _139_/D _174_/B _162_/A _176_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA__123__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_11_158 vpwr vgnd scs8hd_fill_2
XFILLER_11_169 vpwr vgnd scs8hd_fill_2
XFILLER_22_10 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vgnd vpwr scs8hd_decap_3
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XANTENNA__134__A _162_/A vgnd vpwr scs8hd_diode_2
X_159_ _162_/A _159_/B _159_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_239 vgnd vpwr scs8hd_decap_12
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_198 vpwr vgnd scs8hd_fill_2
XFILLER_3_187 vpwr vgnd scs8hd_fill_2
XFILLER_3_176 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _184_/HI _107_/Y mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__129__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_220 vgnd vpwr scs8hd_decap_12
XFILLER_21_275 vpwr vgnd scs8hd_fill_2
XFILLER_0_113 vpwr vgnd scs8hd_fill_2
XFILLER_0_135 vgnd vpwr scs8hd_decap_3
XFILLER_28_86 vgnd vpwr scs8hd_decap_6
XANTENNA__131__B _130_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_35 vpwr vgnd scs8hd_fill_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XFILLER_14_11 vpwr vgnd scs8hd_fill_2
XFILLER_14_22 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XFILLER_39_96 vpwr vgnd scs8hd_fill_2
XFILLER_39_41 vgnd vpwr scs8hd_decap_12
XANTENNA__126__B enable vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_131 vgnd vpwr scs8hd_decap_12
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/HI _192_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_14.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_track_13.LATCH_0_.latch data_in _116_/A _172_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XANTENNA__137__A _162_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _101_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_156 vgnd vpwr scs8hd_decap_12
XFILLER_23_112 vpwr vgnd scs8hd_fill_2
XFILLER_11_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__123__C _142_/C vgnd vpwr scs8hd_diode_2
X_175_ _161_/D _174_/B address[0] _175_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_104 vpwr vgnd scs8hd_fill_2
XFILLER_11_115 vpwr vgnd scs8hd_fill_2
XFILLER_22_44 vpwr vgnd scs8hd_fill_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
X_089_ _089_/A _089_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__134__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_163 vpwr vgnd scs8hd_fill_2
XFILLER_6_174 vpwr vgnd scs8hd_fill_2
X_158_ address[3] _142_/B _161_/C _139_/D _159_/B vgnd vpwr scs8hd_or4_4
XFILLER_26_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _109_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__150__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_66 vpwr vgnd scs8hd_fill_2
XFILLER_17_99 vpwr vgnd scs8hd_fill_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _113_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_155 vpwr vgnd scs8hd_fill_2
XANTENNA__129__B _129_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A _161_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _106_/A mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_232 vgnd vpwr scs8hd_decap_8
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_8_258 vgnd vpwr scs8hd_decap_12
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_14 vpwr vgnd scs8hd_fill_2
XFILLER_38_151 vpwr vgnd scs8hd_fill_2
XFILLER_30_11 vgnd vpwr scs8hd_decap_4
XFILLER_5_217 vgnd vpwr scs8hd_decap_12
XFILLER_14_45 vgnd vpwr scs8hd_fill_1
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XFILLER_39_53 vgnd vpwr scs8hd_decap_8
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__B _142_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_132 vgnd vpwr scs8hd_decap_12
XFILLER_35_110 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _110_/Y mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_2_209 vgnd vpwr scs8hd_decap_4
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vgnd vpwr scs8hd_decap_12
XFILLER_26_143 vgnd vpwr scs8hd_decap_8
XFILLER_25_88 vpwr vgnd scs8hd_fill_2
XFILLER_25_77 vpwr vgnd scs8hd_fill_2
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
X_191_ _191_/HI _191_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_231 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _111_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__137__B _138_/B vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_168 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _115_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_102 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_0_.latch data_in _104_/A _154_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_157 vgnd vpwr scs8hd_decap_12
XFILLER_22_190 vgnd vpwr scs8hd_decap_12
XANTENNA__123__D _161_/D vgnd vpwr scs8hd_diode_2
X_174_ _161_/D _174_/B _162_/A _174_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_28_7 vgnd vpwr scs8hd_fill_1
XANTENNA__148__A address[4] vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_172 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XFILLER_7_109 vpwr vgnd scs8hd_fill_2
XFILLER_11_127 vpwr vgnd scs8hd_fill_2
XFILLER_22_23 vgnd vpwr scs8hd_decap_8
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
XFILLER_19_249 vgnd vpwr scs8hd_decap_12
X_157_ address[0] _156_/B _157_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_69 vpwr vgnd scs8hd_fill_2
X_088_ _088_/A _088_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__150__B _151_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_208 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _085_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_263 vgnd vpwr scs8hd_decap_12
XFILLER_17_45 vpwr vgnd scs8hd_fill_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_11 vgnd vpwr scs8hd_decap_12
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_16.LATCH_0_.latch data_in _102_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_123 vpwr vgnd scs8hd_fill_2
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
X_209_ _209_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__145__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_211 vgnd vpwr scs8hd_decap_3
XFILLER_8_204 vgnd vpwr scs8hd_decap_8
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XFILLER_39_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _186_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_10.tap_buf4_0_.scs8hd_inv_1 mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _199_/A vgnd vpwr scs8hd_inv_1
XANTENNA__156__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_163 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _192_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_5_229 vgnd vpwr scs8hd_decap_12
XFILLER_39_10 vgnd vpwr scs8hd_decap_8
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
XANTENNA__142__C _142_/C vgnd vpwr scs8hd_diode_2
XFILLER_35_144 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_45 vpwr vgnd scs8hd_fill_2
XFILLER_25_34 vpwr vgnd scs8hd_fill_2
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
X_190_ _190_/HI _190_/LO vgnd vpwr scs8hd_conb_1
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_2_27 vpwr vgnd scs8hd_fill_2
XFILLER_1_243 vgnd vpwr scs8hd_fill_1
XFILLER_17_133 vpwr vgnd scs8hd_fill_2
XANTENNA__153__B _153_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _088_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_69 vgnd vpwr scs8hd_decap_3
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XFILLER_14_125 vpwr vgnd scs8hd_fill_2
X_173_ address[3] address[2] address[4] _080_/Y _174_/B vgnd vpwr scs8hd_or4_4
XFILLER_14_169 vgnd vpwr scs8hd_decap_12
XANTENNA__148__B _080_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_106 vgnd vpwr scs8hd_decap_3
XFILLER_20_139 vgnd vpwr scs8hd_decap_3
XFILLER_9_151 vgnd vpwr scs8hd_decap_3
XFILLER_9_184 vgnd vpwr scs8hd_decap_12
XANTENNA__164__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
X_156_ _162_/A _156_/B _156_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_150 vgnd vpwr scs8hd_fill_1
X_087_ _087_/A _087_/Y vgnd vpwr scs8hd_inv_8
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XANTENNA__159__A _162_/A vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_23 vgnd vpwr scs8hd_decap_12
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_10.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_24 vpwr vgnd scs8hd_fill_2
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XFILLER_17_79 vpwr vgnd scs8hd_fill_2
XFILLER_3_102 vpwr vgnd scs8hd_fill_2
XFILLER_3_113 vgnd vpwr scs8hd_decap_3
XFILLER_15_220 vgnd vpwr scs8hd_decap_12
XANTENNA__145__C _142_/C vgnd vpwr scs8hd_diode_2
XANTENNA__161__B address[2] vgnd vpwr scs8hd_diode_2
X_208_ _208_/A chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
X_139_ _161_/A address[2] _142_/C _139_/D _140_/B vgnd vpwr scs8hd_or4_4
Xmux_right_track_4.tap_buf4_0_.scs8hd_inv_1 mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _202_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_245 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_67 vgnd vpwr scs8hd_decap_3
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _182_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__172__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _156_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_175 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _183_/HI _105_/Y mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _212_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_69 vpwr vgnd scs8hd_fill_2
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XFILLER_5_208 vpwr vgnd scs8hd_fill_2
XANTENNA__082__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_39_88 vgnd vpwr scs8hd_decap_4
XFILLER_39_66 vpwr vgnd scs8hd_fill_2
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XANTENNA__142__D _161_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_156 vgnd vpwr scs8hd_decap_12
XANTENNA__167__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_178 vgnd vpwr scs8hd_decap_12
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_255 vpwr vgnd scs8hd_fill_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_3
XFILLER_40_170 vgnd vpwr scs8hd_decap_12
XFILLER_15_90 vgnd vpwr scs8hd_decap_3
Xmem_bottom_track_9.LATCH_1_.latch data_in _111_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _093_/A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
X_172_ address[0] _172_/B _172_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__164__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_9_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_60 vgnd vpwr scs8hd_fill_1
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XANTENNA__090__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
XFILLER_8_38 vgnd vpwr scs8hd_fill_1
X_086_ _086_/A _086_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_100 vgnd vpwr scs8hd_decap_4
X_155_ address[3] _142_/B _161_/C _161_/D _156_/B vgnd vpwr scs8hd_or4_4
XFILLER_12_91 vgnd vpwr scs8hd_fill_1
XFILLER_33_7 vpwr vgnd scs8hd_fill_2
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_251 vgnd vpwr scs8hd_decap_12
XANTENNA__175__A _161_/D vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_35 vgnd vpwr scs8hd_decap_12
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XANTENNA__085__A _085_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_232 vgnd vpwr scs8hd_decap_12
X_207_ _207_/A chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_30_202 vgnd vpwr scs8hd_decap_12
XANTENNA__145__D _139_/D vgnd vpwr scs8hd_diode_2
XANTENNA__161__C _161_/C vgnd vpwr scs8hd_diode_2
X_138_ address[0] _138_/B _138_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_180 vgnd vpwr scs8hd_decap_8
XFILLER_0_72 vpwr vgnd scs8hd_fill_2
XFILLER_0_94 vpwr vgnd scs8hd_fill_2
XFILLER_0_117 vgnd vpwr scs8hd_decap_4
XFILLER_28_35 vgnd vpwr scs8hd_decap_12
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_39 vpwr vgnd scs8hd_fill_2
Xmem_right_track_12.LATCH_0_.latch data_in _098_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__172__B _172_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_187 vgnd vpwr scs8hd_decap_12
XFILLER_14_26 vpwr vgnd scs8hd_fill_2
XFILLER_14_48 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _104_/A mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_39_78 vgnd vpwr scs8hd_decap_3
XFILLER_29_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _112_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _101_/A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_35_168 vgnd vpwr scs8hd_decap_12
XANTENNA__167__B _142_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _116_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_102 vgnd vpwr scs8hd_decap_8
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XANTENNA__093__A _093_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_6
XFILLER_17_146 vgnd vpwr scs8hd_decap_8
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XFILLER_17_157 vpwr vgnd scs8hd_fill_2
XFILLER_40_182 vgnd vpwr scs8hd_decap_12
XFILLER_23_116 vgnd vpwr scs8hd_decap_4
XFILLER_31_171 vgnd vpwr scs8hd_decap_12
XFILLER_16_190 vgnd vpwr scs8hd_decap_12
XFILLER_11_38 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A _088_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XFILLER_14_138 vpwr vgnd scs8hd_fill_2
X_171_ _162_/A _172_/B _171_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _108_/Y mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_1_.latch data_in _119_/A _176_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__164__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_13_171 vpwr vgnd scs8hd_fill_2
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XFILLER_11_119 vgnd vpwr scs8hd_decap_3
XFILLER_22_48 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_19_208 vgnd vpwr scs8hd_decap_12
X_154_ address[0] _153_/B _154_/Y vgnd vpwr scs8hd_nor2_4
X_085_ _085_/A _085_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_134 vpwr vgnd scs8hd_fill_2
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
XFILLER_6_167 vgnd vpwr scs8hd_decap_4
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
XFILLER_10_163 vgnd vpwr scs8hd_decap_12
XANTENNA__175__B _174_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _208_/A vgnd vpwr scs8hd_inv_1
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_47 vgnd vpwr scs8hd_decap_12
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_159 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_0_.latch data_in _094_/A _138_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_206_ _206_/A chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
X_137_ _162_/A _138_/B _137_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__161__D _161_/D vgnd vpwr scs8hd_diode_2
XFILLER_17_3 vpwr vgnd scs8hd_fill_2
XFILLER_0_84 vpwr vgnd scs8hd_fill_2
XFILLER_9_60 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _118_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_82 vpwr vgnd scs8hd_fill_2
XFILLER_28_47 vgnd vpwr scs8hd_decap_12
XFILLER_0_129 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _096_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__096__A _096_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_18 vpwr vgnd scs8hd_fill_2
XFILLER_38_199 vgnd vpwr scs8hd_decap_12
XFILLER_38_133 vgnd vpwr scs8hd_decap_12
XFILLER_39_24 vpwr vgnd scs8hd_fill_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XANTENNA__167__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_61 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _104_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_40_194 vgnd vpwr scs8hd_decap_12
XFILLER_32_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _086_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_17 vpwr vgnd scs8hd_fill_2
XFILLER_14_106 vgnd vpwr scs8hd_decap_4
X_170_ _161_/A _142_/B _161_/C _139_/D _172_/B vgnd vpwr scs8hd_or4_4
XFILLER_22_150 vgnd vpwr scs8hd_decap_3
XANTENNA__164__D _139_/D vgnd vpwr scs8hd_diode_2
XFILLER_3_73 vgnd vpwr scs8hd_fill_1
XFILLER_3_51 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_7_ mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__099__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_220 vgnd vpwr scs8hd_decap_12
X_153_ _162_/A _153_/B _153_/Y vgnd vpwr scs8hd_nor2_4
Xmem_bottom_track_5.LATCH_1_.latch data_in _107_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_142 vgnd vpwr scs8hd_decap_8
XFILLER_10_175 vgnd vpwr scs8hd_decap_12
X_084_ address[0] _162_/A vgnd vpwr scs8hd_inv_8
XFILLER_12_60 vpwr vgnd scs8hd_fill_2
XFILLER_12_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
XANTENNA__175__C address[0] vgnd vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_16 vpwr vgnd scs8hd_fill_2
XFILLER_17_49 vpwr vgnd scs8hd_fill_2
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_138 vpwr vgnd scs8hd_fill_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_15_245 vgnd vpwr scs8hd_decap_12
X_205_ _205_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
X_136_ _161_/A address[2] _142_/C _161_/D _138_/B vgnd vpwr scs8hd_or4_4
XFILLER_31_6 vpwr vgnd scs8hd_fill_2
XFILLER_0_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_259 vpwr vgnd scs8hd_fill_2
XFILLER_28_59 vgnd vpwr scs8hd_decap_8
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _087_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
X_119_ _119_/A _119_/Y vgnd vpwr scs8hd_inv_8
XFILLER_38_145 vgnd vpwr scs8hd_decap_4
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _193_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XANTENNA__167__D _161_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XFILLER_25_49 vpwr vgnd scs8hd_fill_2
XFILLER_25_27 vgnd vpwr scs8hd_decap_4
XFILLER_25_16 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_9_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _178_/HI _103_/Y mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_32_129 vgnd vpwr scs8hd_decap_12
XFILLER_40_151 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_184 vgnd vpwr scs8hd_decap_12
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XFILLER_3_85 vpwr vgnd scs8hd_fill_2
XFILLER_27_232 vgnd vpwr scs8hd_decap_12
X_083_ enable _122_/B vgnd vpwr scs8hd_inv_8
XFILLER_10_110 vgnd vpwr scs8hd_decap_8
XFILLER_10_187 vgnd vpwr scs8hd_decap_12
X_152_ address[3] address[2] _161_/C _139_/D _153_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_83 vpwr vgnd scs8hd_fill_2
XFILLER_37_80 vgnd vpwr scs8hd_fill_1
Xmux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _091_/A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_180 vgnd vpwr scs8hd_decap_3
XFILLER_5_191 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_13.LATCH_1_.latch data_in _115_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_28 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_7.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_5_ mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_106 vpwr vgnd scs8hd_fill_2
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
X_204_ _204_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
X_135_ address[0] _135_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_9_51 vgnd vpwr scs8hd_decap_6
XFILLER_9_62 vgnd vpwr scs8hd_decap_4
XFILLER_0_109 vpwr vgnd scs8hd_fill_2
XFILLER_12_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_271 vgnd vpwr scs8hd_decap_4
XFILLER_18_71 vpwr vgnd scs8hd_fill_2
X_118_ _118_/A _118_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_253 vpwr vgnd scs8hd_fill_2
Xmem_right_track_4.LATCH_0_.latch data_in _090_/A _132_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_39_37 vpwr vgnd scs8hd_fill_2
XFILLER_29_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_83 vgnd vpwr scs8hd_decap_6
XFILLER_28_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_1_215 vpwr vgnd scs8hd_fill_2
XFILLER_1_204 vpwr vgnd scs8hd_fill_2
XFILLER_1_259 vgnd vpwr scs8hd_decap_12
XFILLER_25_171 vgnd vpwr scs8hd_decap_12
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
XFILLER_39_252 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _099_/A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_263 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_9_101 vpwr vgnd scs8hd_fill_2
XFILLER_9_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_156 vgnd vpwr scs8hd_decap_3
XFILLER_13_196 vgnd vpwr scs8hd_decap_12
X_151_ address[0] _151_/B _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_104 vgnd vpwr scs8hd_fill_1
X_082_ address[2] _142_/B vgnd vpwr scs8hd_inv_8
XFILLER_10_199 vgnd vpwr scs8hd_decap_12
XFILLER_18_211 vgnd vpwr scs8hd_decap_3
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _106_/Y mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _111_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
X_203_ _203_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
XFILLER_23_94 vgnd vpwr scs8hd_decap_3
XFILLER_2_140 vgnd vpwr scs8hd_decap_6
X_134_ _162_/A _135_/B _134_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_10 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_1_.latch data_in _103_/A _153_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _115_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_0_76 vpwr vgnd scs8hd_fill_2
XFILLER_0_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_17 vgnd vpwr scs8hd_decap_12
XFILLER_12_239 vgnd vpwr scs8hd_decap_12
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
X_117_ _117_/A _117_/Y vgnd vpwr scs8hd_inv_8
Xmux_bottom_track_5.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_3_ mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_3 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _094_/A mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_30_18 vgnd vpwr scs8hd_decap_12
XFILLER_29_103 vgnd vpwr scs8hd_decap_12
XFILLER_29_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_213 vgnd vpwr scs8hd_fill_1
XFILLER_20_62 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_1_.latch data_in _101_/A _150_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_42 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_40_131 vgnd vpwr scs8hd_decap_12
XFILLER_40_120 vgnd vpwr scs8hd_decap_3
XFILLER_15_73 vpwr vgnd scs8hd_fill_2
XFILLER_15_95 vpwr vgnd scs8hd_fill_2
XANTENNA__102__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_275 vpwr vgnd scs8hd_fill_2
XFILLER_39_242 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_153 vgnd vpwr scs8hd_fill_1
XFILLER_13_175 vgnd vpwr scs8hd_decap_8
XFILLER_9_168 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _117_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_65 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _095_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_12
X_150_ _162_/A _151_/B _150_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_138 vgnd vpwr scs8hd_decap_4
XFILLER_6_149 vpwr vgnd scs8hd_fill_2
X_081_ address[3] _161_/A vgnd vpwr scs8hd_inv_8
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _088_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_62 vpwr vgnd scs8hd_fill_2
X_202_ _202_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
X_133_ address[3] _142_/B _142_/C _139_/D _135_/B vgnd vpwr scs8hd_or4_4
XFILLER_2_163 vpwr vgnd scs8hd_fill_2
XFILLER_2_152 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ _102_/A mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_88 vgnd vpwr scs8hd_decap_3
XFILLER_9_97 vpwr vgnd scs8hd_fill_2
XFILLER_28_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _103_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_84 vgnd vpwr scs8hd_decap_6
XFILLER_7_200 vgnd vpwr scs8hd_decap_12
XANTENNA__105__A _105_/A vgnd vpwr scs8hd_diode_2
X_116_ _116_/A _116_/Y vgnd vpwr scs8hd_inv_8
XFILLER_39_28 vgnd vpwr scs8hd_decap_6
XFILLER_29_159 vgnd vpwr scs8hd_decap_12
XFILLER_29_115 vgnd vpwr scs8hd_decap_6
XFILLER_35_118 vpwr vgnd scs8hd_fill_2
XFILLER_29_94 vpwr vgnd scs8hd_fill_2
XFILLER_6_10 vpwr vgnd scs8hd_fill_2
XFILLER_6_32 vgnd vpwr scs8hd_fill_1
XFILLER_6_65 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_1_ mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_right_track_0.LATCH_0_.latch data_in _085_/A _125_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_17_129 vpwr vgnd scs8hd_fill_2
XFILLER_40_143 vgnd vpwr scs8hd_decap_8
XFILLER_25_184 vgnd vpwr scs8hd_decap_12
XFILLER_15_52 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XFILLER_31_110 vgnd vpwr scs8hd_decap_12
XFILLER_16_140 vpwr vgnd scs8hd_fill_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_121 vpwr vgnd scs8hd_fill_2
XFILLER_22_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _090_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_33 vgnd vpwr scs8hd_decap_3
XFILLER_8_180 vgnd vpwr scs8hd_decap_12
XFILLER_27_257 vgnd vpwr scs8hd_decap_12
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
X_080_ address[5] _080_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_117 vgnd vpwr scs8hd_decap_6
XFILLER_12_20 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _204_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_3 vpwr vgnd scs8hd_fill_2
XFILLER_12_75 vpwr vgnd scs8hd_fill_2
XFILLER_37_83 vgnd vpwr scs8hd_decap_12
XANTENNA__108__A _108_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_172 vgnd vpwr scs8hd_decap_8
XFILLER_24_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_201_ _201_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
X_132_ address[0] _130_/X _132_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_197 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _196_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_9_10 vgnd vpwr scs8hd_decap_4
XFILLER_21_208 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _089_/A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__211__A _211_/A vgnd vpwr scs8hd_diode_2
X_115_ _115_/A _115_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_212 vgnd vpwr scs8hd_decap_12
XFILLER_7_245 vgnd vpwr scs8hd_decap_8
XFILLER_38_116 vgnd vpwr scs8hd_decap_8
XFILLER_38_105 vgnd vpwr scs8hd_decap_8
XANTENNA__121__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_22_6 vpwr vgnd scs8hd_fill_2
XFILLER_37_182 vgnd vpwr scs8hd_fill_1
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _194_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_decap_12
XANTENNA__116__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_119 vgnd vpwr scs8hd_decap_12
XFILLER_20_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _195_/HI _093_/Y mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_196 vgnd vpwr scs8hd_decap_12
XFILLER_15_20 vpwr vgnd scs8hd_fill_2
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XFILLER_0_262 vgnd vpwr scs8hd_decap_12
XFILLER_0_240 vpwr vgnd scs8hd_fill_2
XFILLER_16_152 vgnd vpwr scs8hd_fill_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

