magic
tech EFS8A
magscale 1 2
timestamp 1604349141
<< locali >>
rect 26525 13175 26559 13277
rect 16037 12631 16071 12869
rect 32413 12631 32447 12733
rect 2973 10999 3007 11101
rect 3709 10999 3743 11101
rect 8953 10455 8987 10557
rect 3065 8823 3099 9061
rect 26801 5015 26835 5253
rect 25697 4675 25731 4777
rect 26985 3927 27019 4165
<< viali >>
rect 4261 13481 4295 13515
rect 5365 13481 5399 13515
rect 31585 13481 31619 13515
rect 34437 13481 34471 13515
rect 36737 13481 36771 13515
rect 1685 13413 1719 13447
rect 2329 13413 2363 13447
rect 21649 13413 21683 13447
rect 25697 13413 25731 13447
rect 27445 13413 27479 13447
rect 30297 13413 30331 13447
rect 4077 13345 4111 13379
rect 5181 13345 5215 13379
rect 6929 13345 6963 13379
rect 21373 13345 21407 13379
rect 22661 13345 22695 13379
rect 22937 13345 22971 13379
rect 30113 13345 30147 13379
rect 31401 13345 31435 13379
rect 33149 13345 33183 13379
rect 34253 13345 34287 13379
rect 35449 13345 35483 13379
rect 36553 13345 36587 13379
rect 2237 13277 2271 13311
rect 2421 13277 2455 13311
rect 25697 13277 25731 13311
rect 25789 13277 25823 13311
rect 26525 13277 26559 13311
rect 27353 13277 27387 13311
rect 27537 13277 27571 13311
rect 30389 13277 30423 13311
rect 31217 13277 31251 13311
rect 2789 13209 2823 13243
rect 7113 13209 7147 13243
rect 33333 13209 33367 13243
rect 1869 13141 1903 13175
rect 14749 13141 14783 13175
rect 16497 13141 16531 13175
rect 24317 13141 24351 13175
rect 24685 13141 24719 13175
rect 25053 13141 25087 13175
rect 25237 13141 25271 13175
rect 26249 13141 26283 13175
rect 26525 13141 26559 13175
rect 26617 13141 26651 13175
rect 26985 13141 27019 13175
rect 29469 13141 29503 13175
rect 29837 13141 29871 13175
rect 35633 13141 35667 13175
rect 4629 12937 4663 12971
rect 5181 12937 5215 12971
rect 7021 12937 7055 12971
rect 7481 12937 7515 12971
rect 25513 12937 25547 12971
rect 35633 12937 35667 12971
rect 37105 12937 37139 12971
rect 2329 12869 2363 12903
rect 7849 12869 7883 12903
rect 14841 12869 14875 12903
rect 15853 12869 15887 12903
rect 16037 12869 16071 12903
rect 16497 12869 16531 12903
rect 21557 12869 21591 12903
rect 24041 12869 24075 12903
rect 24593 12869 24627 12903
rect 27629 12869 27663 12903
rect 29009 12869 29043 12903
rect 29653 12869 29687 12903
rect 31217 12869 31251 12903
rect 3985 12801 4019 12835
rect 5733 12801 5767 12835
rect 10333 12801 10367 12835
rect 13645 12801 13679 12835
rect 3617 12733 3651 12767
rect 3801 12733 3835 12767
rect 5457 12733 5491 12767
rect 6285 12733 6319 12767
rect 6837 12733 6871 12767
rect 10057 12733 10091 12767
rect 13369 12733 13403 12767
rect 2605 12665 2639 12699
rect 2881 12665 2915 12699
rect 14289 12665 14323 12699
rect 15117 12665 15151 12699
rect 15301 12665 15335 12699
rect 15393 12665 15427 12699
rect 24869 12801 24903 12835
rect 26433 12801 26467 12835
rect 28089 12801 28123 12835
rect 30205 12801 30239 12835
rect 30665 12801 30699 12835
rect 30941 12801 30975 12835
rect 32873 12801 32907 12835
rect 36001 12801 36035 12835
rect 16313 12733 16347 12767
rect 17049 12733 17083 12767
rect 22937 12733 22971 12767
rect 24685 12733 24719 12767
rect 26047 12733 26081 12767
rect 28641 12733 28675 12767
rect 31493 12733 31527 12767
rect 32137 12733 32171 12767
rect 32413 12733 32447 12767
rect 32689 12733 32723 12767
rect 35449 12733 35483 12767
rect 36553 12733 36587 12767
rect 16773 12665 16807 12699
rect 21005 12665 21039 12699
rect 21833 12665 21867 12699
rect 22109 12665 22143 12699
rect 26617 12665 26651 12699
rect 27077 12665 27111 12699
rect 28181 12665 28215 12699
rect 29929 12665 29963 12699
rect 30113 12665 30147 12699
rect 31677 12665 31711 12699
rect 31769 12665 31803 12699
rect 36369 12665 36403 12699
rect 1685 12597 1719 12631
rect 2145 12597 2179 12631
rect 2789 12597 2823 12631
rect 3341 12597 3375 12631
rect 10885 12597 10919 12631
rect 13185 12597 13219 12631
rect 14657 12597 14691 12631
rect 16037 12597 16071 12631
rect 16957 12597 16991 12631
rect 20545 12597 20579 12631
rect 21281 12597 21315 12631
rect 22017 12597 22051 12631
rect 22569 12597 22603 12631
rect 25881 12597 25915 12631
rect 26525 12597 26559 12631
rect 27445 12597 27479 12631
rect 28089 12597 28123 12631
rect 32413 12597 32447 12631
rect 32505 12597 32539 12631
rect 33425 12597 33459 12631
rect 34253 12597 34287 12631
rect 35265 12597 35299 12631
rect 36737 12597 36771 12631
rect 5365 12393 5399 12427
rect 6469 12393 6503 12427
rect 7573 12393 7607 12427
rect 25421 12393 25455 12427
rect 28273 12393 28307 12427
rect 30389 12393 30423 12427
rect 31125 12393 31159 12427
rect 31585 12393 31619 12427
rect 32873 12393 32907 12427
rect 2697 12325 2731 12359
rect 12541 12325 12575 12359
rect 13829 12325 13863 12359
rect 16957 12325 16991 12359
rect 18245 12325 18279 12359
rect 19809 12325 19843 12359
rect 21741 12325 21775 12359
rect 23305 12325 23339 12359
rect 25237 12325 25271 12359
rect 28365 12325 28399 12359
rect 28825 12325 28859 12359
rect 29837 12325 29871 12359
rect 34069 12325 34103 12359
rect 4077 12257 4111 12291
rect 5181 12257 5215 12291
rect 6285 12257 6319 12291
rect 7389 12257 7423 12291
rect 12357 12257 12391 12291
rect 13553 12257 13587 12291
rect 17969 12257 18003 12291
rect 18797 12257 18831 12291
rect 19533 12257 19567 12291
rect 21557 12257 21591 12291
rect 23121 12257 23155 12291
rect 25513 12257 25547 12291
rect 30665 12257 30699 12291
rect 30941 12257 30975 12291
rect 32689 12257 32723 12291
rect 33793 12257 33827 12291
rect 35449 12257 35483 12291
rect 36553 12257 36587 12291
rect 2697 12189 2731 12223
rect 2789 12189 2823 12223
rect 3249 12189 3283 12223
rect 4629 12189 4663 12223
rect 12633 12189 12667 12223
rect 16865 12189 16899 12223
rect 17049 12189 17083 12223
rect 21833 12189 21867 12223
rect 23397 12189 23431 12223
rect 26985 12189 27019 12223
rect 28273 12189 28307 12223
rect 29101 12189 29135 12223
rect 29837 12189 29871 12223
rect 29929 12189 29963 12223
rect 1869 12121 1903 12155
rect 4261 12121 4295 12155
rect 16497 12121 16531 12155
rect 24041 12121 24075 12155
rect 24685 12121 24719 12155
rect 24961 12121 24995 12155
rect 27629 12121 27663 12155
rect 29377 12121 29411 12155
rect 2237 12053 2271 12087
rect 3617 12053 3651 12087
rect 6837 12053 6871 12087
rect 9229 12053 9263 12087
rect 12081 12053 12115 12087
rect 13001 12053 13035 12087
rect 14933 12053 14967 12087
rect 16221 12053 16255 12087
rect 20729 12053 20763 12087
rect 21281 12053 21315 12087
rect 22845 12053 22879 12087
rect 24409 12053 24443 12087
rect 25973 12053 26007 12087
rect 27813 12053 27847 12087
rect 33333 12053 33367 12087
rect 33701 12053 33735 12087
rect 35633 12053 35667 12087
rect 36737 12053 36771 12087
rect 5457 11849 5491 11883
rect 5825 11849 5859 11883
rect 12081 11849 12115 11883
rect 13921 11849 13955 11883
rect 14749 11849 14783 11883
rect 19625 11849 19659 11883
rect 20913 11849 20947 11883
rect 21833 11849 21867 11883
rect 23305 11849 23339 11883
rect 29469 11849 29503 11883
rect 31769 11849 31803 11883
rect 33241 11849 33275 11883
rect 34161 11849 34195 11883
rect 1593 11781 1627 11815
rect 2605 11781 2639 11815
rect 4169 11781 4203 11815
rect 9229 11781 9263 11815
rect 12541 11781 12575 11815
rect 14933 11781 14967 11815
rect 16497 11781 16531 11815
rect 18153 11781 18187 11815
rect 20361 11781 20395 11815
rect 24041 11781 24075 11815
rect 26893 11781 26927 11815
rect 29101 11781 29135 11815
rect 3985 11713 4019 11747
rect 4537 11713 4571 11747
rect 6285 11713 6319 11747
rect 7113 11713 7147 11747
rect 9781 11713 9815 11747
rect 11713 11713 11747 11747
rect 12909 11713 12943 11747
rect 15393 11713 15427 11747
rect 16957 11713 16991 11747
rect 21281 11713 21315 11747
rect 22385 11713 22419 11747
rect 24593 11713 24627 11747
rect 28181 11713 28215 11747
rect 33701 11713 33735 11747
rect 1409 11645 1443 11679
rect 5181 11645 5215 11679
rect 5641 11645 5675 11679
rect 6837 11645 6871 11679
rect 17877 11645 17911 11679
rect 22937 11645 22971 11679
rect 24317 11645 24351 11679
rect 25513 11645 25547 11679
rect 29285 11645 29319 11679
rect 29837 11645 29871 11679
rect 30389 11645 30423 11679
rect 30656 11645 30690 11679
rect 35449 11645 35483 11679
rect 36001 11645 36035 11679
rect 36553 11645 36587 11679
rect 37105 11645 37139 11679
rect 2053 11577 2087 11611
rect 2881 11577 2915 11611
rect 3157 11577 3191 11611
rect 4629 11577 4663 11611
rect 4721 11577 4755 11611
rect 9505 11577 9539 11611
rect 9689 11577 9723 11611
rect 11345 11577 11379 11611
rect 13001 11577 13035 11611
rect 13093 11577 13127 11611
rect 15485 11577 15519 11611
rect 16957 11577 16991 11611
rect 17049 11577 17083 11611
rect 17509 11577 17543 11611
rect 18429 11577 18463 11611
rect 18613 11577 18647 11611
rect 18705 11577 18739 11611
rect 19073 11577 19107 11611
rect 19993 11577 20027 11611
rect 20729 11577 20763 11611
rect 21465 11577 21499 11611
rect 24501 11577 24535 11611
rect 25780 11577 25814 11611
rect 27813 11577 27847 11611
rect 33793 11577 33827 11611
rect 2421 11509 2455 11543
rect 3065 11509 3099 11543
rect 3525 11509 3559 11543
rect 6561 11509 6595 11543
rect 7665 11509 7699 11543
rect 8953 11509 8987 11543
rect 13461 11509 13495 11543
rect 15393 11509 15427 11543
rect 15945 11509 15979 11543
rect 16221 11509 16255 11543
rect 21373 11509 21407 11543
rect 22201 11509 22235 11543
rect 24961 11509 24995 11543
rect 25329 11509 25363 11543
rect 28733 11509 28767 11543
rect 30297 11509 30331 11543
rect 32413 11509 32447 11543
rect 32689 11509 32723 11543
rect 33701 11509 33735 11543
rect 34713 11509 34747 11543
rect 35265 11509 35299 11543
rect 35633 11509 35667 11543
rect 36461 11509 36495 11543
rect 36737 11509 36771 11543
rect 2605 11305 2639 11339
rect 3801 11305 3835 11339
rect 4629 11305 4663 11339
rect 9137 11305 9171 11339
rect 12081 11305 12115 11339
rect 15945 11305 15979 11339
rect 17049 11305 17083 11339
rect 20729 11305 20763 11339
rect 22753 11305 22787 11339
rect 25237 11305 25271 11339
rect 25789 11305 25823 11339
rect 26249 11305 26283 11339
rect 28457 11305 28491 11339
rect 28825 11305 28859 11339
rect 30757 11305 30791 11339
rect 31125 11305 31159 11339
rect 4721 11237 4755 11271
rect 10241 11237 10275 11271
rect 16589 11237 16623 11271
rect 17846 11237 17880 11271
rect 21281 11237 21315 11271
rect 26792 11237 26826 11271
rect 29561 11237 29595 11271
rect 32413 11237 32447 11271
rect 33425 11237 33459 11271
rect 35173 11237 35207 11271
rect 2421 11169 2455 11203
rect 3433 11169 3467 11203
rect 5089 11169 5123 11203
rect 5641 11169 5675 11203
rect 10057 11169 10091 11203
rect 12521 11169 12555 11203
rect 21640 11169 21674 11203
rect 24124 11169 24158 11203
rect 29377 11169 29411 11203
rect 30941 11169 30975 11203
rect 35265 11169 35299 11203
rect 35633 11169 35667 11203
rect 36185 11169 36219 11203
rect 1685 11101 1719 11135
rect 2697 11101 2731 11135
rect 2973 11101 3007 11135
rect 2145 11033 2179 11067
rect 3709 11101 3743 11135
rect 4629 11101 4663 11135
rect 8585 11101 8619 11135
rect 10333 11101 10367 11135
rect 12265 11101 12299 11135
rect 16497 11101 16531 11135
rect 16681 11101 16715 11135
rect 17601 11101 17635 11135
rect 21373 11101 21407 11135
rect 23857 11101 23891 11135
rect 26525 11101 26559 11135
rect 29653 11101 29687 11135
rect 32781 11101 32815 11135
rect 33333 11101 33367 11135
rect 33517 11101 33551 11135
rect 34529 11101 34563 11135
rect 35173 11101 35207 11135
rect 5825 11033 5859 11067
rect 9781 11033 9815 11067
rect 14933 11033 14967 11067
rect 16129 11033 16163 11067
rect 27905 11033 27939 11067
rect 29101 11033 29135 11067
rect 30389 11033 30423 11067
rect 32965 11033 32999 11067
rect 34713 11033 34747 11067
rect 36369 11033 36403 11067
rect 2973 10965 3007 10999
rect 3157 10965 3191 10999
rect 3709 10965 3743 10999
rect 4169 10965 4203 10999
rect 5457 10965 5491 10999
rect 6929 10965 6963 10999
rect 13645 10965 13679 10999
rect 18981 10965 19015 10999
rect 23305 10965 23339 10999
rect 23765 10965 23799 10999
rect 30021 10965 30055 10999
rect 33885 10965 33919 10999
rect 36829 10965 36863 10999
rect 2513 10761 2547 10795
rect 4077 10761 4111 10795
rect 5733 10761 5767 10795
rect 8769 10761 8803 10795
rect 10609 10761 10643 10795
rect 11253 10761 11287 10795
rect 11897 10761 11931 10795
rect 12541 10761 12575 10795
rect 16129 10761 16163 10795
rect 17141 10761 17175 10795
rect 18245 10761 18279 10795
rect 18705 10761 18739 10795
rect 21833 10761 21867 10795
rect 26617 10761 26651 10795
rect 30665 10761 30699 10795
rect 31677 10761 31711 10795
rect 33333 10761 33367 10795
rect 34713 10761 34747 10795
rect 36553 10761 36587 10795
rect 6929 10693 6963 10727
rect 23765 10693 23799 10727
rect 27169 10693 27203 10727
rect 32321 10693 32355 10727
rect 34989 10693 35023 10727
rect 1409 10625 1443 10659
rect 1961 10625 1995 10659
rect 2881 10625 2915 10659
rect 4537 10625 4571 10659
rect 13829 10625 13863 10659
rect 14013 10625 14047 10659
rect 16405 10625 16439 10659
rect 16681 10625 16715 10659
rect 22293 10625 22327 10659
rect 22385 10625 22419 10659
rect 22845 10625 22879 10659
rect 24317 10625 24351 10659
rect 33885 10625 33919 10659
rect 35357 10625 35391 10659
rect 36921 10625 36955 10659
rect 4629 10557 4663 10591
rect 4997 10557 5031 10591
rect 5549 10557 5583 10591
rect 7481 10557 7515 10591
rect 8953 10557 8987 10591
rect 9229 10557 9263 10591
rect 12817 10557 12851 10591
rect 19257 10557 19291 10591
rect 19513 10557 19547 10591
rect 23489 10557 23523 10591
rect 24685 10557 24719 10591
rect 25053 10557 25087 10591
rect 25237 10557 25271 10591
rect 29285 10557 29319 10591
rect 32137 10557 32171 10591
rect 32689 10557 32723 10591
rect 37473 10557 37507 10591
rect 2329 10489 2363 10523
rect 2973 10489 3007 10523
rect 3065 10489 3099 10523
rect 4537 10489 4571 10523
rect 7205 10489 7239 10523
rect 8401 10489 8435 10523
rect 9496 10489 9530 10523
rect 13093 10489 13127 10523
rect 13461 10489 13495 10523
rect 14258 10489 14292 10523
rect 22293 10489 22327 10523
rect 24041 10489 24075 10523
rect 25504 10489 25538 10523
rect 29530 10489 29564 10523
rect 33057 10489 33091 10523
rect 33609 10489 33643 10523
rect 35541 10489 35575 10523
rect 37013 10489 37047 10523
rect 37105 10489 37139 10523
rect 3433 10421 3467 10455
rect 3801 10421 3835 10455
rect 5457 10421 5491 10455
rect 6193 10421 6227 10455
rect 6561 10421 6595 10455
rect 7389 10421 7423 10455
rect 8953 10421 8987 10455
rect 9045 10421 9079 10455
rect 12173 10421 12207 10455
rect 13001 10421 13035 10455
rect 15393 10421 15427 10455
rect 17601 10421 17635 10455
rect 19073 10421 19107 10455
rect 20637 10421 20671 10455
rect 21373 10421 21407 10455
rect 24225 10421 24259 10455
rect 28365 10421 28399 10455
rect 28641 10421 28675 10455
rect 29009 10421 29043 10455
rect 31217 10421 31251 10455
rect 32045 10421 32079 10455
rect 33793 10421 33827 10455
rect 34345 10421 34379 10455
rect 35449 10421 35483 10455
rect 36185 10421 36219 10455
rect 2513 10217 2547 10251
rect 4353 10217 4387 10251
rect 5917 10217 5951 10251
rect 10241 10217 10275 10251
rect 12081 10217 12115 10251
rect 13001 10217 13035 10251
rect 16129 10217 16163 10251
rect 17785 10217 17819 10251
rect 20729 10217 20763 10251
rect 22661 10217 22695 10251
rect 24133 10217 24167 10251
rect 25237 10217 25271 10251
rect 26065 10217 26099 10251
rect 26985 10217 27019 10251
rect 29837 10217 29871 10251
rect 36553 10217 36587 10251
rect 37105 10217 37139 10251
rect 1869 10149 1903 10183
rect 2605 10149 2639 10183
rect 3433 10149 3467 10183
rect 4782 10149 4816 10183
rect 7266 10149 7300 10183
rect 12633 10149 12667 10183
rect 14197 10149 14231 10183
rect 19809 10149 19843 10183
rect 25697 10149 25731 10183
rect 28273 10149 28307 10183
rect 29359 10149 29393 10183
rect 32597 10149 32631 10183
rect 32956 10149 32990 10183
rect 35418 10149 35452 10183
rect 7021 10081 7055 10115
rect 10057 10081 10091 10115
rect 11437 10081 11471 10115
rect 13277 10081 13311 10115
rect 14289 10081 14323 10115
rect 16661 10081 16695 10115
rect 21189 10081 21223 10115
rect 21548 10081 21582 10115
rect 25053 10081 25087 10115
rect 25329 10081 25363 10115
rect 32689 10081 32723 10115
rect 2421 10013 2455 10047
rect 4537 10013 4571 10047
rect 9321 10013 9355 10047
rect 10333 10013 10367 10047
rect 12081 10013 12115 10047
rect 12173 10013 12207 10047
rect 14197 10013 14231 10047
rect 16405 10013 16439 10047
rect 19165 10013 19199 10047
rect 19809 10013 19843 10047
rect 19901 10013 19935 10047
rect 21281 10013 21315 10047
rect 23489 10013 23523 10047
rect 26525 10013 26559 10047
rect 28181 10013 28215 10047
rect 28365 10013 28399 10047
rect 29745 10013 29779 10047
rect 29929 10013 29963 10047
rect 35173 10013 35207 10047
rect 2053 9945 2087 9979
rect 9781 9945 9815 9979
rect 11621 9945 11655 9979
rect 13737 9945 13771 9979
rect 19349 9945 19383 9979
rect 24501 9945 24535 9979
rect 3065 9877 3099 9911
rect 3893 9877 3927 9911
rect 6469 9877 6503 9911
rect 6929 9877 6963 9911
rect 8401 9877 8435 9911
rect 10885 9877 10919 9911
rect 18797 9877 18831 9911
rect 20361 9877 20395 9911
rect 23857 9877 23891 9911
rect 24777 9877 24811 9911
rect 27813 9877 27847 9911
rect 29193 9877 29227 9911
rect 30389 9877 30423 9911
rect 34069 9877 34103 9911
rect 34989 9877 35023 9911
rect 4261 9673 4295 9707
rect 5181 9673 5215 9707
rect 6561 9673 6595 9707
rect 10057 9673 10091 9707
rect 14381 9673 14415 9707
rect 15117 9673 15151 9707
rect 17233 9673 17267 9707
rect 17601 9673 17635 9707
rect 25145 9673 25179 9707
rect 33057 9673 33091 9707
rect 5549 9605 5583 9639
rect 9781 9605 9815 9639
rect 10885 9605 10919 9639
rect 13829 9605 13863 9639
rect 14841 9605 14875 9639
rect 18797 9605 18831 9639
rect 20361 9605 20395 9639
rect 21925 9605 21959 9639
rect 23857 9605 23891 9639
rect 26709 9605 26743 9639
rect 27445 9605 27479 9639
rect 28641 9605 28675 9639
rect 33333 9605 33367 9639
rect 34989 9605 35023 9639
rect 35909 9605 35943 9639
rect 1869 9537 1903 9571
rect 2881 9537 2915 9571
rect 7021 9537 7055 9571
rect 7481 9537 7515 9571
rect 7665 9537 7699 9571
rect 11437 9537 11471 9571
rect 11897 9537 11931 9571
rect 19349 9537 19383 9571
rect 19809 9537 19843 9571
rect 20085 9537 20119 9571
rect 22477 9537 22511 9571
rect 23489 9537 23523 9571
rect 24317 9537 24351 9571
rect 29101 9537 29135 9571
rect 29561 9537 29595 9571
rect 32045 9537 32079 9571
rect 37565 9537 37599 9571
rect 1593 9469 1627 9503
rect 3148 9469 3182 9503
rect 4813 9469 4847 9503
rect 5365 9469 5399 9503
rect 7932 9469 7966 9503
rect 12173 9469 12207 9503
rect 12449 9469 12483 9503
rect 15301 9469 15335 9503
rect 15557 9469 15591 9503
rect 20913 9469 20947 9503
rect 23121 9469 23155 9503
rect 24409 9469 24443 9503
rect 25329 9469 25363 9503
rect 25596 9469 25630 9503
rect 29828 9469 29862 9503
rect 32137 9469 32171 9503
rect 35541 9469 35575 9503
rect 36277 9469 36311 9503
rect 36461 9469 36495 9503
rect 37013 9469 37047 9503
rect 2421 9401 2455 9435
rect 11161 9401 11195 9435
rect 12716 9401 12750 9435
rect 19073 9401 19107 9435
rect 20637 9401 20671 9435
rect 22201 9401 22235 9435
rect 24317 9401 24351 9435
rect 28089 9401 28123 9435
rect 33609 9401 33643 9435
rect 33885 9401 33919 9435
rect 35265 9401 35299 9435
rect 35449 9401 35483 9435
rect 2697 9333 2731 9367
rect 6009 9333 6043 9367
rect 9045 9333 9079 9367
rect 10609 9333 10643 9367
rect 11345 9333 11379 9367
rect 16681 9333 16715 9367
rect 18521 9333 18555 9367
rect 19257 9333 19291 9367
rect 20821 9333 20855 9367
rect 21281 9333 21315 9367
rect 21741 9333 21775 9367
rect 22385 9333 22419 9367
rect 24869 9333 24903 9367
rect 27721 9333 27755 9367
rect 30941 9333 30975 9367
rect 32321 9333 32355 9367
rect 32781 9333 32815 9367
rect 33793 9333 33827 9367
rect 34345 9333 34379 9367
rect 34621 9333 34655 9367
rect 36645 9333 36679 9367
rect 4261 9129 4295 9163
rect 4629 9129 4663 9163
rect 4997 9129 5031 9163
rect 8217 9129 8251 9163
rect 9505 9129 9539 9163
rect 11345 9129 11379 9163
rect 14105 9129 14139 9163
rect 17877 9129 17911 9163
rect 19165 9129 19199 9163
rect 20637 9129 20671 9163
rect 22293 9129 22327 9163
rect 25605 9129 25639 9163
rect 27169 9129 27203 9163
rect 27721 9129 27755 9163
rect 30941 9129 30975 9163
rect 36461 9129 36495 9163
rect 1961 9061 1995 9095
rect 3065 9061 3099 9095
rect 6101 9061 6135 9095
rect 7665 9061 7699 9095
rect 7757 9061 7791 9095
rect 10241 9061 10275 9095
rect 11693 9061 11727 9095
rect 19809 9061 19843 9095
rect 21281 9061 21315 9095
rect 21465 9061 21499 9095
rect 22845 9061 22879 9095
rect 23489 9061 23523 9095
rect 24575 9061 24609 9095
rect 25053 9061 25087 9095
rect 26065 9061 26099 9095
rect 28089 9061 28123 9095
rect 33149 9061 33183 9095
rect 1961 8925 1995 8959
rect 2053 8925 2087 8959
rect 2421 8925 2455 8959
rect 1501 8857 1535 8891
rect 2881 8857 2915 8891
rect 3525 8993 3559 9027
rect 4077 8993 4111 9027
rect 5457 8993 5491 9027
rect 6193 8993 6227 9027
rect 6929 8993 6963 9027
rect 8585 8993 8619 9027
rect 10333 8993 10367 9027
rect 10885 8993 10919 9027
rect 16764 8993 16798 9027
rect 19625 8993 19659 9027
rect 21557 8993 21591 9027
rect 23305 8993 23339 9027
rect 26985 8993 27019 9027
rect 28365 8993 28399 9027
rect 29817 8993 29851 9027
rect 32505 8993 32539 9027
rect 32965 8993 32999 9027
rect 34428 8993 34462 9027
rect 6101 8925 6135 8959
rect 7665 8925 7699 8959
rect 10241 8925 10275 8959
rect 11437 8925 11471 8959
rect 16497 8925 16531 8959
rect 19901 8925 19935 8959
rect 23581 8925 23615 8959
rect 24961 8925 24995 8959
rect 25145 8925 25179 8959
rect 27261 8925 27295 8959
rect 29561 8925 29595 8959
rect 33241 8925 33275 8959
rect 34161 8925 34195 8959
rect 36645 8925 36679 8959
rect 5641 8857 5675 8891
rect 19349 8857 19383 8891
rect 23029 8857 23063 8891
rect 35541 8857 35575 8891
rect 36093 8857 36127 8891
rect 3065 8789 3099 8823
rect 3249 8789 3283 8823
rect 6653 8789 6687 8823
rect 7205 8789 7239 8823
rect 9781 8789 9815 8823
rect 12817 8789 12851 8823
rect 13737 8789 13771 8823
rect 18797 8789 18831 8823
rect 20361 8789 20395 8823
rect 21005 8789 21039 8823
rect 21925 8789 21959 8823
rect 24225 8789 24259 8823
rect 26709 8789 26743 8823
rect 28917 8789 28951 8823
rect 29377 8789 29411 8823
rect 32689 8789 32723 8823
rect 33609 8789 33643 8823
rect 34069 8789 34103 8823
rect 2053 8585 2087 8619
rect 3985 8585 4019 8619
rect 4629 8585 4663 8619
rect 5089 8585 5123 8619
rect 6285 8585 6319 8619
rect 7021 8585 7055 8619
rect 8401 8585 8435 8619
rect 10977 8585 11011 8619
rect 11437 8585 11471 8619
rect 12173 8585 12207 8619
rect 13921 8585 13955 8619
rect 16773 8585 16807 8619
rect 18705 8585 18739 8619
rect 19073 8585 19107 8619
rect 19349 8585 19383 8619
rect 23489 8585 23523 8619
rect 24317 8585 24351 8619
rect 25237 8585 25271 8619
rect 26157 8585 26191 8619
rect 27721 8585 27755 8619
rect 30297 8585 30331 8619
rect 33701 8585 33735 8619
rect 35909 8585 35943 8619
rect 1593 8517 1627 8551
rect 5273 8517 5307 8551
rect 7941 8517 7975 8551
rect 9965 8517 9999 8551
rect 11805 8517 11839 8551
rect 28733 8517 28767 8551
rect 29377 8517 29411 8551
rect 34989 8517 35023 8551
rect 5733 8449 5767 8483
rect 6653 8449 6687 8483
rect 7481 8449 7515 8483
rect 8585 8449 8619 8483
rect 13369 8449 13403 8483
rect 14473 8449 14507 8483
rect 15393 8449 15427 8483
rect 19901 8449 19935 8483
rect 24869 8449 24903 8483
rect 26525 8449 26559 8483
rect 26709 8449 26743 8483
rect 28181 8449 28215 8483
rect 29101 8449 29135 8483
rect 29929 8449 29963 8483
rect 31309 8449 31343 8483
rect 35449 8449 35483 8483
rect 36737 8449 36771 8483
rect 1409 8381 1443 8415
rect 2605 8381 2639 8415
rect 7573 8381 7607 8415
rect 13737 8381 13771 8415
rect 20821 8381 20855 8415
rect 27169 8381 27203 8415
rect 27537 8381 27571 8415
rect 31033 8381 31067 8415
rect 32229 8381 32263 8415
rect 32321 8381 32355 8415
rect 34345 8381 34379 8415
rect 36277 8381 36311 8415
rect 36461 8381 36495 8415
rect 37197 8381 37231 8415
rect 2872 8313 2906 8347
rect 5733 8313 5767 8347
rect 5825 8313 5859 8347
rect 8830 8313 8864 8347
rect 10517 8313 10551 8347
rect 14197 8313 14231 8347
rect 14381 8313 14415 8347
rect 14933 8313 14967 8347
rect 15660 8313 15694 8347
rect 18061 8313 18095 8347
rect 19625 8313 19659 8347
rect 19809 8313 19843 8347
rect 20361 8313 20395 8347
rect 21088 8313 21122 8347
rect 24041 8313 24075 8347
rect 24593 8313 24627 8347
rect 25973 8313 26007 8347
rect 26617 8313 26651 8347
rect 28181 8313 28215 8347
rect 28273 8313 28307 8347
rect 29653 8313 29687 8347
rect 29837 8313 29871 8347
rect 31861 8313 31895 8347
rect 32588 8313 32622 8347
rect 34713 8313 34747 8347
rect 35449 8313 35483 8347
rect 35541 8313 35575 8347
rect 2421 8245 2455 8279
rect 7481 8245 7515 8279
rect 12725 8245 12759 8279
rect 15209 8245 15243 8279
rect 17325 8245 17359 8279
rect 20729 8245 20763 8279
rect 22201 8245 22235 8279
rect 22937 8245 22971 8279
rect 24777 8245 24811 8279
rect 30941 8245 30975 8279
rect 3801 8041 3835 8075
rect 4261 8041 4295 8075
rect 4905 8041 4939 8075
rect 6377 8041 6411 8075
rect 8033 8041 8067 8075
rect 9413 8041 9447 8075
rect 10241 8041 10275 8075
rect 16313 8041 16347 8075
rect 17141 8041 17175 8075
rect 18705 8041 18739 8075
rect 19993 8041 20027 8075
rect 20913 8041 20947 8075
rect 21465 8041 21499 8075
rect 22109 8041 22143 8075
rect 24685 8041 24719 8075
rect 26157 8041 26191 8075
rect 27997 8041 28031 8075
rect 30665 8041 30699 8075
rect 34897 8041 34931 8075
rect 36461 8041 36495 8075
rect 36829 8041 36863 8075
rect 2973 7973 3007 8007
rect 5181 7973 5215 8007
rect 5917 7973 5951 8007
rect 6745 7973 6779 8007
rect 7481 7973 7515 8007
rect 8493 7973 8527 8007
rect 11774 7973 11808 8007
rect 19717 7973 19751 8007
rect 25329 7973 25363 8007
rect 27077 7973 27111 8007
rect 29000 7973 29034 8007
rect 32781 7973 32815 8007
rect 33232 7973 33266 8007
rect 36001 7973 36035 8007
rect 3433 7905 3467 7939
rect 4077 7905 4111 7939
rect 8309 7905 8343 7939
rect 11529 7905 11563 7939
rect 15669 7905 15703 7939
rect 16405 7905 16439 7939
rect 16773 7905 16807 7939
rect 17592 7905 17626 7939
rect 20729 7905 20763 7939
rect 21833 7905 21867 7939
rect 22560 7905 22594 7939
rect 25145 7905 25179 7939
rect 28733 7905 28767 7939
rect 32965 7905 32999 7939
rect 1409 7837 1443 7871
rect 2237 7837 2271 7871
rect 2881 7837 2915 7871
rect 3065 7837 3099 7871
rect 5917 7837 5951 7871
rect 6009 7837 6043 7871
rect 7389 7837 7423 7871
rect 7573 7837 7607 7871
rect 10241 7837 10275 7871
rect 10333 7837 10367 7871
rect 16313 7837 16347 7871
rect 17325 7837 17359 7871
rect 22293 7837 22327 7871
rect 25421 7837 25455 7871
rect 26985 7837 27019 7871
rect 27169 7837 27203 7871
rect 36001 7837 36035 7871
rect 36093 7837 36127 7871
rect 5457 7769 5491 7803
rect 7021 7769 7055 7803
rect 11345 7769 11379 7803
rect 24869 7769 24903 7803
rect 27537 7769 27571 7803
rect 32413 7769 32447 7803
rect 35541 7769 35575 7803
rect 1869 7701 1903 7735
rect 2513 7701 2547 7735
rect 9781 7701 9815 7735
rect 10793 7701 10827 7735
rect 12909 7701 12943 7735
rect 13921 7701 13955 7735
rect 15853 7701 15887 7735
rect 19349 7701 19383 7735
rect 23673 7701 23707 7735
rect 24317 7701 24351 7735
rect 26617 7701 26651 7735
rect 28641 7701 28675 7735
rect 30113 7701 30147 7735
rect 34345 7701 34379 7735
rect 35265 7701 35299 7735
rect 3157 7497 3191 7531
rect 4169 7497 4203 7531
rect 6193 7497 6227 7531
rect 7113 7497 7147 7531
rect 10149 7497 10183 7531
rect 15117 7497 15151 7531
rect 20913 7497 20947 7531
rect 23489 7497 23523 7531
rect 25973 7497 26007 7531
rect 28089 7497 28123 7531
rect 28733 7497 28767 7531
rect 29009 7497 29043 7531
rect 32229 7497 32263 7531
rect 33701 7497 33735 7531
rect 36553 7497 36587 7531
rect 6653 7429 6687 7463
rect 10701 7429 10735 7463
rect 11621 7429 11655 7463
rect 12173 7429 12207 7463
rect 15761 7429 15795 7463
rect 16221 7429 16255 7463
rect 17141 7429 17175 7463
rect 19625 7429 19659 7463
rect 27169 7429 27203 7463
rect 34989 7429 35023 7463
rect 36001 7429 36035 7463
rect 16589 7361 16623 7395
rect 16773 7361 16807 7395
rect 19441 7361 19475 7395
rect 20085 7361 20119 7395
rect 21097 7361 21131 7395
rect 29285 7361 29319 7395
rect 32321 7361 32355 7395
rect 37105 7361 37139 7395
rect 1777 7293 1811 7327
rect 2044 7293 2078 7327
rect 4261 7293 4295 7327
rect 7481 7293 7515 7327
rect 11253 7293 11287 7327
rect 12449 7293 12483 7327
rect 15485 7293 15519 7327
rect 19073 7293 19107 7327
rect 24593 7293 24627 7327
rect 24860 7293 24894 7327
rect 29552 7293 29586 7327
rect 35265 7293 35299 7327
rect 36829 7293 36863 7327
rect 1685 7225 1719 7259
rect 4528 7225 4562 7259
rect 7748 7225 7782 7259
rect 10977 7225 11011 7259
rect 11161 7225 11195 7259
rect 12694 7225 12728 7259
rect 16681 7225 16715 7259
rect 18705 7225 18739 7259
rect 20177 7225 20211 7259
rect 21342 7225 21376 7259
rect 24133 7225 24167 7259
rect 26617 7225 26651 7259
rect 27445 7225 27479 7259
rect 27721 7225 27755 7259
rect 31861 7225 31895 7259
rect 32566 7225 32600 7259
rect 35541 7225 35575 7259
rect 37013 7225 37047 7259
rect 3801 7157 3835 7191
rect 5641 7157 5675 7191
rect 8861 7157 8895 7191
rect 9781 7157 9815 7191
rect 10425 7157 10459 7191
rect 13829 7157 13863 7191
rect 17601 7157 17635 7191
rect 20085 7157 20119 7191
rect 22477 7157 22511 7191
rect 23121 7157 23155 7191
rect 24501 7157 24535 7191
rect 26893 7157 26927 7191
rect 27629 7157 27663 7191
rect 30665 7157 30699 7191
rect 34345 7157 34379 7191
rect 34713 7157 34747 7191
rect 35449 7157 35483 7191
rect 36369 7157 36403 7191
rect 2881 6953 2915 6987
rect 3801 6953 3835 6987
rect 6745 6953 6779 6987
rect 7941 6953 7975 6987
rect 10241 6953 10275 6987
rect 11897 6953 11931 6987
rect 17141 6953 17175 6987
rect 21189 6953 21223 6987
rect 23673 6953 23707 6987
rect 24685 6953 24719 6987
rect 25973 6953 26007 6987
rect 27077 6953 27111 6987
rect 28089 6953 28123 6987
rect 32321 6953 32355 6987
rect 33793 6953 33827 6987
rect 5917 6885 5951 6919
rect 7297 6885 7331 6919
rect 7481 6885 7515 6919
rect 10057 6885 10091 6919
rect 13461 6885 13495 6919
rect 25421 6885 25455 6919
rect 33333 6885 33367 6919
rect 33425 6885 33459 6919
rect 34897 6885 34931 6919
rect 36461 6885 36495 6919
rect 1501 6817 1535 6851
rect 1768 6817 1802 6851
rect 4077 6817 4111 6851
rect 5733 6817 5767 6851
rect 8493 6817 8527 6851
rect 8953 6817 8987 6851
rect 10701 6817 10735 6851
rect 11713 6817 11747 6851
rect 16028 6817 16062 6851
rect 18501 6817 18535 6851
rect 22293 6817 22327 6851
rect 22549 6817 22583 6851
rect 24225 6817 24259 6851
rect 26893 6817 26927 6851
rect 28825 6817 28859 6851
rect 29357 6817 29391 6851
rect 34989 6817 35023 6851
rect 35725 6817 35759 6851
rect 36553 6817 36587 6851
rect 4721 6749 4755 6783
rect 5273 6749 5307 6783
rect 6009 6749 6043 6783
rect 6377 6749 6411 6783
rect 7573 6749 7607 6783
rect 8309 6749 8343 6783
rect 9413 6749 9447 6783
rect 10333 6749 10367 6783
rect 11989 6749 12023 6783
rect 13369 6749 13403 6783
rect 13553 6749 13587 6783
rect 15761 6749 15795 6783
rect 18245 6749 18279 6783
rect 25421 6749 25455 6783
rect 25513 6749 25547 6783
rect 27169 6749 27203 6783
rect 27537 6749 27571 6783
rect 29101 6749 29135 6783
rect 33333 6749 33367 6783
rect 34897 6749 34931 6783
rect 36369 6749 36403 6783
rect 4261 6681 4295 6715
rect 7021 6681 7055 6715
rect 11437 6681 11471 6715
rect 13001 6681 13035 6715
rect 24961 6681 24995 6715
rect 26249 6681 26283 6715
rect 32873 6681 32907 6715
rect 3525 6613 3559 6647
rect 5457 6613 5491 6647
rect 9781 6613 9815 6647
rect 11161 6613 11195 6647
rect 12633 6613 12667 6647
rect 15485 6613 15519 6647
rect 17785 6613 17819 6647
rect 18061 6613 18095 6647
rect 19625 6613 19659 6647
rect 26617 6613 26651 6647
rect 27905 6613 27939 6647
rect 30481 6613 30515 6647
rect 34437 6613 34471 6647
rect 35357 6613 35391 6647
rect 36001 6613 36035 6647
rect 36921 6613 36955 6647
rect 1593 6409 1627 6443
rect 2053 6409 2087 6443
rect 4537 6409 4571 6443
rect 5089 6409 5123 6443
rect 6285 6409 6319 6443
rect 6653 6409 6687 6443
rect 9413 6409 9447 6443
rect 10149 6409 10183 6443
rect 11805 6409 11839 6443
rect 12173 6409 12207 6443
rect 14565 6409 14599 6443
rect 17417 6409 17451 6443
rect 19073 6409 19107 6443
rect 21005 6409 21039 6443
rect 22477 6409 22511 6443
rect 23121 6409 23155 6443
rect 23949 6409 23983 6443
rect 24133 6409 24167 6443
rect 25145 6409 25179 6443
rect 27537 6409 27571 6443
rect 29009 6409 29043 6443
rect 33333 6409 33367 6443
rect 34069 6409 34103 6443
rect 36645 6409 36679 6443
rect 5273 6341 5307 6375
rect 10885 6341 10919 6375
rect 14013 6341 14047 6375
rect 18153 6341 18187 6375
rect 27905 6341 27939 6375
rect 29377 6341 29411 6375
rect 33057 6341 33091 6375
rect 5733 6273 5767 6307
rect 9781 6273 9815 6307
rect 11345 6273 11379 6307
rect 12633 6273 12667 6307
rect 21097 6273 21131 6307
rect 24501 6273 24535 6307
rect 24685 6273 24719 6307
rect 25421 6273 25455 6307
rect 29837 6273 29871 6307
rect 34345 6273 34379 6307
rect 35081 6273 35115 6307
rect 1409 6205 1443 6239
rect 2421 6205 2455 6239
rect 2605 6205 2639 6239
rect 5825 6205 5859 6239
rect 6837 6205 6871 6239
rect 8769 6205 8803 6239
rect 10701 6205 10735 6239
rect 11437 6205 11471 6239
rect 14933 6205 14967 6239
rect 15117 6205 15151 6239
rect 15373 6205 15407 6239
rect 19441 6205 19475 6239
rect 23489 6205 23523 6239
rect 25605 6205 25639 6239
rect 28733 6205 28767 6239
rect 29929 6205 29963 6239
rect 30941 6205 30975 6239
rect 31033 6205 31067 6239
rect 35265 6205 35299 6239
rect 35532 6205 35566 6239
rect 37197 6205 37231 6239
rect 2872 6137 2906 6171
rect 5733 6137 5767 6171
rect 7082 6137 7116 6171
rect 11345 6137 11379 6171
rect 12900 6137 12934 6171
rect 18429 6137 18463 6171
rect 18613 6137 18647 6171
rect 18705 6137 18739 6171
rect 20637 6137 20671 6171
rect 21342 6137 21376 6171
rect 24593 6137 24627 6171
rect 25872 6137 25906 6171
rect 28181 6137 28215 6171
rect 31278 6137 31312 6171
rect 3985 6069 4019 6103
rect 8217 6069 8251 6103
rect 16497 6069 16531 6103
rect 17049 6069 17083 6103
rect 17785 6069 17819 6103
rect 26985 6069 27019 6103
rect 29837 6069 29871 6103
rect 30297 6069 30331 6103
rect 32413 6069 32447 6103
rect 4261 5865 4295 5899
rect 5457 5865 5491 5899
rect 6101 5865 6135 5899
rect 7021 5865 7055 5899
rect 10057 5865 10091 5899
rect 11971 5865 12005 5899
rect 12449 5865 12483 5899
rect 13001 5865 13035 5899
rect 13369 5865 13403 5899
rect 15761 5865 15795 5899
rect 16681 5865 16715 5899
rect 21649 5865 21683 5899
rect 22385 5865 22419 5899
rect 24869 5865 24903 5899
rect 26801 5865 26835 5899
rect 27445 5865 27479 5899
rect 28539 5865 28573 5899
rect 29837 5865 29871 5899
rect 30573 5865 30607 5899
rect 33149 5865 33183 5899
rect 35541 5865 35575 5899
rect 36093 5865 36127 5899
rect 2789 5797 2823 5831
rect 3617 5797 3651 5831
rect 4629 5797 4663 5831
rect 7380 5797 7414 5831
rect 10701 5797 10735 5831
rect 10793 5797 10827 5831
rect 12265 5797 12299 5831
rect 12541 5797 12575 5831
rect 14013 5797 14047 5831
rect 14197 5797 14231 5831
rect 14289 5797 14323 5831
rect 16773 5797 16807 5831
rect 18061 5797 18095 5831
rect 18245 5797 18279 5831
rect 21741 5797 21775 5831
rect 29009 5797 29043 5831
rect 29469 5797 29503 5831
rect 32505 5797 32539 5831
rect 32965 5797 32999 5831
rect 33241 5797 33275 5831
rect 33701 5797 33735 5831
rect 34406 5797 34440 5831
rect 2605 5729 2639 5763
rect 4077 5729 4111 5763
rect 6193 5729 6227 5763
rect 6561 5729 6595 5763
rect 10517 5729 10551 5763
rect 11437 5729 11471 5763
rect 20729 5729 20763 5763
rect 22661 5729 22695 5763
rect 22928 5729 22962 5763
rect 27537 5729 27571 5763
rect 27905 5729 27939 5763
rect 28825 5729 28859 5763
rect 30665 5729 30699 5763
rect 31033 5729 31067 5763
rect 2881 5661 2915 5695
rect 6009 5661 6043 5695
rect 7113 5661 7147 5695
rect 16681 5661 16715 5695
rect 18337 5661 18371 5695
rect 19809 5661 19843 5695
rect 21557 5661 21591 5695
rect 25237 5661 25271 5695
rect 27445 5661 27479 5695
rect 29101 5661 29135 5695
rect 30481 5661 30515 5695
rect 34161 5661 34195 5695
rect 5641 5593 5675 5627
rect 13737 5593 13771 5627
rect 21189 5593 21223 5627
rect 26065 5593 26099 5627
rect 26985 5593 27019 5627
rect 32689 5593 32723 5627
rect 36461 5593 36495 5627
rect 1685 5525 1719 5559
rect 2145 5525 2179 5559
rect 2329 5525 2363 5559
rect 3249 5525 3283 5559
rect 4997 5525 5031 5559
rect 8493 5525 8527 5559
rect 10241 5525 10275 5559
rect 16221 5525 16255 5559
rect 17785 5525 17819 5559
rect 18705 5525 18739 5559
rect 24041 5525 24075 5559
rect 25697 5525 25731 5559
rect 30113 5525 30147 5559
rect 1593 5321 1627 5355
rect 2329 5321 2363 5355
rect 2881 5321 2915 5355
rect 4445 5321 4479 5355
rect 5641 5321 5675 5355
rect 6561 5321 6595 5355
rect 10885 5321 10919 5355
rect 11989 5321 12023 5355
rect 12909 5321 12943 5355
rect 13737 5321 13771 5355
rect 14105 5321 14139 5355
rect 15761 5321 15795 5355
rect 17049 5321 17083 5355
rect 17417 5321 17451 5355
rect 17785 5321 17819 5355
rect 19533 5321 19567 5355
rect 20821 5321 20855 5355
rect 21097 5321 21131 5355
rect 22385 5321 22419 5355
rect 22753 5321 22787 5355
rect 24685 5321 24719 5355
rect 25605 5321 25639 5355
rect 26617 5321 26651 5355
rect 28181 5321 28215 5355
rect 30941 5321 30975 5355
rect 31861 5321 31895 5355
rect 35633 5321 35667 5355
rect 6193 5253 6227 5287
rect 7389 5253 7423 5287
rect 8953 5253 8987 5287
rect 10241 5253 10275 5287
rect 14381 5253 14415 5287
rect 15577 5253 15611 5287
rect 18153 5253 18187 5287
rect 19809 5253 19843 5287
rect 21373 5253 21407 5287
rect 23765 5253 23799 5287
rect 26801 5253 26835 5287
rect 26893 5253 26927 5287
rect 27169 5253 27203 5287
rect 29653 5253 29687 5287
rect 4997 5185 5031 5219
rect 7757 5185 7791 5219
rect 10701 5185 10735 5219
rect 11437 5185 11471 5219
rect 12449 5185 12483 5219
rect 14841 5185 14875 5219
rect 16129 5185 16163 5219
rect 16773 5185 16807 5219
rect 18521 5185 18555 5219
rect 24225 5185 24259 5219
rect 26065 5185 26099 5219
rect 1409 5117 1443 5151
rect 3157 5117 3191 5151
rect 4169 5117 4203 5151
rect 9505 5117 9539 5151
rect 11161 5117 11195 5151
rect 15209 5117 15243 5151
rect 19257 5117 19291 5151
rect 20085 5117 20119 5151
rect 20361 5117 20395 5151
rect 21649 5117 21683 5151
rect 23489 5117 23523 5151
rect 3433 5049 3467 5083
rect 4721 5049 4755 5083
rect 7941 5049 7975 5083
rect 8309 5049 8343 5083
rect 9229 5049 9263 5083
rect 9413 5049 9447 5083
rect 16221 5049 16255 5083
rect 16313 5049 16347 5083
rect 18613 5049 18647 5083
rect 18705 5049 18739 5083
rect 21925 5049 21959 5083
rect 24317 5049 24351 5083
rect 26065 5049 26099 5083
rect 26157 5049 26191 5083
rect 27721 5185 27755 5219
rect 30205 5185 30239 5219
rect 28825 5117 28859 5151
rect 31309 5117 31343 5151
rect 32229 5117 32263 5151
rect 32321 5117 32355 5151
rect 32577 5117 32611 5151
rect 35449 5117 35483 5151
rect 36001 5117 36035 5151
rect 27445 5049 27479 5083
rect 28457 5049 28491 5083
rect 29929 5049 29963 5083
rect 30113 5049 30147 5083
rect 34621 5049 34655 5083
rect 2697 4981 2731 5015
rect 3341 4981 3375 5015
rect 4905 4981 4939 5015
rect 7113 4981 7147 5015
rect 7849 4981 7883 5015
rect 8769 4981 8803 5015
rect 11345 4981 11379 5015
rect 20269 4981 20303 5015
rect 21833 4981 21867 5015
rect 23121 4981 23155 5015
rect 24225 4981 24259 5015
rect 25421 4981 25455 5015
rect 26801 4981 26835 5015
rect 27629 4981 27663 5015
rect 30573 4981 30607 5015
rect 33701 4981 33735 5015
rect 34345 4981 34379 5015
rect 1685 4777 1719 4811
rect 2145 4777 2179 4811
rect 3893 4777 3927 4811
rect 6009 4777 6043 4811
rect 7757 4777 7791 4811
rect 10885 4777 10919 4811
rect 11253 4777 11287 4811
rect 11989 4777 12023 4811
rect 15761 4777 15795 4811
rect 16405 4777 16439 4811
rect 17785 4777 17819 4811
rect 18153 4777 18187 4811
rect 19809 4777 19843 4811
rect 20729 4777 20763 4811
rect 23765 4777 23799 4811
rect 25697 4777 25731 4811
rect 25881 4777 25915 4811
rect 28641 4777 28675 4811
rect 29653 4777 29687 4811
rect 30297 4777 30331 4811
rect 30757 4777 30791 4811
rect 32321 4777 32355 4811
rect 32781 4777 32815 4811
rect 33425 4777 33459 4811
rect 2881 4709 2915 4743
rect 7573 4709 7607 4743
rect 18429 4709 18463 4743
rect 21465 4709 21499 4743
rect 23581 4709 23615 4743
rect 25329 4709 25363 4743
rect 25421 4709 25455 4743
rect 26801 4709 26835 4743
rect 27528 4709 27562 4743
rect 30389 4709 30423 4743
rect 33241 4709 33275 4743
rect 3433 4641 3467 4675
rect 4344 4641 4378 4675
rect 12357 4641 12391 4675
rect 16497 4641 16531 4675
rect 21281 4641 21315 4675
rect 23121 4641 23155 4675
rect 25145 4641 25179 4675
rect 25697 4641 25731 4675
rect 27077 4641 27111 4675
rect 33517 4641 33551 4675
rect 2881 4573 2915 4607
rect 2973 4573 3007 4607
rect 4077 4573 4111 4607
rect 7849 4573 7883 4607
rect 10149 4573 10183 4607
rect 16405 4573 16439 4607
rect 19809 4573 19843 4607
rect 19901 4573 19935 4607
rect 21557 4573 21591 4607
rect 23857 4573 23891 4607
rect 27261 4573 27295 4607
rect 30297 4573 30331 4607
rect 2421 4505 2455 4539
rect 15945 4505 15979 4539
rect 19349 4505 19383 4539
rect 23305 4505 23339 4539
rect 24593 4505 24627 4539
rect 29837 4505 29871 4539
rect 32965 4505 32999 4539
rect 5457 4437 5491 4471
rect 6653 4437 6687 4471
rect 7021 4437 7055 4471
rect 7297 4437 7331 4471
rect 8953 4437 8987 4471
rect 10517 4437 10551 4471
rect 20269 4437 20303 4471
rect 21005 4437 21039 4471
rect 21925 4437 21959 4471
rect 24317 4437 24351 4471
rect 24869 4437 24903 4471
rect 29193 4437 29227 4471
rect 31125 4437 31159 4471
rect 4077 4233 4111 4267
rect 6653 4233 6687 4267
rect 7205 4233 7239 4267
rect 7389 4233 7423 4267
rect 15853 4233 15887 4267
rect 16313 4233 16347 4267
rect 19717 4233 19751 4267
rect 23765 4233 23799 4267
rect 25605 4233 25639 4267
rect 26801 4233 26835 4267
rect 27353 4233 27387 4267
rect 29929 4233 29963 4267
rect 33333 4233 33367 4267
rect 33609 4233 33643 4267
rect 2513 4165 2547 4199
rect 8953 4165 8987 4199
rect 19349 4165 19383 4199
rect 22845 4165 22879 4199
rect 23213 4165 23247 4199
rect 24869 4165 24903 4199
rect 26985 4165 27019 4199
rect 27077 4165 27111 4199
rect 2881 4097 2915 4131
rect 3065 4097 3099 4131
rect 3525 4097 3559 4131
rect 4537 4097 4571 4131
rect 6009 4097 6043 4131
rect 7941 4097 7975 4131
rect 16589 4097 16623 4131
rect 20085 4097 20119 4131
rect 25145 4097 25179 4131
rect 26433 4097 26467 4131
rect 1961 4029 1995 4063
rect 5641 4029 5675 4063
rect 7665 4029 7699 4063
rect 8309 4029 8343 4063
rect 9505 4029 9539 4063
rect 20821 4029 20855 4063
rect 21088 4029 21122 4063
rect 24041 4029 24075 4063
rect 2329 3961 2363 3995
rect 3893 3961 3927 3995
rect 4537 3961 4571 3995
rect 4629 3961 4663 3995
rect 7849 3961 7883 3995
rect 9229 3961 9263 3995
rect 9413 3961 9447 3995
rect 20729 3961 20763 3995
rect 24225 3961 24259 3995
rect 24317 3961 24351 3995
rect 27905 4097 27939 4131
rect 29101 4097 29135 4131
rect 30849 4097 30883 4131
rect 32965 4097 32999 4131
rect 30481 4029 30515 4063
rect 27629 3961 27663 3995
rect 30205 3961 30239 3995
rect 2973 3893 3007 3927
rect 4997 3893 5031 3927
rect 8677 3893 8711 3927
rect 22201 3893 22235 3927
rect 26985 3893 27019 3927
rect 27813 3893 27847 3927
rect 29653 3893 29687 3927
rect 30389 3893 30423 3927
rect 3249 3689 3283 3723
rect 3617 3689 3651 3723
rect 7205 3689 7239 3723
rect 7941 3689 7975 3723
rect 9321 3689 9355 3723
rect 20361 3689 20395 3723
rect 20729 3689 20763 3723
rect 21097 3689 21131 3723
rect 23765 3689 23799 3723
rect 24685 3689 24719 3723
rect 25145 3689 25179 3723
rect 27629 3689 27663 3723
rect 29837 3689 29871 3723
rect 30573 3689 30607 3723
rect 2421 3621 2455 3655
rect 7665 3621 7699 3655
rect 8953 3621 8987 3655
rect 24777 3621 24811 3655
rect 30297 3621 30331 3655
rect 1777 3553 1811 3587
rect 21557 3553 21591 3587
rect 21916 3553 21950 3587
rect 2329 3485 2363 3519
rect 2513 3485 2547 3519
rect 21649 3485 21683 3519
rect 24685 3485 24719 3519
rect 1961 3417 1995 3451
rect 24225 3417 24259 3451
rect 2973 3349 3007 3383
rect 4261 3349 4295 3383
rect 4721 3349 4755 3383
rect 23029 3349 23063 3383
rect 27353 3349 27387 3383
rect 2421 3145 2455 3179
rect 2973 3145 3007 3179
rect 21649 3145 21683 3179
rect 22017 3145 22051 3179
rect 24593 3145 24627 3179
rect 24869 3145 24903 3179
rect 20545 3077 20579 3111
rect 1961 3009 1995 3043
rect 3433 3009 3467 3043
rect 5273 3009 5307 3043
rect 20361 3009 20395 3043
rect 21097 3009 21131 3043
rect 24225 3009 24259 3043
rect 4445 2941 4479 2975
rect 19993 2941 20027 2975
rect 20821 2941 20855 2975
rect 3525 2873 3559 2907
rect 4721 2873 4755 2907
rect 21005 2873 21039 2907
rect 2697 2805 2731 2839
rect 3433 2805 3467 2839
rect 1961 2601 1995 2635
rect 2329 2601 2363 2635
rect 2973 2601 3007 2635
rect 5457 2601 5491 2635
rect 20545 2601 20579 2635
rect 3893 2465 3927 2499
rect 4344 2465 4378 2499
rect 3525 2397 3559 2431
rect 4077 2397 4111 2431
<< metal1 >>
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 7190 14056 7196 14068
rect 3476 14028 7196 14056
rect 3476 14016 3482 14028
rect 7190 14016 7196 14028
rect 7248 14016 7254 14068
rect 4062 13948 4068 14000
rect 4120 13988 4126 14000
rect 6454 13988 6460 14000
rect 4120 13960 6460 13988
rect 4120 13948 4126 13960
rect 6454 13948 6460 13960
rect 6512 13948 6518 14000
rect 3326 13880 3332 13932
rect 3384 13920 3390 13932
rect 7006 13920 7012 13932
rect 3384 13892 7012 13920
rect 3384 13880 3390 13892
rect 7006 13880 7012 13892
rect 7064 13880 7070 13932
rect 32858 13880 32864 13932
rect 32916 13920 32922 13932
rect 34790 13920 34796 13932
rect 32916 13892 34796 13920
rect 32916 13880 32922 13892
rect 34790 13880 34796 13892
rect 34848 13880 34854 13932
rect 3050 13812 3056 13864
rect 3108 13852 3114 13864
rect 7098 13852 7104 13864
rect 3108 13824 7104 13852
rect 3108 13812 3114 13824
rect 7098 13812 7104 13824
rect 7156 13812 7162 13864
rect 25406 13812 25412 13864
rect 25464 13852 25470 13864
rect 25464 13824 26648 13852
rect 25464 13812 25470 13824
rect 26620 13784 26648 13824
rect 31754 13812 31760 13864
rect 31812 13852 31818 13864
rect 34606 13852 34612 13864
rect 31812 13824 34612 13852
rect 31812 13812 31818 13824
rect 34606 13812 34612 13824
rect 34664 13812 34670 13864
rect 35158 13784 35164 13796
rect 26620 13756 35164 13784
rect 35158 13744 35164 13756
rect 35216 13744 35222 13796
rect 23566 13676 23572 13728
rect 23624 13716 23630 13728
rect 30926 13716 30932 13728
rect 23624 13688 30932 13716
rect 23624 13676 23630 13688
rect 30926 13676 30932 13688
rect 30984 13676 30990 13728
rect 31202 13676 31208 13728
rect 31260 13716 31266 13728
rect 31662 13716 31668 13728
rect 31260 13688 31668 13716
rect 31260 13676 31266 13688
rect 31662 13676 31668 13688
rect 31720 13676 31726 13728
rect 1104 13626 38824 13648
rect 1104 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 27648 13626
rect 27700 13574 27712 13626
rect 27764 13574 27776 13626
rect 27828 13574 27840 13626
rect 27892 13574 38824 13626
rect 1104 13552 38824 13574
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 4249 13515 4307 13521
rect 4249 13512 4261 13515
rect 2832 13484 4261 13512
rect 2832 13472 2838 13484
rect 4249 13481 4261 13484
rect 4295 13481 4307 13515
rect 4249 13475 4307 13481
rect 4338 13472 4344 13524
rect 4396 13512 4402 13524
rect 5353 13515 5411 13521
rect 5353 13512 5365 13515
rect 4396 13484 5365 13512
rect 4396 13472 4402 13484
rect 5353 13481 5365 13484
rect 5399 13481 5411 13515
rect 24026 13512 24032 13524
rect 5353 13475 5411 13481
rect 5460 13484 24032 13512
rect 1673 13447 1731 13453
rect 1673 13413 1685 13447
rect 1719 13444 1731 13447
rect 2130 13444 2136 13456
rect 1719 13416 2136 13444
rect 1719 13413 1731 13416
rect 1673 13407 1731 13413
rect 2130 13404 2136 13416
rect 2188 13444 2194 13456
rect 2317 13447 2375 13453
rect 2317 13444 2329 13447
rect 2188 13416 2329 13444
rect 2188 13404 2194 13416
rect 2317 13413 2329 13416
rect 2363 13413 2375 13447
rect 4614 13444 4620 13456
rect 2317 13407 2375 13413
rect 4080 13416 4620 13444
rect 4080 13385 4108 13416
rect 4614 13404 4620 13416
rect 4672 13444 4678 13456
rect 5460 13444 5488 13484
rect 24026 13472 24032 13484
rect 24084 13472 24090 13524
rect 26142 13512 26148 13524
rect 24136 13484 26148 13512
rect 4672 13416 5488 13444
rect 21637 13447 21695 13453
rect 4672 13404 4678 13416
rect 21637 13413 21649 13447
rect 21683 13444 21695 13447
rect 24136 13444 24164 13484
rect 26142 13472 26148 13484
rect 26200 13472 26206 13524
rect 28534 13512 28540 13524
rect 26528 13484 28540 13512
rect 21683 13416 24164 13444
rect 21683 13413 21695 13416
rect 21637 13407 21695 13413
rect 25498 13404 25504 13456
rect 25556 13444 25562 13456
rect 25685 13447 25743 13453
rect 25685 13444 25697 13447
rect 25556 13416 25697 13444
rect 25556 13404 25562 13416
rect 25685 13413 25697 13416
rect 25731 13444 25743 13447
rect 26528 13444 26556 13484
rect 28534 13472 28540 13484
rect 28592 13472 28598 13524
rect 31573 13515 31631 13521
rect 31573 13481 31585 13515
rect 31619 13512 31631 13515
rect 31754 13512 31760 13524
rect 31619 13484 31760 13512
rect 31619 13481 31631 13484
rect 31573 13475 31631 13481
rect 31754 13472 31760 13484
rect 31812 13472 31818 13524
rect 34425 13515 34483 13521
rect 34425 13481 34437 13515
rect 34471 13512 34483 13515
rect 34514 13512 34520 13524
rect 34471 13484 34520 13512
rect 34471 13481 34483 13484
rect 34425 13475 34483 13481
rect 34514 13472 34520 13484
rect 34572 13472 34578 13524
rect 36722 13512 36728 13524
rect 36683 13484 36728 13512
rect 36722 13472 36728 13484
rect 36780 13472 36786 13524
rect 25731 13416 26556 13444
rect 25731 13413 25743 13416
rect 25685 13407 25743 13413
rect 26602 13404 26608 13456
rect 26660 13444 26666 13456
rect 27433 13447 27491 13453
rect 27433 13444 27445 13447
rect 26660 13416 27445 13444
rect 26660 13404 26666 13416
rect 27433 13413 27445 13416
rect 27479 13413 27491 13447
rect 27433 13407 27491 13413
rect 28902 13404 28908 13456
rect 28960 13444 28966 13456
rect 30285 13447 30343 13453
rect 30285 13444 30297 13447
rect 28960 13416 30297 13444
rect 28960 13404 28966 13416
rect 30285 13413 30297 13416
rect 30331 13444 30343 13447
rect 35066 13444 35072 13456
rect 30331 13416 35072 13444
rect 30331 13413 30343 13416
rect 30285 13407 30343 13413
rect 35066 13404 35072 13416
rect 35124 13404 35130 13456
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13345 4123 13379
rect 5166 13376 5172 13388
rect 5127 13348 5172 13376
rect 4065 13339 4123 13345
rect 5166 13336 5172 13348
rect 5224 13336 5230 13388
rect 6917 13379 6975 13385
rect 6917 13345 6929 13379
rect 6963 13376 6975 13379
rect 8018 13376 8024 13388
rect 6963 13348 8024 13376
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 8018 13336 8024 13348
rect 8076 13376 8082 13388
rect 17862 13376 17868 13388
rect 8076 13348 17868 13376
rect 8076 13336 8082 13348
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 21361 13379 21419 13385
rect 21361 13345 21373 13379
rect 21407 13376 21419 13379
rect 22462 13376 22468 13388
rect 21407 13348 22468 13376
rect 21407 13345 21419 13348
rect 21361 13339 21419 13345
rect 22462 13336 22468 13348
rect 22520 13336 22526 13388
rect 22646 13376 22652 13388
rect 22607 13348 22652 13376
rect 22646 13336 22652 13348
rect 22704 13336 22710 13388
rect 22925 13379 22983 13385
rect 22925 13345 22937 13379
rect 22971 13376 22983 13379
rect 28718 13376 28724 13388
rect 22971 13348 28724 13376
rect 22971 13345 22983 13348
rect 22925 13339 22983 13345
rect 28718 13336 28724 13348
rect 28776 13336 28782 13388
rect 30098 13336 30104 13388
rect 30156 13376 30162 13388
rect 31389 13379 31447 13385
rect 30156 13348 30201 13376
rect 30156 13336 30162 13348
rect 31389 13345 31401 13379
rect 31435 13376 31447 13379
rect 32122 13376 32128 13388
rect 31435 13348 32128 13376
rect 31435 13345 31447 13348
rect 31389 13339 31447 13345
rect 2038 13268 2044 13320
rect 2096 13308 2102 13320
rect 2225 13311 2283 13317
rect 2225 13308 2237 13311
rect 2096 13280 2237 13308
rect 2096 13268 2102 13280
rect 2225 13277 2237 13280
rect 2271 13277 2283 13311
rect 2225 13271 2283 13277
rect 2240 13240 2268 13271
rect 2314 13268 2320 13320
rect 2372 13308 2378 13320
rect 2409 13311 2467 13317
rect 2409 13308 2421 13311
rect 2372 13280 2421 13308
rect 2372 13268 2378 13280
rect 2409 13277 2421 13280
rect 2455 13277 2467 13311
rect 2409 13271 2467 13277
rect 22830 13268 22836 13320
rect 22888 13308 22894 13320
rect 25406 13308 25412 13320
rect 22888 13280 25412 13308
rect 22888 13268 22894 13280
rect 25406 13268 25412 13280
rect 25464 13268 25470 13320
rect 25682 13308 25688 13320
rect 25643 13280 25688 13308
rect 25682 13268 25688 13280
rect 25740 13268 25746 13320
rect 25777 13311 25835 13317
rect 25777 13277 25789 13311
rect 25823 13277 25835 13311
rect 25777 13271 25835 13277
rect 26513 13311 26571 13317
rect 26513 13277 26525 13311
rect 26559 13308 26571 13311
rect 27341 13311 27399 13317
rect 27341 13308 27353 13311
rect 26559 13280 27353 13308
rect 26559 13277 26571 13280
rect 26513 13271 26571 13277
rect 27341 13277 27353 13280
rect 27387 13277 27399 13311
rect 27341 13271 27399 13277
rect 2777 13243 2835 13249
rect 2777 13240 2789 13243
rect 2240 13212 2789 13240
rect 2777 13209 2789 13212
rect 2823 13209 2835 13243
rect 7098 13240 7104 13252
rect 7059 13212 7104 13240
rect 2777 13203 2835 13209
rect 7098 13200 7104 13212
rect 7156 13200 7162 13252
rect 24578 13200 24584 13252
rect 24636 13240 24642 13252
rect 25792 13240 25820 13271
rect 27430 13268 27436 13320
rect 27488 13308 27494 13320
rect 27525 13311 27583 13317
rect 27525 13308 27537 13311
rect 27488 13280 27537 13308
rect 27488 13268 27494 13280
rect 27525 13277 27537 13280
rect 27571 13277 27583 13311
rect 27525 13271 27583 13277
rect 27982 13268 27988 13320
rect 28040 13308 28046 13320
rect 30116 13308 30144 13336
rect 30374 13308 30380 13320
rect 28040 13280 30144 13308
rect 30335 13280 30380 13308
rect 28040 13268 28046 13280
rect 30374 13268 30380 13280
rect 30432 13268 30438 13320
rect 31202 13308 31208 13320
rect 31163 13280 31208 13308
rect 31202 13268 31208 13280
rect 31260 13268 31266 13320
rect 25958 13240 25964 13252
rect 24636 13212 25964 13240
rect 24636 13200 24642 13212
rect 25958 13200 25964 13212
rect 26016 13200 26022 13252
rect 26050 13200 26056 13252
rect 26108 13240 26114 13252
rect 31404 13240 31432 13339
rect 32122 13336 32128 13348
rect 32180 13336 32186 13388
rect 33137 13379 33195 13385
rect 33137 13345 33149 13379
rect 33183 13376 33195 13379
rect 33410 13376 33416 13388
rect 33183 13348 33416 13376
rect 33183 13345 33195 13348
rect 33137 13339 33195 13345
rect 33410 13336 33416 13348
rect 33468 13336 33474 13388
rect 34146 13336 34152 13388
rect 34204 13376 34210 13388
rect 34241 13379 34299 13385
rect 34241 13376 34253 13379
rect 34204 13348 34253 13376
rect 34204 13336 34210 13348
rect 34241 13345 34253 13348
rect 34287 13345 34299 13379
rect 34241 13339 34299 13345
rect 35437 13379 35495 13385
rect 35437 13345 35449 13379
rect 35483 13376 35495 13379
rect 35526 13376 35532 13388
rect 35483 13348 35532 13376
rect 35483 13345 35495 13348
rect 35437 13339 35495 13345
rect 35526 13336 35532 13348
rect 35584 13336 35590 13388
rect 36538 13376 36544 13388
rect 36499 13348 36544 13376
rect 36538 13336 36544 13348
rect 36596 13336 36602 13388
rect 26108 13212 31432 13240
rect 33321 13243 33379 13249
rect 26108 13200 26114 13212
rect 33321 13209 33333 13243
rect 33367 13240 33379 13243
rect 34698 13240 34704 13252
rect 33367 13212 34704 13240
rect 33367 13209 33379 13212
rect 33321 13203 33379 13209
rect 34698 13200 34704 13212
rect 34756 13200 34762 13252
rect 1670 13132 1676 13184
rect 1728 13172 1734 13184
rect 1857 13175 1915 13181
rect 1857 13172 1869 13175
rect 1728 13144 1869 13172
rect 1728 13132 1734 13144
rect 1857 13141 1869 13144
rect 1903 13141 1915 13175
rect 1857 13135 1915 13141
rect 13722 13132 13728 13184
rect 13780 13172 13786 13184
rect 14737 13175 14795 13181
rect 14737 13172 14749 13175
rect 13780 13144 14749 13172
rect 13780 13132 13786 13144
rect 14737 13141 14749 13144
rect 14783 13141 14795 13175
rect 14737 13135 14795 13141
rect 16485 13175 16543 13181
rect 16485 13141 16497 13175
rect 16531 13172 16543 13175
rect 16942 13172 16948 13184
rect 16531 13144 16948 13172
rect 16531 13141 16543 13144
rect 16485 13135 16543 13141
rect 16942 13132 16948 13144
rect 17000 13132 17006 13184
rect 24302 13172 24308 13184
rect 24263 13144 24308 13172
rect 24302 13132 24308 13144
rect 24360 13132 24366 13184
rect 24673 13175 24731 13181
rect 24673 13141 24685 13175
rect 24719 13172 24731 13175
rect 24854 13172 24860 13184
rect 24719 13144 24860 13172
rect 24719 13141 24731 13144
rect 24673 13135 24731 13141
rect 24854 13132 24860 13144
rect 24912 13132 24918 13184
rect 25038 13172 25044 13184
rect 24999 13144 25044 13172
rect 25038 13132 25044 13144
rect 25096 13132 25102 13184
rect 25222 13172 25228 13184
rect 25183 13144 25228 13172
rect 25222 13132 25228 13144
rect 25280 13132 25286 13184
rect 25590 13132 25596 13184
rect 25648 13172 25654 13184
rect 26237 13175 26295 13181
rect 26237 13172 26249 13175
rect 25648 13144 26249 13172
rect 25648 13132 25654 13144
rect 26237 13141 26249 13144
rect 26283 13172 26295 13175
rect 26513 13175 26571 13181
rect 26513 13172 26525 13175
rect 26283 13144 26525 13172
rect 26283 13141 26295 13144
rect 26237 13135 26295 13141
rect 26513 13141 26525 13144
rect 26559 13141 26571 13175
rect 26513 13135 26571 13141
rect 26602 13132 26608 13184
rect 26660 13172 26666 13184
rect 26970 13172 26976 13184
rect 26660 13144 26705 13172
rect 26931 13144 26976 13172
rect 26660 13132 26666 13144
rect 26970 13132 26976 13144
rect 27028 13132 27034 13184
rect 27062 13132 27068 13184
rect 27120 13172 27126 13184
rect 28902 13172 28908 13184
rect 27120 13144 28908 13172
rect 27120 13132 27126 13144
rect 28902 13132 28908 13144
rect 28960 13132 28966 13184
rect 28994 13132 29000 13184
rect 29052 13172 29058 13184
rect 29457 13175 29515 13181
rect 29457 13172 29469 13175
rect 29052 13144 29469 13172
rect 29052 13132 29058 13144
rect 29457 13141 29469 13144
rect 29503 13141 29515 13175
rect 29822 13172 29828 13184
rect 29783 13144 29828 13172
rect 29457 13135 29515 13141
rect 29822 13132 29828 13144
rect 29880 13132 29886 13184
rect 35618 13172 35624 13184
rect 35579 13144 35624 13172
rect 35618 13132 35624 13144
rect 35676 13132 35682 13184
rect 1104 13082 38824 13104
rect 1104 13030 7648 13082
rect 7700 13030 7712 13082
rect 7764 13030 7776 13082
rect 7828 13030 7840 13082
rect 7892 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 34315 13082
rect 34367 13030 34379 13082
rect 34431 13030 34443 13082
rect 34495 13030 34507 13082
rect 34559 13030 38824 13082
rect 1104 13008 38824 13030
rect 4614 12968 4620 12980
rect 4575 12940 4620 12968
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 5166 12968 5172 12980
rect 5127 12940 5172 12968
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 7006 12968 7012 12980
rect 6967 12940 7012 12968
rect 7006 12928 7012 12940
rect 7064 12928 7070 12980
rect 7469 12971 7527 12977
rect 7469 12937 7481 12971
rect 7515 12968 7527 12971
rect 22830 12968 22836 12980
rect 7515 12940 22836 12968
rect 7515 12937 7527 12940
rect 7469 12931 7527 12937
rect 2317 12903 2375 12909
rect 2317 12869 2329 12903
rect 2363 12900 2375 12903
rect 2406 12900 2412 12912
rect 2363 12872 2412 12900
rect 2363 12869 2375 12872
rect 2317 12863 2375 12869
rect 2406 12860 2412 12872
rect 2464 12860 2470 12912
rect 1210 12792 1216 12844
rect 1268 12832 1274 12844
rect 3973 12835 4031 12841
rect 3973 12832 3985 12835
rect 1268 12804 3985 12832
rect 1268 12792 1274 12804
rect 3973 12801 3985 12804
rect 4019 12801 4031 12835
rect 3973 12795 4031 12801
rect 4062 12792 4068 12844
rect 4120 12832 4126 12844
rect 5626 12832 5632 12844
rect 4120 12804 5632 12832
rect 4120 12792 4126 12804
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 5721 12835 5779 12841
rect 5721 12801 5733 12835
rect 5767 12832 5779 12835
rect 6178 12832 6184 12844
rect 5767 12804 6184 12832
rect 5767 12801 5779 12804
rect 5721 12795 5779 12801
rect 6178 12792 6184 12804
rect 6236 12792 6242 12844
rect 1486 12724 1492 12776
rect 1544 12764 1550 12776
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 1544 12736 3617 12764
rect 1544 12724 1550 12736
rect 3605 12733 3617 12736
rect 3651 12764 3663 12767
rect 3789 12767 3847 12773
rect 3789 12764 3801 12767
rect 3651 12736 3801 12764
rect 3651 12733 3663 12736
rect 3605 12727 3663 12733
rect 3789 12733 3801 12736
rect 3835 12733 3847 12767
rect 3789 12727 3847 12733
rect 5350 12724 5356 12776
rect 5408 12764 5414 12776
rect 5445 12767 5503 12773
rect 5445 12764 5457 12767
rect 5408 12736 5457 12764
rect 5408 12724 5414 12736
rect 5445 12733 5457 12736
rect 5491 12764 5503 12767
rect 6273 12767 6331 12773
rect 6273 12764 6285 12767
rect 5491 12736 6285 12764
rect 5491 12733 5503 12736
rect 5445 12727 5503 12733
rect 6273 12733 6285 12736
rect 6319 12733 6331 12767
rect 6273 12727 6331 12733
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 7484 12764 7512 12931
rect 22830 12928 22836 12940
rect 22888 12928 22894 12980
rect 25498 12928 25504 12980
rect 25556 12968 25562 12980
rect 29362 12968 29368 12980
rect 25556 12940 25601 12968
rect 27724 12940 29368 12968
rect 25556 12928 25562 12940
rect 7837 12903 7895 12909
rect 7837 12869 7849 12903
rect 7883 12900 7895 12903
rect 8018 12900 8024 12912
rect 7883 12872 8024 12900
rect 7883 12869 7895 12872
rect 7837 12863 7895 12869
rect 8018 12860 8024 12872
rect 8076 12860 8082 12912
rect 14826 12900 14832 12912
rect 14787 12872 14832 12900
rect 14826 12860 14832 12872
rect 14884 12860 14890 12912
rect 14918 12860 14924 12912
rect 14976 12900 14982 12912
rect 15841 12903 15899 12909
rect 15841 12900 15853 12903
rect 14976 12872 15853 12900
rect 14976 12860 14982 12872
rect 15841 12869 15853 12872
rect 15887 12900 15899 12903
rect 16025 12903 16083 12909
rect 16025 12900 16037 12903
rect 15887 12872 16037 12900
rect 15887 12869 15899 12872
rect 15841 12863 15899 12869
rect 16025 12869 16037 12872
rect 16071 12869 16083 12903
rect 16025 12863 16083 12869
rect 16485 12903 16543 12909
rect 16485 12869 16497 12903
rect 16531 12900 16543 12903
rect 17034 12900 17040 12912
rect 16531 12872 17040 12900
rect 16531 12869 16543 12872
rect 16485 12863 16543 12869
rect 17034 12860 17040 12872
rect 17092 12860 17098 12912
rect 21542 12900 21548 12912
rect 21503 12872 21548 12900
rect 21542 12860 21548 12872
rect 21600 12860 21606 12912
rect 24026 12900 24032 12912
rect 23987 12872 24032 12900
rect 24026 12860 24032 12872
rect 24084 12860 24090 12912
rect 24578 12900 24584 12912
rect 24539 12872 24584 12900
rect 24578 12860 24584 12872
rect 24636 12860 24642 12912
rect 26234 12860 26240 12912
rect 26292 12900 26298 12912
rect 27617 12903 27675 12909
rect 27617 12900 27629 12903
rect 26292 12872 27629 12900
rect 26292 12860 26298 12872
rect 27617 12869 27629 12872
rect 27663 12869 27675 12903
rect 27617 12863 27675 12869
rect 10321 12835 10379 12841
rect 10321 12801 10333 12835
rect 10367 12832 10379 12835
rect 11146 12832 11152 12844
rect 10367 12804 11152 12832
rect 10367 12801 10379 12804
rect 10321 12795 10379 12801
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 13633 12835 13691 12841
rect 13633 12801 13645 12835
rect 13679 12832 13691 12835
rect 16206 12832 16212 12844
rect 13679 12804 16212 12832
rect 13679 12801 13691 12804
rect 13633 12795 13691 12801
rect 16206 12792 16212 12804
rect 16264 12792 16270 12844
rect 18414 12792 18420 12844
rect 18472 12832 18478 12844
rect 23566 12832 23572 12844
rect 18472 12804 23572 12832
rect 18472 12792 18478 12804
rect 23566 12792 23572 12804
rect 23624 12792 23630 12844
rect 23658 12792 23664 12844
rect 23716 12832 23722 12844
rect 24857 12835 24915 12841
rect 24857 12832 24869 12835
rect 23716 12804 24869 12832
rect 23716 12792 23722 12804
rect 24857 12801 24869 12804
rect 24903 12801 24915 12835
rect 24857 12795 24915 12801
rect 24946 12792 24952 12844
rect 25004 12832 25010 12844
rect 26421 12835 26479 12841
rect 26421 12832 26433 12835
rect 25004 12804 26433 12832
rect 25004 12792 25010 12804
rect 26421 12801 26433 12804
rect 26467 12832 26479 12835
rect 27724 12832 27752 12940
rect 29362 12928 29368 12940
rect 29420 12928 29426 12980
rect 29454 12928 29460 12980
rect 29512 12968 29518 12980
rect 34606 12968 34612 12980
rect 29512 12940 34612 12968
rect 29512 12928 29518 12940
rect 34606 12928 34612 12940
rect 34664 12928 34670 12980
rect 35621 12971 35679 12977
rect 35621 12937 35633 12971
rect 35667 12968 35679 12971
rect 35802 12968 35808 12980
rect 35667 12940 35808 12968
rect 35667 12937 35679 12940
rect 35621 12931 35679 12937
rect 35802 12928 35808 12940
rect 35860 12928 35866 12980
rect 36538 12928 36544 12980
rect 36596 12968 36602 12980
rect 37093 12971 37151 12977
rect 37093 12968 37105 12971
rect 36596 12940 37105 12968
rect 36596 12928 36602 12940
rect 37093 12937 37105 12940
rect 37139 12937 37151 12971
rect 37093 12931 37151 12937
rect 27798 12860 27804 12912
rect 27856 12900 27862 12912
rect 27856 12872 28580 12900
rect 27856 12860 27862 12872
rect 26467 12804 27752 12832
rect 28077 12835 28135 12841
rect 26467 12801 26479 12804
rect 26421 12795 26479 12801
rect 28077 12801 28089 12835
rect 28123 12832 28135 12835
rect 28442 12832 28448 12844
rect 28123 12804 28448 12832
rect 28123 12801 28135 12804
rect 28077 12795 28135 12801
rect 28442 12792 28448 12804
rect 28500 12792 28506 12844
rect 28552 12832 28580 12872
rect 28902 12860 28908 12912
rect 28960 12900 28966 12912
rect 28997 12903 29055 12909
rect 28997 12900 29009 12903
rect 28960 12872 29009 12900
rect 28960 12860 28966 12872
rect 28997 12869 29009 12872
rect 29043 12869 29055 12903
rect 28997 12863 29055 12869
rect 29641 12903 29699 12909
rect 29641 12869 29653 12903
rect 29687 12900 29699 12903
rect 29730 12900 29736 12912
rect 29687 12872 29736 12900
rect 29687 12869 29699 12872
rect 29641 12863 29699 12869
rect 29730 12860 29736 12872
rect 29788 12860 29794 12912
rect 31205 12903 31263 12909
rect 31205 12900 31217 12903
rect 29840 12872 31217 12900
rect 29840 12832 29868 12872
rect 31205 12869 31217 12872
rect 31251 12869 31263 12903
rect 31205 12863 31263 12869
rect 31386 12860 31392 12912
rect 31444 12900 31450 12912
rect 34790 12900 34796 12912
rect 31444 12872 34796 12900
rect 31444 12860 31450 12872
rect 34790 12860 34796 12872
rect 34848 12860 34854 12912
rect 30190 12832 30196 12844
rect 28552 12804 29868 12832
rect 30103 12804 30196 12832
rect 30190 12792 30196 12804
rect 30248 12832 30254 12844
rect 30374 12832 30380 12844
rect 30248 12804 30380 12832
rect 30248 12792 30254 12804
rect 30374 12792 30380 12804
rect 30432 12792 30438 12844
rect 30650 12832 30656 12844
rect 30611 12804 30656 12832
rect 30650 12792 30656 12804
rect 30708 12792 30714 12844
rect 30926 12832 30932 12844
rect 30887 12804 30932 12832
rect 30926 12792 30932 12804
rect 30984 12792 30990 12844
rect 31662 12792 31668 12844
rect 31720 12832 31726 12844
rect 32861 12835 32919 12841
rect 32861 12832 32873 12835
rect 31720 12804 32873 12832
rect 31720 12792 31726 12804
rect 32861 12801 32873 12804
rect 32907 12801 32919 12835
rect 32861 12795 32919 12801
rect 33594 12792 33600 12844
rect 33652 12832 33658 12844
rect 35526 12832 35532 12844
rect 33652 12804 35532 12832
rect 33652 12792 33658 12804
rect 35526 12792 35532 12804
rect 35584 12832 35590 12844
rect 35989 12835 36047 12841
rect 35989 12832 36001 12835
rect 35584 12804 36001 12832
rect 35584 12792 35590 12804
rect 35989 12801 36001 12804
rect 36035 12801 36047 12835
rect 35989 12795 36047 12801
rect 6871 12736 7512 12764
rect 10045 12767 10103 12773
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 10045 12733 10057 12767
rect 10091 12764 10103 12767
rect 13357 12767 13415 12773
rect 13357 12764 13369 12767
rect 10091 12736 10916 12764
rect 10091 12733 10103 12736
rect 10045 12727 10103 12733
rect 2593 12699 2651 12705
rect 2593 12696 2605 12699
rect 1688 12668 2605 12696
rect 1394 12588 1400 12640
rect 1452 12628 1458 12640
rect 1688 12637 1716 12668
rect 2593 12665 2605 12668
rect 2639 12665 2651 12699
rect 2866 12696 2872 12708
rect 2827 12668 2872 12696
rect 2593 12659 2651 12665
rect 2866 12656 2872 12668
rect 2924 12656 2930 12708
rect 6840 12696 6868 12727
rect 3160 12668 6868 12696
rect 1673 12631 1731 12637
rect 1673 12628 1685 12631
rect 1452 12600 1685 12628
rect 1452 12588 1458 12600
rect 1673 12597 1685 12600
rect 1719 12597 1731 12631
rect 1673 12591 1731 12597
rect 2133 12631 2191 12637
rect 2133 12597 2145 12631
rect 2179 12628 2191 12631
rect 2777 12631 2835 12637
rect 2777 12628 2789 12631
rect 2179 12600 2789 12628
rect 2179 12597 2191 12600
rect 2133 12591 2191 12597
rect 2777 12597 2789 12600
rect 2823 12628 2835 12631
rect 3160 12628 3188 12668
rect 10888 12640 10916 12736
rect 13188 12736 13369 12764
rect 2823 12600 3188 12628
rect 3329 12631 3387 12637
rect 2823 12597 2835 12600
rect 2777 12591 2835 12597
rect 3329 12597 3341 12631
rect 3375 12628 3387 12631
rect 3510 12628 3516 12640
rect 3375 12600 3516 12628
rect 3375 12597 3387 12600
rect 3329 12591 3387 12597
rect 3510 12588 3516 12600
rect 3568 12588 3574 12640
rect 10870 12628 10876 12640
rect 10831 12600 10876 12628
rect 10870 12588 10876 12600
rect 10928 12588 10934 12640
rect 12526 12588 12532 12640
rect 12584 12628 12590 12640
rect 13188 12637 13216 12736
rect 13357 12733 13369 12736
rect 13403 12733 13415 12767
rect 13357 12727 13415 12733
rect 13722 12724 13728 12776
rect 13780 12764 13786 12776
rect 16301 12767 16359 12773
rect 13780 12736 15332 12764
rect 13780 12724 13786 12736
rect 15304 12705 15332 12736
rect 16301 12733 16313 12767
rect 16347 12764 16359 12767
rect 16347 12736 16804 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 14277 12699 14335 12705
rect 14277 12665 14289 12699
rect 14323 12696 14335 12699
rect 15105 12699 15163 12705
rect 15105 12696 15117 12699
rect 14323 12668 15117 12696
rect 14323 12665 14335 12668
rect 14277 12659 14335 12665
rect 15105 12665 15117 12668
rect 15151 12665 15163 12699
rect 15105 12659 15163 12665
rect 15289 12699 15347 12705
rect 15289 12665 15301 12699
rect 15335 12665 15347 12699
rect 15289 12659 15347 12665
rect 13173 12631 13231 12637
rect 13173 12628 13185 12631
rect 12584 12600 13185 12628
rect 12584 12588 12590 12600
rect 13173 12597 13185 12600
rect 13219 12597 13231 12631
rect 13173 12591 13231 12597
rect 14645 12631 14703 12637
rect 14645 12597 14657 12631
rect 14691 12628 14703 12631
rect 15010 12628 15016 12640
rect 14691 12600 15016 12628
rect 14691 12597 14703 12600
rect 14645 12591 14703 12597
rect 15010 12588 15016 12600
rect 15068 12588 15074 12640
rect 15120 12628 15148 12659
rect 15378 12656 15384 12708
rect 15436 12696 15442 12708
rect 16776 12705 16804 12736
rect 16942 12724 16948 12776
rect 17000 12764 17006 12776
rect 17037 12767 17095 12773
rect 17037 12764 17049 12767
rect 17000 12736 17049 12764
rect 17000 12724 17006 12736
rect 17037 12733 17049 12736
rect 17083 12733 17095 12767
rect 22370 12764 22376 12776
rect 17037 12727 17095 12733
rect 21836 12736 22376 12764
rect 16761 12699 16819 12705
rect 15436 12668 15481 12696
rect 15436 12656 15442 12668
rect 16761 12665 16773 12699
rect 16807 12696 16819 12699
rect 20438 12696 20444 12708
rect 16807 12668 20444 12696
rect 16807 12665 16819 12668
rect 16761 12659 16819 12665
rect 20438 12656 20444 12668
rect 20496 12656 20502 12708
rect 21836 12705 21864 12736
rect 22370 12724 22376 12736
rect 22428 12724 22434 12776
rect 22646 12724 22652 12776
rect 22704 12764 22710 12776
rect 22925 12767 22983 12773
rect 22925 12764 22937 12767
rect 22704 12736 22937 12764
rect 22704 12724 22710 12736
rect 22925 12733 22937 12736
rect 22971 12764 22983 12767
rect 22971 12736 24072 12764
rect 22971 12733 22983 12736
rect 22925 12727 22983 12733
rect 20993 12699 21051 12705
rect 20993 12665 21005 12699
rect 21039 12696 21051 12699
rect 21821 12699 21879 12705
rect 21821 12696 21833 12699
rect 21039 12668 21833 12696
rect 21039 12665 21051 12668
rect 20993 12659 21051 12665
rect 21821 12665 21833 12668
rect 21867 12665 21879 12699
rect 21821 12659 21879 12665
rect 22097 12699 22155 12705
rect 22097 12665 22109 12699
rect 22143 12696 22155 12699
rect 22186 12696 22192 12708
rect 22143 12668 22192 12696
rect 22143 12665 22155 12668
rect 22097 12659 22155 12665
rect 22186 12656 22192 12668
rect 22244 12656 22250 12708
rect 15746 12628 15752 12640
rect 15120 12600 15752 12628
rect 15746 12588 15752 12600
rect 15804 12588 15810 12640
rect 16025 12631 16083 12637
rect 16025 12597 16037 12631
rect 16071 12628 16083 12631
rect 16945 12631 17003 12637
rect 16945 12628 16957 12631
rect 16071 12600 16957 12628
rect 16071 12597 16083 12600
rect 16025 12591 16083 12597
rect 16945 12597 16957 12600
rect 16991 12597 17003 12631
rect 20530 12628 20536 12640
rect 20491 12600 20536 12628
rect 16945 12591 17003 12597
rect 20530 12588 20536 12600
rect 20588 12588 20594 12640
rect 20806 12588 20812 12640
rect 20864 12628 20870 12640
rect 21269 12631 21327 12637
rect 21269 12628 21281 12631
rect 20864 12600 21281 12628
rect 20864 12588 20870 12600
rect 21269 12597 21281 12600
rect 21315 12628 21327 12631
rect 22005 12631 22063 12637
rect 22005 12628 22017 12631
rect 21315 12600 22017 12628
rect 21315 12597 21327 12600
rect 21269 12591 21327 12597
rect 22005 12597 22017 12600
rect 22051 12597 22063 12631
rect 22005 12591 22063 12597
rect 22462 12588 22468 12640
rect 22520 12628 22526 12640
rect 22557 12631 22615 12637
rect 22557 12628 22569 12631
rect 22520 12600 22569 12628
rect 22520 12588 22526 12600
rect 22557 12597 22569 12600
rect 22603 12628 22615 12631
rect 23014 12628 23020 12640
rect 22603 12600 23020 12628
rect 22603 12597 22615 12600
rect 22557 12591 22615 12597
rect 23014 12588 23020 12600
rect 23072 12588 23078 12640
rect 24044 12628 24072 12736
rect 24302 12724 24308 12776
rect 24360 12764 24366 12776
rect 24673 12767 24731 12773
rect 24673 12764 24685 12767
rect 24360 12736 24685 12764
rect 24360 12724 24366 12736
rect 24673 12733 24685 12736
rect 24719 12764 24731 12767
rect 26035 12767 26093 12773
rect 26035 12764 26047 12767
rect 24719 12736 26047 12764
rect 24719 12733 24731 12736
rect 24673 12727 24731 12733
rect 26035 12733 26047 12736
rect 26081 12733 26093 12767
rect 26035 12727 26093 12733
rect 26694 12724 26700 12776
rect 26752 12764 26758 12776
rect 28629 12767 28687 12773
rect 28629 12764 28641 12767
rect 26752 12736 28641 12764
rect 26752 12724 26758 12736
rect 28629 12733 28641 12736
rect 28675 12764 28687 12767
rect 28675 12736 30144 12764
rect 28675 12733 28687 12736
rect 28629 12727 28687 12733
rect 25038 12656 25044 12708
rect 25096 12696 25102 12708
rect 25096 12668 26188 12696
rect 25096 12656 25102 12668
rect 25774 12628 25780 12640
rect 24044 12600 25780 12628
rect 25774 12588 25780 12600
rect 25832 12588 25838 12640
rect 25866 12588 25872 12640
rect 25924 12628 25930 12640
rect 26160 12628 26188 12668
rect 26418 12656 26424 12708
rect 26476 12696 26482 12708
rect 26605 12699 26663 12705
rect 26605 12696 26617 12699
rect 26476 12668 26617 12696
rect 26476 12656 26482 12668
rect 26605 12665 26617 12668
rect 26651 12665 26663 12699
rect 26605 12659 26663 12665
rect 27065 12699 27123 12705
rect 27065 12665 27077 12699
rect 27111 12696 27123 12699
rect 28169 12699 28227 12705
rect 28169 12696 28181 12699
rect 27111 12668 28181 12696
rect 27111 12665 27123 12668
rect 27065 12659 27123 12665
rect 28169 12665 28181 12668
rect 28215 12696 28227 12699
rect 28350 12696 28356 12708
rect 28215 12668 28356 12696
rect 28215 12665 28227 12668
rect 28169 12659 28227 12665
rect 28350 12656 28356 12668
rect 28408 12656 28414 12708
rect 29086 12656 29092 12708
rect 29144 12696 29150 12708
rect 29914 12696 29920 12708
rect 29144 12668 29920 12696
rect 29144 12656 29150 12668
rect 29914 12656 29920 12668
rect 29972 12656 29978 12708
rect 30116 12705 30144 12736
rect 30101 12699 30159 12705
rect 30101 12665 30113 12699
rect 30147 12665 30159 12699
rect 30944 12696 30972 12792
rect 31202 12724 31208 12776
rect 31260 12764 31266 12776
rect 31481 12767 31539 12773
rect 31481 12764 31493 12767
rect 31260 12736 31493 12764
rect 31260 12724 31266 12736
rect 31481 12733 31493 12736
rect 31527 12733 31539 12767
rect 32122 12764 32128 12776
rect 31481 12727 31539 12733
rect 31680 12736 31984 12764
rect 32083 12736 32128 12764
rect 31680 12705 31708 12736
rect 31665 12699 31723 12705
rect 31665 12696 31677 12699
rect 30944 12668 31677 12696
rect 30101 12659 30159 12665
rect 31665 12665 31677 12668
rect 31711 12665 31723 12699
rect 31665 12659 31723 12665
rect 31754 12656 31760 12708
rect 31812 12696 31818 12708
rect 31956 12696 31984 12736
rect 32122 12724 32128 12736
rect 32180 12724 32186 12776
rect 32401 12767 32459 12773
rect 32401 12733 32413 12767
rect 32447 12764 32459 12767
rect 32677 12767 32735 12773
rect 32677 12764 32689 12767
rect 32447 12736 32689 12764
rect 32447 12733 32459 12736
rect 32401 12727 32459 12733
rect 32677 12733 32689 12736
rect 32723 12733 32735 12767
rect 35434 12764 35440 12776
rect 35395 12736 35440 12764
rect 32677 12727 32735 12733
rect 35434 12724 35440 12736
rect 35492 12724 35498 12776
rect 36541 12767 36599 12773
rect 36541 12733 36553 12767
rect 36587 12733 36599 12767
rect 36541 12727 36599 12733
rect 36357 12699 36415 12705
rect 36357 12696 36369 12699
rect 31812 12668 31857 12696
rect 31956 12668 36369 12696
rect 31812 12656 31818 12668
rect 36357 12665 36369 12668
rect 36403 12696 36415 12699
rect 36556 12696 36584 12727
rect 36403 12668 36584 12696
rect 36403 12665 36415 12668
rect 36357 12659 36415 12665
rect 26513 12631 26571 12637
rect 26513 12628 26525 12631
rect 25924 12600 25969 12628
rect 26160 12600 26525 12628
rect 25924 12588 25930 12600
rect 26513 12597 26525 12600
rect 26559 12628 26571 12631
rect 26970 12628 26976 12640
rect 26559 12600 26976 12628
rect 26559 12597 26571 12600
rect 26513 12591 26571 12597
rect 26970 12588 26976 12600
rect 27028 12588 27034 12640
rect 27433 12631 27491 12637
rect 27433 12597 27445 12631
rect 27479 12628 27491 12631
rect 28077 12631 28135 12637
rect 28077 12628 28089 12631
rect 27479 12600 28089 12628
rect 27479 12597 27491 12600
rect 27433 12591 27491 12597
rect 28077 12597 28089 12600
rect 28123 12628 28135 12631
rect 28258 12628 28264 12640
rect 28123 12600 28264 12628
rect 28123 12597 28135 12600
rect 28077 12591 28135 12597
rect 28258 12588 28264 12600
rect 28316 12588 28322 12640
rect 29638 12588 29644 12640
rect 29696 12628 29702 12640
rect 32401 12631 32459 12637
rect 32401 12628 32413 12631
rect 29696 12600 32413 12628
rect 29696 12588 29702 12600
rect 32401 12597 32413 12600
rect 32447 12628 32459 12631
rect 32493 12631 32551 12637
rect 32493 12628 32505 12631
rect 32447 12600 32505 12628
rect 32447 12597 32459 12600
rect 32401 12591 32459 12597
rect 32493 12597 32505 12600
rect 32539 12597 32551 12631
rect 33410 12628 33416 12640
rect 33371 12600 33416 12628
rect 32493 12591 32551 12597
rect 33410 12588 33416 12600
rect 33468 12588 33474 12640
rect 34238 12628 34244 12640
rect 34199 12600 34244 12628
rect 34238 12588 34244 12600
rect 34296 12588 34302 12640
rect 34790 12588 34796 12640
rect 34848 12628 34854 12640
rect 35253 12631 35311 12637
rect 35253 12628 35265 12631
rect 34848 12600 35265 12628
rect 34848 12588 34854 12600
rect 35253 12597 35265 12600
rect 35299 12628 35311 12631
rect 35434 12628 35440 12640
rect 35299 12600 35440 12628
rect 35299 12597 35311 12600
rect 35253 12591 35311 12597
rect 35434 12588 35440 12600
rect 35492 12588 35498 12640
rect 36722 12628 36728 12640
rect 36683 12600 36728 12628
rect 36722 12588 36728 12600
rect 36780 12588 36786 12640
rect 1104 12538 38824 12560
rect 1104 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 27648 12538
rect 27700 12486 27712 12538
rect 27764 12486 27776 12538
rect 27828 12486 27840 12538
rect 27892 12486 38824 12538
rect 1104 12464 38824 12486
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 5353 12427 5411 12433
rect 5353 12424 5365 12427
rect 4212 12396 5365 12424
rect 4212 12384 4218 12396
rect 5353 12393 5365 12396
rect 5399 12393 5411 12427
rect 6454 12424 6460 12436
rect 6415 12396 6460 12424
rect 5353 12387 5411 12393
rect 6454 12384 6460 12396
rect 6512 12384 6518 12436
rect 7190 12384 7196 12436
rect 7248 12424 7254 12436
rect 7561 12427 7619 12433
rect 7561 12424 7573 12427
rect 7248 12396 7573 12424
rect 7248 12384 7254 12396
rect 7561 12393 7573 12396
rect 7607 12393 7619 12427
rect 7561 12387 7619 12393
rect 20530 12384 20536 12436
rect 20588 12424 20594 12436
rect 22186 12424 22192 12436
rect 20588 12396 22192 12424
rect 20588 12384 20594 12396
rect 22186 12384 22192 12396
rect 22244 12384 22250 12436
rect 25409 12427 25467 12433
rect 25409 12393 25421 12427
rect 25455 12424 25467 12427
rect 26326 12424 26332 12436
rect 25455 12396 26332 12424
rect 25455 12393 25467 12396
rect 25409 12387 25467 12393
rect 26326 12384 26332 12396
rect 26384 12424 26390 12436
rect 27522 12424 27528 12436
rect 26384 12396 27528 12424
rect 26384 12384 26390 12396
rect 27522 12384 27528 12396
rect 27580 12384 27586 12436
rect 28258 12424 28264 12436
rect 28219 12396 28264 12424
rect 28258 12384 28264 12396
rect 28316 12384 28322 12436
rect 29914 12384 29920 12436
rect 29972 12424 29978 12436
rect 30377 12427 30435 12433
rect 30377 12424 30389 12427
rect 29972 12396 30389 12424
rect 29972 12384 29978 12396
rect 30377 12393 30389 12396
rect 30423 12393 30435 12427
rect 30377 12387 30435 12393
rect 31113 12427 31171 12433
rect 31113 12393 31125 12427
rect 31159 12424 31171 12427
rect 31386 12424 31392 12436
rect 31159 12396 31392 12424
rect 31159 12393 31171 12396
rect 31113 12387 31171 12393
rect 31386 12384 31392 12396
rect 31444 12384 31450 12436
rect 31573 12427 31631 12433
rect 31573 12393 31585 12427
rect 31619 12424 31631 12427
rect 31662 12424 31668 12436
rect 31619 12396 31668 12424
rect 31619 12393 31631 12396
rect 31573 12387 31631 12393
rect 31662 12384 31668 12396
rect 31720 12384 31726 12436
rect 32858 12424 32864 12436
rect 32819 12396 32864 12424
rect 32858 12384 32864 12396
rect 32916 12384 32922 12436
rect 2498 12316 2504 12368
rect 2556 12356 2562 12368
rect 2685 12359 2743 12365
rect 2685 12356 2697 12359
rect 2556 12328 2697 12356
rect 2556 12316 2562 12328
rect 2685 12325 2697 12328
rect 2731 12325 2743 12359
rect 2685 12319 2743 12325
rect 12066 12316 12072 12368
rect 12124 12356 12130 12368
rect 12529 12359 12587 12365
rect 12529 12356 12541 12359
rect 12124 12328 12541 12356
rect 12124 12316 12130 12328
rect 12529 12325 12541 12328
rect 12575 12325 12587 12359
rect 12529 12319 12587 12325
rect 13630 12316 13636 12368
rect 13688 12356 13694 12368
rect 13817 12359 13875 12365
rect 13817 12356 13829 12359
rect 13688 12328 13829 12356
rect 13688 12316 13694 12328
rect 13817 12325 13829 12328
rect 13863 12325 13875 12359
rect 13817 12319 13875 12325
rect 16945 12359 17003 12365
rect 16945 12325 16957 12359
rect 16991 12356 17003 12359
rect 17034 12356 17040 12368
rect 16991 12328 17040 12356
rect 16991 12325 17003 12328
rect 16945 12319 17003 12325
rect 17034 12316 17040 12328
rect 17092 12316 17098 12368
rect 18233 12359 18291 12365
rect 18233 12325 18245 12359
rect 18279 12356 18291 12359
rect 18690 12356 18696 12368
rect 18279 12328 18696 12356
rect 18279 12325 18291 12328
rect 18233 12319 18291 12325
rect 18690 12316 18696 12328
rect 18748 12316 18754 12368
rect 19797 12359 19855 12365
rect 19797 12325 19809 12359
rect 19843 12356 19855 12359
rect 20622 12356 20628 12368
rect 19843 12328 20628 12356
rect 19843 12325 19855 12328
rect 19797 12319 19855 12325
rect 20622 12316 20628 12328
rect 20680 12316 20686 12368
rect 21726 12356 21732 12368
rect 21687 12328 21732 12356
rect 21726 12316 21732 12328
rect 21784 12316 21790 12368
rect 23290 12356 23296 12368
rect 23251 12328 23296 12356
rect 23290 12316 23296 12328
rect 23348 12316 23354 12368
rect 24946 12316 24952 12368
rect 25004 12356 25010 12368
rect 25225 12359 25283 12365
rect 25225 12356 25237 12359
rect 25004 12328 25237 12356
rect 25004 12316 25010 12328
rect 25225 12325 25237 12328
rect 25271 12325 25283 12359
rect 25225 12319 25283 12325
rect 25774 12316 25780 12368
rect 25832 12356 25838 12368
rect 26234 12356 26240 12368
rect 25832 12328 26240 12356
rect 25832 12316 25838 12328
rect 26234 12316 26240 12328
rect 26292 12316 26298 12368
rect 28350 12356 28356 12368
rect 28311 12328 28356 12356
rect 28350 12316 28356 12328
rect 28408 12316 28414 12368
rect 28813 12359 28871 12365
rect 28813 12325 28825 12359
rect 28859 12356 28871 12359
rect 29822 12356 29828 12368
rect 28859 12328 29828 12356
rect 28859 12325 28871 12328
rect 28813 12319 28871 12325
rect 29822 12316 29828 12328
rect 29880 12316 29886 12368
rect 34054 12356 34060 12368
rect 34015 12328 34060 12356
rect 34054 12316 34060 12328
rect 34112 12316 34118 12368
rect 3418 12248 3424 12300
rect 3476 12288 3482 12300
rect 4065 12291 4123 12297
rect 4065 12288 4077 12291
rect 3476 12260 4077 12288
rect 3476 12248 3482 12260
rect 4065 12257 4077 12260
rect 4111 12257 4123 12291
rect 5166 12288 5172 12300
rect 5127 12260 5172 12288
rect 4065 12251 4123 12257
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 6178 12248 6184 12300
rect 6236 12288 6242 12300
rect 6273 12291 6331 12297
rect 6273 12288 6285 12291
rect 6236 12260 6285 12288
rect 6236 12248 6242 12260
rect 6273 12257 6285 12260
rect 6319 12257 6331 12291
rect 7374 12288 7380 12300
rect 7335 12260 7380 12288
rect 6273 12251 6331 12257
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 12342 12288 12348 12300
rect 12303 12260 12348 12288
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 13541 12291 13599 12297
rect 13541 12257 13553 12291
rect 13587 12288 13599 12291
rect 13906 12288 13912 12300
rect 13587 12260 13912 12288
rect 13587 12257 13599 12260
rect 13541 12251 13599 12257
rect 13906 12248 13912 12260
rect 13964 12288 13970 12300
rect 14826 12288 14832 12300
rect 13964 12260 14832 12288
rect 13964 12248 13970 12260
rect 14826 12248 14832 12260
rect 14884 12248 14890 12300
rect 17954 12288 17960 12300
rect 17915 12260 17960 12288
rect 17954 12248 17960 12260
rect 18012 12288 18018 12300
rect 18785 12291 18843 12297
rect 18785 12288 18797 12291
rect 18012 12260 18797 12288
rect 18012 12248 18018 12260
rect 18785 12257 18797 12260
rect 18831 12257 18843 12291
rect 19518 12288 19524 12300
rect 19479 12260 19524 12288
rect 18785 12251 18843 12257
rect 19518 12248 19524 12260
rect 19576 12248 19582 12300
rect 21542 12288 21548 12300
rect 21503 12260 21548 12288
rect 21542 12248 21548 12260
rect 21600 12248 21606 12300
rect 22922 12248 22928 12300
rect 22980 12288 22986 12300
rect 23109 12291 23167 12297
rect 23109 12288 23121 12291
rect 22980 12260 23121 12288
rect 22980 12248 22986 12260
rect 23109 12257 23121 12260
rect 23155 12257 23167 12291
rect 25498 12288 25504 12300
rect 23109 12251 23167 12257
rect 24688 12260 25504 12288
rect 2685 12223 2743 12229
rect 2685 12189 2697 12223
rect 2731 12189 2743 12223
rect 2685 12183 2743 12189
rect 2777 12223 2835 12229
rect 2777 12189 2789 12223
rect 2823 12220 2835 12223
rect 2866 12220 2872 12232
rect 2823 12192 2872 12220
rect 2823 12189 2835 12192
rect 2777 12183 2835 12189
rect 1857 12155 1915 12161
rect 1857 12121 1869 12155
rect 1903 12152 1915 12155
rect 2314 12152 2320 12164
rect 1903 12124 2320 12152
rect 1903 12121 1915 12124
rect 1857 12115 1915 12121
rect 2314 12112 2320 12124
rect 2372 12112 2378 12164
rect 2700 12152 2728 12183
rect 2866 12180 2872 12192
rect 2924 12220 2930 12232
rect 3237 12223 3295 12229
rect 3237 12220 3249 12223
rect 2924 12192 3249 12220
rect 2924 12180 2930 12192
rect 3237 12189 3249 12192
rect 3283 12220 3295 12223
rect 3510 12220 3516 12232
rect 3283 12192 3516 12220
rect 3283 12189 3295 12192
rect 3237 12183 3295 12189
rect 3510 12180 3516 12192
rect 3568 12220 3574 12232
rect 3878 12220 3884 12232
rect 3568 12192 3884 12220
rect 3568 12180 3574 12192
rect 3878 12180 3884 12192
rect 3936 12220 3942 12232
rect 4617 12223 4675 12229
rect 4617 12220 4629 12223
rect 3936 12192 4629 12220
rect 3936 12180 3942 12192
rect 4617 12189 4629 12192
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12220 12679 12223
rect 12710 12220 12716 12232
rect 12667 12192 12716 12220
rect 12667 12189 12679 12192
rect 12621 12183 12679 12189
rect 12710 12180 12716 12192
rect 12768 12180 12774 12232
rect 16853 12223 16911 12229
rect 16853 12189 16865 12223
rect 16899 12189 16911 12223
rect 16853 12183 16911 12189
rect 17037 12223 17095 12229
rect 17037 12189 17049 12223
rect 17083 12220 17095 12223
rect 17126 12220 17132 12232
rect 17083 12192 17132 12220
rect 17083 12189 17095 12192
rect 17037 12183 17095 12189
rect 4246 12152 4252 12164
rect 2700 12124 3648 12152
rect 4207 12124 4252 12152
rect 3620 12096 3648 12124
rect 4246 12112 4252 12124
rect 4304 12112 4310 12164
rect 16114 12112 16120 12164
rect 16172 12152 16178 12164
rect 16485 12155 16543 12161
rect 16485 12152 16497 12155
rect 16172 12124 16497 12152
rect 16172 12112 16178 12124
rect 16485 12121 16497 12124
rect 16531 12121 16543 12155
rect 16485 12115 16543 12121
rect 2222 12084 2228 12096
rect 2183 12056 2228 12084
rect 2222 12044 2228 12056
rect 2280 12044 2286 12096
rect 3602 12084 3608 12096
rect 3563 12056 3608 12084
rect 3602 12044 3608 12056
rect 3660 12044 3666 12096
rect 6822 12084 6828 12096
rect 6783 12056 6828 12084
rect 6822 12044 6828 12056
rect 6880 12044 6886 12096
rect 9217 12087 9275 12093
rect 9217 12053 9229 12087
rect 9263 12084 9275 12087
rect 9490 12084 9496 12096
rect 9263 12056 9496 12084
rect 9263 12053 9275 12056
rect 9217 12047 9275 12053
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 12069 12087 12127 12093
rect 12069 12053 12081 12087
rect 12115 12084 12127 12087
rect 12986 12084 12992 12096
rect 12115 12056 12992 12084
rect 12115 12053 12127 12056
rect 12069 12047 12127 12053
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 14921 12087 14979 12093
rect 14921 12053 14933 12087
rect 14967 12084 14979 12087
rect 15102 12084 15108 12096
rect 14967 12056 15108 12084
rect 14967 12053 14979 12056
rect 14921 12047 14979 12053
rect 15102 12044 15108 12056
rect 15160 12044 15166 12096
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 16209 12087 16267 12093
rect 16209 12084 16221 12087
rect 16080 12056 16221 12084
rect 16080 12044 16086 12056
rect 16209 12053 16221 12056
rect 16255 12084 16267 12087
rect 16868 12084 16896 12183
rect 17126 12180 17132 12192
rect 17184 12180 17190 12232
rect 21818 12220 21824 12232
rect 21779 12192 21824 12220
rect 21818 12180 21824 12192
rect 21876 12180 21882 12232
rect 23385 12223 23443 12229
rect 23385 12189 23397 12223
rect 23431 12220 23443 12223
rect 23842 12220 23848 12232
rect 23431 12192 23848 12220
rect 23431 12189 23443 12192
rect 23385 12183 23443 12189
rect 23842 12180 23848 12192
rect 23900 12180 23906 12232
rect 24029 12155 24087 12161
rect 24029 12121 24041 12155
rect 24075 12152 24087 12155
rect 24578 12152 24584 12164
rect 24075 12124 24584 12152
rect 24075 12121 24087 12124
rect 24029 12115 24087 12121
rect 24578 12112 24584 12124
rect 24636 12152 24642 12164
rect 24688 12161 24716 12260
rect 25498 12248 25504 12260
rect 25556 12248 25562 12300
rect 30190 12288 30196 12300
rect 29104 12260 30196 12288
rect 26970 12220 26976 12232
rect 26883 12192 26976 12220
rect 26970 12180 26976 12192
rect 27028 12220 27034 12232
rect 27430 12220 27436 12232
rect 27028 12192 27436 12220
rect 27028 12180 27034 12192
rect 27430 12180 27436 12192
rect 27488 12180 27494 12232
rect 28261 12223 28319 12229
rect 28261 12189 28273 12223
rect 28307 12220 28319 12223
rect 28810 12220 28816 12232
rect 28307 12192 28816 12220
rect 28307 12189 28319 12192
rect 28261 12183 28319 12189
rect 28810 12180 28816 12192
rect 28868 12180 28874 12232
rect 28994 12180 29000 12232
rect 29052 12220 29058 12232
rect 29104 12229 29132 12260
rect 30190 12248 30196 12260
rect 30248 12288 30254 12300
rect 30650 12288 30656 12300
rect 30248 12260 30656 12288
rect 30248 12248 30254 12260
rect 30650 12248 30656 12260
rect 30708 12248 30714 12300
rect 30929 12291 30987 12297
rect 30929 12257 30941 12291
rect 30975 12257 30987 12291
rect 32674 12288 32680 12300
rect 32635 12260 32680 12288
rect 30929 12251 30987 12257
rect 29089 12223 29147 12229
rect 29089 12220 29101 12223
rect 29052 12192 29101 12220
rect 29052 12180 29058 12192
rect 29089 12189 29101 12192
rect 29135 12189 29147 12223
rect 29822 12220 29828 12232
rect 29783 12192 29828 12220
rect 29089 12183 29147 12189
rect 29822 12180 29828 12192
rect 29880 12180 29886 12232
rect 29914 12180 29920 12232
rect 29972 12220 29978 12232
rect 29972 12192 30017 12220
rect 29972 12180 29978 12192
rect 30558 12180 30564 12232
rect 30616 12220 30622 12232
rect 30944 12220 30972 12251
rect 32674 12248 32680 12260
rect 32732 12248 32738 12300
rect 33778 12288 33784 12300
rect 33739 12260 33784 12288
rect 33778 12248 33784 12260
rect 33836 12248 33842 12300
rect 34974 12248 34980 12300
rect 35032 12288 35038 12300
rect 35437 12291 35495 12297
rect 35437 12288 35449 12291
rect 35032 12260 35449 12288
rect 35032 12248 35038 12260
rect 35437 12257 35449 12260
rect 35483 12257 35495 12291
rect 35437 12251 35495 12257
rect 36446 12248 36452 12300
rect 36504 12288 36510 12300
rect 36541 12291 36599 12297
rect 36541 12288 36553 12291
rect 36504 12260 36553 12288
rect 36504 12248 36510 12260
rect 36541 12257 36553 12260
rect 36587 12257 36599 12291
rect 36541 12251 36599 12257
rect 30616 12192 30972 12220
rect 30616 12180 30622 12192
rect 24673 12155 24731 12161
rect 24673 12152 24685 12155
rect 24636 12124 24685 12152
rect 24636 12112 24642 12124
rect 24673 12121 24685 12124
rect 24719 12121 24731 12155
rect 24673 12115 24731 12121
rect 24949 12155 25007 12161
rect 24949 12121 24961 12155
rect 24995 12152 25007 12155
rect 25590 12152 25596 12164
rect 24995 12124 25596 12152
rect 24995 12121 25007 12124
rect 24949 12115 25007 12121
rect 25590 12112 25596 12124
rect 25648 12112 25654 12164
rect 27617 12155 27675 12161
rect 27617 12121 27629 12155
rect 27663 12152 27675 12155
rect 28442 12152 28448 12164
rect 27663 12124 28448 12152
rect 27663 12121 27675 12124
rect 27617 12115 27675 12121
rect 28442 12112 28448 12124
rect 28500 12152 28506 12164
rect 28626 12152 28632 12164
rect 28500 12124 28632 12152
rect 28500 12112 28506 12124
rect 28626 12112 28632 12124
rect 28684 12112 28690 12164
rect 29362 12152 29368 12164
rect 29323 12124 29368 12152
rect 29362 12112 29368 12124
rect 29420 12112 29426 12164
rect 16255 12056 16896 12084
rect 20717 12087 20775 12093
rect 16255 12053 16267 12056
rect 16209 12047 16267 12053
rect 20717 12053 20729 12087
rect 20763 12084 20775 12087
rect 21266 12084 21272 12096
rect 20763 12056 21272 12084
rect 20763 12053 20775 12056
rect 20717 12047 20775 12053
rect 21266 12044 21272 12056
rect 21324 12044 21330 12096
rect 21726 12044 21732 12096
rect 21784 12084 21790 12096
rect 22833 12087 22891 12093
rect 22833 12084 22845 12087
rect 21784 12056 22845 12084
rect 21784 12044 21790 12056
rect 22833 12053 22845 12056
rect 22879 12053 22891 12087
rect 24394 12084 24400 12096
rect 24355 12056 24400 12084
rect 22833 12047 22891 12053
rect 24394 12044 24400 12056
rect 24452 12044 24458 12096
rect 25682 12044 25688 12096
rect 25740 12084 25746 12096
rect 25961 12087 26019 12093
rect 25961 12084 25973 12087
rect 25740 12056 25973 12084
rect 25740 12044 25746 12056
rect 25961 12053 25973 12056
rect 26007 12084 26019 12087
rect 26418 12084 26424 12096
rect 26007 12056 26424 12084
rect 26007 12053 26019 12056
rect 25961 12047 26019 12053
rect 26418 12044 26424 12056
rect 26476 12044 26482 12096
rect 27798 12084 27804 12096
rect 27759 12056 27804 12084
rect 27798 12044 27804 12056
rect 27856 12044 27862 12096
rect 33318 12084 33324 12096
rect 33279 12056 33324 12084
rect 33318 12044 33324 12056
rect 33376 12044 33382 12096
rect 33686 12084 33692 12096
rect 33647 12056 33692 12084
rect 33686 12044 33692 12056
rect 33744 12044 33750 12096
rect 35618 12084 35624 12096
rect 35579 12056 35624 12084
rect 35618 12044 35624 12056
rect 35676 12044 35682 12096
rect 36725 12087 36783 12093
rect 36725 12053 36737 12087
rect 36771 12084 36783 12087
rect 37182 12084 37188 12096
rect 36771 12056 37188 12084
rect 36771 12053 36783 12056
rect 36725 12047 36783 12053
rect 37182 12044 37188 12056
rect 37240 12044 37246 12096
rect 1104 11994 38824 12016
rect 1104 11942 7648 11994
rect 7700 11942 7712 11994
rect 7764 11942 7776 11994
rect 7828 11942 7840 11994
rect 7892 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 34315 11994
rect 34367 11942 34379 11994
rect 34431 11942 34443 11994
rect 34495 11942 34507 11994
rect 34559 11942 38824 11994
rect 1104 11920 38824 11942
rect 5166 11840 5172 11892
rect 5224 11880 5230 11892
rect 5445 11883 5503 11889
rect 5445 11880 5457 11883
rect 5224 11852 5457 11880
rect 5224 11840 5230 11852
rect 5445 11849 5457 11852
rect 5491 11849 5503 11883
rect 5445 11843 5503 11849
rect 5626 11840 5632 11892
rect 5684 11880 5690 11892
rect 5813 11883 5871 11889
rect 5813 11880 5825 11883
rect 5684 11852 5825 11880
rect 5684 11840 5690 11852
rect 5813 11849 5825 11852
rect 5859 11849 5871 11883
rect 12066 11880 12072 11892
rect 12027 11852 12072 11880
rect 5813 11843 5871 11849
rect 12066 11840 12072 11852
rect 12124 11840 12130 11892
rect 13906 11880 13912 11892
rect 13867 11852 13912 11880
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 14737 11883 14795 11889
rect 14737 11849 14749 11883
rect 14783 11880 14795 11883
rect 14783 11852 15424 11880
rect 14783 11849 14795 11852
rect 14737 11843 14795 11849
rect 1578 11812 1584 11824
rect 1539 11784 1584 11812
rect 1578 11772 1584 11784
rect 1636 11772 1642 11824
rect 2593 11815 2651 11821
rect 2593 11781 2605 11815
rect 2639 11812 2651 11815
rect 3786 11812 3792 11824
rect 2639 11784 3792 11812
rect 2639 11781 2651 11784
rect 2593 11775 2651 11781
rect 3786 11772 3792 11784
rect 3844 11772 3850 11824
rect 4157 11815 4215 11821
rect 4157 11781 4169 11815
rect 4203 11812 4215 11815
rect 4614 11812 4620 11824
rect 4203 11784 4620 11812
rect 4203 11781 4215 11784
rect 4157 11775 4215 11781
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 9214 11812 9220 11824
rect 9175 11784 9220 11812
rect 9214 11772 9220 11784
rect 9272 11772 9278 11824
rect 12434 11772 12440 11824
rect 12492 11812 12498 11824
rect 12529 11815 12587 11821
rect 12529 11812 12541 11815
rect 12492 11784 12541 11812
rect 12492 11772 12498 11784
rect 12529 11781 12541 11784
rect 12575 11781 12587 11815
rect 12529 11775 12587 11781
rect 14921 11815 14979 11821
rect 14921 11781 14933 11815
rect 14967 11781 14979 11815
rect 14921 11775 14979 11781
rect 3510 11704 3516 11756
rect 3568 11744 3574 11756
rect 3973 11747 4031 11753
rect 3973 11744 3985 11747
rect 3568 11716 3985 11744
rect 3568 11704 3574 11716
rect 3973 11713 3985 11716
rect 4019 11744 4031 11747
rect 4522 11744 4528 11756
rect 4019 11716 4528 11744
rect 4019 11713 4031 11716
rect 3973 11707 4031 11713
rect 4522 11704 4528 11716
rect 4580 11704 4586 11756
rect 6270 11744 6276 11756
rect 5644 11716 6276 11744
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 1578 11676 1584 11688
rect 1443 11648 1584 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 1578 11636 1584 11648
rect 1636 11636 1642 11688
rect 5644 11685 5672 11716
rect 6270 11704 6276 11716
rect 6328 11704 6334 11756
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11744 7159 11747
rect 8662 11744 8668 11756
rect 7147 11716 8668 11744
rect 7147 11713 7159 11716
rect 7101 11707 7159 11713
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 9548 11716 9781 11744
rect 9548 11704 9554 11716
rect 9769 11713 9781 11716
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11744 11759 11747
rect 12894 11744 12900 11756
rect 11747 11716 12900 11744
rect 11747 11713 11759 11716
rect 11701 11707 11759 11713
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 5169 11679 5227 11685
rect 5169 11676 5181 11679
rect 4632 11648 5181 11676
rect 2041 11611 2099 11617
rect 2041 11577 2053 11611
rect 2087 11608 2099 11611
rect 2590 11608 2596 11620
rect 2087 11580 2596 11608
rect 2087 11577 2099 11580
rect 2041 11571 2099 11577
rect 2590 11568 2596 11580
rect 2648 11608 2654 11620
rect 2869 11611 2927 11617
rect 2869 11608 2881 11611
rect 2648 11580 2881 11608
rect 2648 11568 2654 11580
rect 2869 11577 2881 11580
rect 2915 11577 2927 11611
rect 3142 11608 3148 11620
rect 3103 11580 3148 11608
rect 2869 11571 2927 11577
rect 3142 11568 3148 11580
rect 3200 11568 3206 11620
rect 4632 11617 4660 11648
rect 5169 11645 5181 11648
rect 5215 11676 5227 11679
rect 5629 11679 5687 11685
rect 5629 11676 5641 11679
rect 5215 11648 5641 11676
rect 5215 11645 5227 11648
rect 5169 11639 5227 11645
rect 5629 11645 5641 11648
rect 5675 11645 5687 11679
rect 6822 11676 6828 11688
rect 6783 11648 6828 11676
rect 5629 11639 5687 11645
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 9122 11636 9128 11688
rect 9180 11676 9186 11688
rect 14936 11676 14964 11775
rect 15396 11756 15424 11852
rect 19518 11840 19524 11892
rect 19576 11880 19582 11892
rect 19613 11883 19671 11889
rect 19613 11880 19625 11883
rect 19576 11852 19625 11880
rect 19576 11840 19582 11852
rect 19613 11849 19625 11852
rect 19659 11880 19671 11883
rect 20901 11883 20959 11889
rect 20901 11880 20913 11883
rect 19659 11852 20913 11880
rect 19659 11849 19671 11852
rect 19613 11843 19671 11849
rect 20901 11849 20913 11852
rect 20947 11849 20959 11883
rect 21818 11880 21824 11892
rect 21779 11852 21824 11880
rect 20901 11843 20959 11849
rect 21818 11840 21824 11852
rect 21876 11840 21882 11892
rect 23290 11880 23296 11892
rect 23251 11852 23296 11880
rect 23290 11840 23296 11852
rect 23348 11840 23354 11892
rect 26510 11880 26516 11892
rect 25516 11852 26516 11880
rect 16482 11812 16488 11824
rect 16443 11784 16488 11812
rect 16482 11772 16488 11784
rect 16540 11772 16546 11824
rect 18141 11815 18199 11821
rect 18141 11812 18153 11815
rect 16960 11784 18153 11812
rect 15378 11744 15384 11756
rect 15339 11716 15384 11744
rect 15378 11704 15384 11716
rect 15436 11704 15442 11756
rect 15930 11704 15936 11756
rect 15988 11744 15994 11756
rect 16960 11753 16988 11784
rect 18141 11781 18153 11784
rect 18187 11781 18199 11815
rect 18141 11775 18199 11781
rect 20349 11815 20407 11821
rect 20349 11781 20361 11815
rect 20395 11812 20407 11815
rect 21726 11812 21732 11824
rect 20395 11784 21732 11812
rect 20395 11781 20407 11784
rect 20349 11775 20407 11781
rect 21726 11772 21732 11784
rect 21784 11772 21790 11824
rect 24029 11815 24087 11821
rect 24029 11781 24041 11815
rect 24075 11812 24087 11815
rect 25516 11812 25544 11852
rect 26510 11840 26516 11852
rect 26568 11840 26574 11892
rect 29454 11880 29460 11892
rect 29415 11852 29460 11880
rect 29454 11840 29460 11852
rect 29512 11840 29518 11892
rect 31754 11840 31760 11892
rect 31812 11880 31818 11892
rect 33229 11883 33287 11889
rect 31812 11852 31857 11880
rect 31812 11840 31818 11852
rect 33229 11849 33241 11883
rect 33275 11880 33287 11883
rect 33778 11880 33784 11892
rect 33275 11852 33784 11880
rect 33275 11849 33287 11852
rect 33229 11843 33287 11849
rect 33778 11840 33784 11852
rect 33836 11880 33842 11892
rect 34149 11883 34207 11889
rect 34149 11880 34161 11883
rect 33836 11852 34161 11880
rect 33836 11840 33842 11852
rect 34149 11849 34161 11852
rect 34195 11849 34207 11883
rect 34149 11843 34207 11849
rect 24075 11784 25544 11812
rect 26881 11815 26939 11821
rect 24075 11781 24087 11784
rect 24029 11775 24087 11781
rect 26881 11781 26893 11815
rect 26927 11812 26939 11815
rect 28350 11812 28356 11824
rect 26927 11784 28356 11812
rect 26927 11781 26939 11784
rect 26881 11775 26939 11781
rect 28350 11772 28356 11784
rect 28408 11772 28414 11824
rect 29089 11815 29147 11821
rect 29089 11781 29101 11815
rect 29135 11812 29147 11815
rect 29914 11812 29920 11824
rect 29135 11784 29920 11812
rect 29135 11781 29147 11784
rect 29089 11775 29147 11781
rect 29914 11772 29920 11784
rect 29972 11772 29978 11824
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 15988 11716 16957 11744
rect 15988 11704 15994 11716
rect 16945 11713 16957 11716
rect 16991 11713 17003 11747
rect 21266 11744 21272 11756
rect 21227 11716 21272 11744
rect 16945 11707 17003 11713
rect 21266 11704 21272 11716
rect 21324 11704 21330 11756
rect 22370 11744 22376 11756
rect 22331 11716 22376 11744
rect 22370 11704 22376 11716
rect 22428 11704 22434 11756
rect 24578 11744 24584 11756
rect 24539 11716 24584 11744
rect 24578 11704 24584 11716
rect 24636 11704 24642 11756
rect 28169 11747 28227 11753
rect 28169 11713 28181 11747
rect 28215 11744 28227 11747
rect 28902 11744 28908 11756
rect 28215 11716 28908 11744
rect 28215 11713 28227 11716
rect 28169 11707 28227 11713
rect 28902 11704 28908 11716
rect 28960 11704 28966 11756
rect 33686 11744 33692 11756
rect 33647 11716 33692 11744
rect 33686 11704 33692 11716
rect 33744 11704 33750 11756
rect 16298 11676 16304 11688
rect 9180 11648 9720 11676
rect 14936 11648 16304 11676
rect 9180 11636 9186 11648
rect 4617 11611 4675 11617
rect 4617 11577 4629 11611
rect 4663 11577 4675 11611
rect 4617 11571 4675 11577
rect 4706 11568 4712 11620
rect 4764 11608 4770 11620
rect 9493 11611 9551 11617
rect 4764 11580 4809 11608
rect 4764 11568 4770 11580
rect 9493 11577 9505 11611
rect 9539 11608 9551 11611
rect 9582 11608 9588 11620
rect 9539 11580 9588 11608
rect 9539 11577 9551 11580
rect 9493 11571 9551 11577
rect 2409 11543 2467 11549
rect 2409 11509 2421 11543
rect 2455 11540 2467 11543
rect 3053 11543 3111 11549
rect 3053 11540 3065 11543
rect 2455 11512 3065 11540
rect 2455 11509 2467 11512
rect 2409 11503 2467 11509
rect 3053 11509 3065 11512
rect 3099 11540 3111 11543
rect 3326 11540 3332 11552
rect 3099 11512 3332 11540
rect 3099 11509 3111 11512
rect 3053 11503 3111 11509
rect 3326 11500 3332 11512
rect 3384 11500 3390 11552
rect 3418 11500 3424 11552
rect 3476 11540 3482 11552
rect 3513 11543 3571 11549
rect 3513 11540 3525 11543
rect 3476 11512 3525 11540
rect 3476 11500 3482 11512
rect 3513 11509 3525 11512
rect 3559 11509 3571 11543
rect 3513 11503 3571 11509
rect 6270 11500 6276 11552
rect 6328 11540 6334 11552
rect 6549 11543 6607 11549
rect 6549 11540 6561 11543
rect 6328 11512 6561 11540
rect 6328 11500 6334 11512
rect 6549 11509 6561 11512
rect 6595 11509 6607 11543
rect 6549 11503 6607 11509
rect 7374 11500 7380 11552
rect 7432 11540 7438 11552
rect 7653 11543 7711 11549
rect 7653 11540 7665 11543
rect 7432 11512 7665 11540
rect 7432 11500 7438 11512
rect 7653 11509 7665 11512
rect 7699 11540 7711 11543
rect 8018 11540 8024 11552
rect 7699 11512 8024 11540
rect 7699 11509 7711 11512
rect 7653 11503 7711 11509
rect 8018 11500 8024 11512
rect 8076 11500 8082 11552
rect 8938 11540 8944 11552
rect 8899 11512 8944 11540
rect 8938 11500 8944 11512
rect 8996 11540 9002 11552
rect 9508 11540 9536 11571
rect 9582 11568 9588 11580
rect 9640 11568 9646 11620
rect 9692 11617 9720 11648
rect 16298 11636 16304 11648
rect 16356 11676 16362 11688
rect 17862 11676 17868 11688
rect 16356 11648 16988 11676
rect 17775 11648 17868 11676
rect 16356 11636 16362 11648
rect 9677 11611 9735 11617
rect 9677 11577 9689 11611
rect 9723 11608 9735 11611
rect 9858 11608 9864 11620
rect 9723 11580 9864 11608
rect 9723 11577 9735 11580
rect 9677 11571 9735 11577
rect 9858 11568 9864 11580
rect 9916 11568 9922 11620
rect 11333 11611 11391 11617
rect 11333 11577 11345 11611
rect 11379 11608 11391 11611
rect 12710 11608 12716 11620
rect 11379 11580 12716 11608
rect 11379 11577 11391 11580
rect 11333 11571 11391 11577
rect 12710 11568 12716 11580
rect 12768 11568 12774 11620
rect 12986 11608 12992 11620
rect 12947 11580 12992 11608
rect 12986 11568 12992 11580
rect 13044 11568 13050 11620
rect 13081 11611 13139 11617
rect 13081 11577 13093 11611
rect 13127 11577 13139 11611
rect 13081 11571 13139 11577
rect 8996 11512 9536 11540
rect 13096 11540 13124 11571
rect 15102 11568 15108 11620
rect 15160 11608 15166 11620
rect 16960 11617 16988 11648
rect 17862 11636 17868 11648
rect 17920 11676 17926 11688
rect 22922 11676 22928 11688
rect 17920 11648 18644 11676
rect 22883 11648 22928 11676
rect 17920 11636 17926 11648
rect 18616 11620 18644 11648
rect 22922 11636 22928 11648
rect 22980 11636 22986 11688
rect 24026 11636 24032 11688
rect 24084 11676 24090 11688
rect 24305 11679 24363 11685
rect 24305 11676 24317 11679
rect 24084 11648 24317 11676
rect 24084 11636 24090 11648
rect 24305 11645 24317 11648
rect 24351 11645 24363 11679
rect 25501 11679 25559 11685
rect 25501 11676 25513 11679
rect 24305 11639 24363 11645
rect 25332 11648 25513 11676
rect 15473 11611 15531 11617
rect 15473 11608 15485 11611
rect 15160 11580 15485 11608
rect 15160 11568 15166 11580
rect 15473 11577 15485 11580
rect 15519 11577 15531 11611
rect 15473 11571 15531 11577
rect 16945 11611 17003 11617
rect 16945 11577 16957 11611
rect 16991 11577 17003 11611
rect 16945 11571 17003 11577
rect 17037 11611 17095 11617
rect 17037 11577 17049 11611
rect 17083 11608 17095 11611
rect 17126 11608 17132 11620
rect 17083 11580 17132 11608
rect 17083 11577 17095 11580
rect 17037 11571 17095 11577
rect 13446 11540 13452 11552
rect 13096 11512 13452 11540
rect 8996 11500 9002 11512
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 15194 11500 15200 11552
rect 15252 11540 15258 11552
rect 15381 11543 15439 11549
rect 15381 11540 15393 11543
rect 15252 11512 15393 11540
rect 15252 11500 15258 11512
rect 15381 11509 15393 11512
rect 15427 11509 15439 11543
rect 15381 11503 15439 11509
rect 15933 11543 15991 11549
rect 15933 11509 15945 11543
rect 15979 11540 15991 11543
rect 16209 11543 16267 11549
rect 16209 11540 16221 11543
rect 15979 11512 16221 11540
rect 15979 11509 15991 11512
rect 15933 11503 15991 11509
rect 16209 11509 16221 11512
rect 16255 11540 16267 11543
rect 17052 11540 17080 11571
rect 17126 11568 17132 11580
rect 17184 11568 17190 11620
rect 17494 11608 17500 11620
rect 17407 11580 17500 11608
rect 17494 11568 17500 11580
rect 17552 11608 17558 11620
rect 18417 11611 18475 11617
rect 18417 11608 18429 11611
rect 17552 11580 18429 11608
rect 17552 11568 17558 11580
rect 18417 11577 18429 11580
rect 18463 11577 18475 11611
rect 18598 11608 18604 11620
rect 18559 11580 18604 11608
rect 18417 11571 18475 11577
rect 18598 11568 18604 11580
rect 18656 11568 18662 11620
rect 18690 11568 18696 11620
rect 18748 11608 18754 11620
rect 19061 11611 19119 11617
rect 19061 11608 19073 11611
rect 18748 11580 19073 11608
rect 18748 11568 18754 11580
rect 19061 11577 19073 11580
rect 19107 11577 19119 11611
rect 19061 11571 19119 11577
rect 19981 11611 20039 11617
rect 19981 11577 19993 11611
rect 20027 11608 20039 11611
rect 20717 11611 20775 11617
rect 20027 11580 20668 11608
rect 20027 11577 20039 11580
rect 19981 11571 20039 11577
rect 16255 11512 17080 11540
rect 20640 11540 20668 11580
rect 20717 11577 20729 11611
rect 20763 11608 20775 11611
rect 21450 11608 21456 11620
rect 20763 11580 21456 11608
rect 20763 11577 20775 11580
rect 20717 11571 20775 11577
rect 21450 11568 21456 11580
rect 21508 11568 21514 11620
rect 21818 11568 21824 11620
rect 21876 11608 21882 11620
rect 22370 11608 22376 11620
rect 21876 11580 22376 11608
rect 21876 11568 21882 11580
rect 22370 11568 22376 11580
rect 22428 11568 22434 11620
rect 24394 11568 24400 11620
rect 24452 11608 24458 11620
rect 24489 11611 24547 11617
rect 24489 11608 24501 11611
rect 24452 11580 24501 11608
rect 24452 11568 24458 11580
rect 24489 11577 24501 11580
rect 24535 11577 24547 11611
rect 24489 11571 24547 11577
rect 25332 11552 25360 11648
rect 25501 11645 25513 11648
rect 25547 11645 25559 11679
rect 25501 11639 25559 11645
rect 29178 11636 29184 11688
rect 29236 11676 29242 11688
rect 29273 11679 29331 11685
rect 29273 11676 29285 11679
rect 29236 11648 29285 11676
rect 29236 11636 29242 11648
rect 29273 11645 29285 11648
rect 29319 11676 29331 11679
rect 29825 11679 29883 11685
rect 29825 11676 29837 11679
rect 29319 11648 29837 11676
rect 29319 11645 29331 11648
rect 29273 11639 29331 11645
rect 29825 11645 29837 11648
rect 29871 11645 29883 11679
rect 30374 11676 30380 11688
rect 30335 11648 30380 11676
rect 29825 11639 29883 11645
rect 30374 11636 30380 11648
rect 30432 11636 30438 11688
rect 30650 11685 30656 11688
rect 30644 11676 30656 11685
rect 30611 11648 30656 11676
rect 30644 11639 30656 11648
rect 30650 11636 30656 11639
rect 30708 11636 30714 11688
rect 35250 11636 35256 11688
rect 35308 11676 35314 11688
rect 35437 11679 35495 11685
rect 35437 11676 35449 11679
rect 35308 11648 35449 11676
rect 35308 11636 35314 11648
rect 35437 11645 35449 11648
rect 35483 11676 35495 11679
rect 35989 11679 36047 11685
rect 35989 11676 36001 11679
rect 35483 11648 36001 11676
rect 35483 11645 35495 11648
rect 35437 11639 35495 11645
rect 35989 11645 36001 11648
rect 36035 11645 36047 11679
rect 35989 11639 36047 11645
rect 36262 11636 36268 11688
rect 36320 11676 36326 11688
rect 36541 11679 36599 11685
rect 36541 11676 36553 11679
rect 36320 11648 36553 11676
rect 36320 11636 36326 11648
rect 36541 11645 36553 11648
rect 36587 11676 36599 11679
rect 37093 11679 37151 11685
rect 37093 11676 37105 11679
rect 36587 11648 37105 11676
rect 36587 11645 36599 11648
rect 36541 11639 36599 11645
rect 37093 11645 37105 11648
rect 37139 11645 37151 11679
rect 37093 11639 37151 11645
rect 25774 11617 25780 11620
rect 25768 11608 25780 11617
rect 25735 11580 25780 11608
rect 25768 11571 25780 11580
rect 25774 11568 25780 11571
rect 25832 11568 25838 11620
rect 27801 11611 27859 11617
rect 27801 11577 27813 11611
rect 27847 11608 27859 11611
rect 28258 11608 28264 11620
rect 27847 11580 28264 11608
rect 27847 11577 27859 11580
rect 27801 11571 27859 11577
rect 28258 11568 28264 11580
rect 28316 11608 28322 11620
rect 28902 11608 28908 11620
rect 28316 11580 28908 11608
rect 28316 11568 28322 11580
rect 28902 11568 28908 11580
rect 28960 11568 28966 11620
rect 32416 11580 32996 11608
rect 32416 11552 32444 11580
rect 21361 11543 21419 11549
rect 21361 11540 21373 11543
rect 20640 11512 21373 11540
rect 16255 11509 16267 11512
rect 16209 11503 16267 11509
rect 21361 11509 21373 11512
rect 21407 11540 21419 11543
rect 21726 11540 21732 11552
rect 21407 11512 21732 11540
rect 21407 11509 21419 11512
rect 21361 11503 21419 11509
rect 21726 11500 21732 11512
rect 21784 11500 21790 11552
rect 22186 11540 22192 11552
rect 22147 11512 22192 11540
rect 22186 11500 22192 11512
rect 22244 11500 22250 11552
rect 24946 11540 24952 11552
rect 24907 11512 24952 11540
rect 24946 11500 24952 11512
rect 25004 11500 25010 11552
rect 25314 11540 25320 11552
rect 25275 11512 25320 11540
rect 25314 11500 25320 11512
rect 25372 11500 25378 11552
rect 28721 11543 28779 11549
rect 28721 11509 28733 11543
rect 28767 11540 28779 11543
rect 28810 11540 28816 11552
rect 28767 11512 28816 11540
rect 28767 11509 28779 11512
rect 28721 11503 28779 11509
rect 28810 11500 28816 11512
rect 28868 11500 28874 11552
rect 30285 11543 30343 11549
rect 30285 11509 30297 11543
rect 30331 11540 30343 11543
rect 30558 11540 30564 11552
rect 30331 11512 30564 11540
rect 30331 11509 30343 11512
rect 30285 11503 30343 11509
rect 30558 11500 30564 11512
rect 30616 11500 30622 11552
rect 32398 11540 32404 11552
rect 32359 11512 32404 11540
rect 32398 11500 32404 11512
rect 32456 11500 32462 11552
rect 32674 11540 32680 11552
rect 32635 11512 32680 11540
rect 32674 11500 32680 11512
rect 32732 11500 32738 11552
rect 32968 11540 32996 11580
rect 33318 11568 33324 11620
rect 33376 11608 33382 11620
rect 33778 11608 33784 11620
rect 33376 11580 33784 11608
rect 33376 11568 33382 11580
rect 33778 11568 33784 11580
rect 33836 11568 33842 11620
rect 33689 11543 33747 11549
rect 33689 11540 33701 11543
rect 32968 11512 33701 11540
rect 33689 11509 33701 11512
rect 33735 11509 33747 11543
rect 34698 11540 34704 11552
rect 34659 11512 34704 11540
rect 33689 11503 33747 11509
rect 34698 11500 34704 11512
rect 34756 11500 34762 11552
rect 34974 11500 34980 11552
rect 35032 11540 35038 11552
rect 35253 11543 35311 11549
rect 35253 11540 35265 11543
rect 35032 11512 35265 11540
rect 35032 11500 35038 11512
rect 35253 11509 35265 11512
rect 35299 11509 35311 11543
rect 35253 11503 35311 11509
rect 35621 11543 35679 11549
rect 35621 11509 35633 11543
rect 35667 11540 35679 11543
rect 35802 11540 35808 11552
rect 35667 11512 35808 11540
rect 35667 11509 35679 11512
rect 35621 11503 35679 11509
rect 35802 11500 35808 11512
rect 35860 11500 35866 11552
rect 36446 11540 36452 11552
rect 36407 11512 36452 11540
rect 36446 11500 36452 11512
rect 36504 11500 36510 11552
rect 36722 11540 36728 11552
rect 36683 11512 36728 11540
rect 36722 11500 36728 11512
rect 36780 11500 36786 11552
rect 1104 11450 38824 11472
rect 1104 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 27648 11450
rect 27700 11398 27712 11450
rect 27764 11398 27776 11450
rect 27828 11398 27840 11450
rect 27892 11398 38824 11450
rect 1104 11376 38824 11398
rect 2222 11296 2228 11348
rect 2280 11336 2286 11348
rect 2593 11339 2651 11345
rect 2593 11336 2605 11339
rect 2280 11308 2605 11336
rect 2280 11296 2286 11308
rect 2593 11305 2605 11308
rect 2639 11336 2651 11339
rect 3786 11336 3792 11348
rect 2639 11308 3556 11336
rect 3747 11308 3792 11336
rect 2639 11305 2651 11308
rect 2593 11299 2651 11305
rect 2409 11203 2467 11209
rect 2409 11169 2421 11203
rect 2455 11169 2467 11203
rect 2409 11163 2467 11169
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 1673 11135 1731 11141
rect 1673 11132 1685 11135
rect 1636 11104 1685 11132
rect 1636 11092 1642 11104
rect 1673 11101 1685 11104
rect 1719 11132 1731 11135
rect 2314 11132 2320 11144
rect 1719 11104 2320 11132
rect 1719 11101 1731 11104
rect 1673 11095 1731 11101
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 2130 11064 2136 11076
rect 2091 11036 2136 11064
rect 2130 11024 2136 11036
rect 2188 11024 2194 11076
rect 2424 10996 2452 11163
rect 2498 11160 2504 11212
rect 2556 11200 2562 11212
rect 3421 11203 3479 11209
rect 3421 11200 3433 11203
rect 2556 11172 3433 11200
rect 2556 11160 2562 11172
rect 3421 11169 3433 11172
rect 3467 11169 3479 11203
rect 3528 11200 3556 11308
rect 3786 11296 3792 11308
rect 3844 11336 3850 11348
rect 4617 11339 4675 11345
rect 4617 11336 4629 11339
rect 3844 11308 4629 11336
rect 3844 11296 3850 11308
rect 4617 11305 4629 11308
rect 4663 11305 4675 11339
rect 9122 11336 9128 11348
rect 9083 11308 9128 11336
rect 4617 11299 4675 11305
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 12069 11339 12127 11345
rect 12069 11305 12081 11339
rect 12115 11336 12127 11339
rect 12342 11336 12348 11348
rect 12115 11308 12348 11336
rect 12115 11305 12127 11308
rect 12069 11299 12127 11305
rect 12342 11296 12348 11308
rect 12400 11296 12406 11348
rect 15930 11336 15936 11348
rect 15891 11308 15936 11336
rect 15930 11296 15936 11308
rect 15988 11296 15994 11348
rect 17034 11336 17040 11348
rect 16995 11308 17040 11336
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 20717 11339 20775 11345
rect 20717 11305 20729 11339
rect 20763 11336 20775 11339
rect 21542 11336 21548 11348
rect 20763 11308 21548 11336
rect 20763 11305 20775 11308
rect 20717 11299 20775 11305
rect 21542 11296 21548 11308
rect 21600 11296 21606 11348
rect 22741 11339 22799 11345
rect 22741 11305 22753 11339
rect 22787 11305 22799 11339
rect 22741 11299 22799 11305
rect 4338 11228 4344 11280
rect 4396 11268 4402 11280
rect 4706 11268 4712 11280
rect 4396 11240 4712 11268
rect 4396 11228 4402 11240
rect 4706 11228 4712 11240
rect 4764 11228 4770 11280
rect 9214 11228 9220 11280
rect 9272 11268 9278 11280
rect 10229 11271 10287 11277
rect 10229 11268 10241 11271
rect 9272 11240 10241 11268
rect 9272 11228 9278 11240
rect 10229 11237 10241 11240
rect 10275 11237 10287 11271
rect 10229 11231 10287 11237
rect 16114 11228 16120 11280
rect 16172 11268 16178 11280
rect 16577 11271 16635 11277
rect 16577 11268 16589 11271
rect 16172 11240 16589 11268
rect 16172 11228 16178 11240
rect 16577 11237 16589 11240
rect 16623 11237 16635 11271
rect 16577 11231 16635 11237
rect 17126 11228 17132 11280
rect 17184 11268 17190 11280
rect 17862 11277 17868 11280
rect 17834 11271 17868 11277
rect 17834 11268 17846 11271
rect 17184 11240 17846 11268
rect 17184 11228 17190 11240
rect 17834 11237 17846 11240
rect 17920 11268 17926 11280
rect 21269 11271 21327 11277
rect 17920 11240 17982 11268
rect 17834 11231 17868 11237
rect 17862 11228 17868 11231
rect 17920 11228 17926 11240
rect 21269 11237 21281 11271
rect 21315 11268 21327 11271
rect 22370 11268 22376 11280
rect 21315 11240 22376 11268
rect 21315 11237 21327 11240
rect 21269 11231 21327 11237
rect 22370 11228 22376 11240
rect 22428 11268 22434 11280
rect 22756 11268 22784 11299
rect 25130 11296 25136 11348
rect 25188 11336 25194 11348
rect 25225 11339 25283 11345
rect 25225 11336 25237 11339
rect 25188 11308 25237 11336
rect 25188 11296 25194 11308
rect 25225 11305 25237 11308
rect 25271 11336 25283 11339
rect 25774 11336 25780 11348
rect 25271 11308 25780 11336
rect 25271 11305 25283 11308
rect 25225 11299 25283 11305
rect 25774 11296 25780 11308
rect 25832 11296 25838 11348
rect 26237 11339 26295 11345
rect 26237 11305 26249 11339
rect 26283 11336 26295 11339
rect 26326 11336 26332 11348
rect 26283 11308 26332 11336
rect 26283 11305 26295 11308
rect 26237 11299 26295 11305
rect 26326 11296 26332 11308
rect 26384 11296 26390 11348
rect 28350 11296 28356 11348
rect 28408 11336 28414 11348
rect 28445 11339 28503 11345
rect 28445 11336 28457 11339
rect 28408 11308 28457 11336
rect 28408 11296 28414 11308
rect 28445 11305 28457 11308
rect 28491 11336 28503 11339
rect 28813 11339 28871 11345
rect 28813 11336 28825 11339
rect 28491 11308 28825 11336
rect 28491 11305 28503 11308
rect 28445 11299 28503 11305
rect 28813 11305 28825 11308
rect 28859 11336 28871 11339
rect 29086 11336 29092 11348
rect 28859 11308 29092 11336
rect 28859 11305 28871 11308
rect 28813 11299 28871 11305
rect 29086 11296 29092 11308
rect 29144 11296 29150 11348
rect 29822 11296 29828 11348
rect 29880 11336 29886 11348
rect 30745 11339 30803 11345
rect 30745 11336 30757 11339
rect 29880 11308 30757 11336
rect 29880 11296 29886 11308
rect 30745 11305 30757 11308
rect 30791 11305 30803 11339
rect 30745 11299 30803 11305
rect 31113 11339 31171 11345
rect 31113 11305 31125 11339
rect 31159 11336 31171 11339
rect 35894 11336 35900 11348
rect 31159 11308 35900 11336
rect 31159 11305 31171 11308
rect 31113 11299 31171 11305
rect 35894 11296 35900 11308
rect 35952 11296 35958 11348
rect 22428 11240 22784 11268
rect 22428 11228 22434 11240
rect 5077 11203 5135 11209
rect 5077 11200 5089 11203
rect 3528 11172 5089 11200
rect 3421 11163 3479 11169
rect 5077 11169 5089 11172
rect 5123 11169 5135 11203
rect 5077 11163 5135 11169
rect 5629 11203 5687 11209
rect 5629 11169 5641 11203
rect 5675 11200 5687 11203
rect 6178 11200 6184 11212
rect 5675 11172 6184 11200
rect 5675 11169 5687 11172
rect 5629 11163 5687 11169
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 10042 11200 10048 11212
rect 10003 11172 10048 11200
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 12342 11160 12348 11212
rect 12400 11200 12406 11212
rect 12509 11203 12567 11209
rect 12509 11200 12521 11203
rect 12400 11172 12521 11200
rect 12400 11160 12406 11172
rect 12509 11169 12521 11172
rect 12555 11169 12567 11203
rect 12509 11163 12567 11169
rect 21628 11203 21686 11209
rect 21628 11169 21640 11203
rect 21674 11200 21686 11203
rect 22186 11200 22192 11212
rect 21674 11172 22192 11200
rect 21674 11169 21686 11172
rect 21628 11163 21686 11169
rect 22186 11160 22192 11172
rect 22244 11200 22250 11212
rect 22646 11200 22652 11212
rect 22244 11172 22652 11200
rect 22244 11160 22250 11172
rect 22646 11160 22652 11172
rect 22704 11160 22710 11212
rect 22756 11200 22784 11240
rect 22922 11228 22928 11280
rect 22980 11268 22986 11280
rect 25866 11268 25872 11280
rect 22980 11240 25872 11268
rect 22980 11228 22986 11240
rect 25866 11228 25872 11240
rect 25924 11228 25930 11280
rect 26780 11271 26838 11277
rect 26780 11237 26792 11271
rect 26826 11268 26838 11271
rect 26970 11268 26976 11280
rect 26826 11240 26976 11268
rect 26826 11237 26838 11240
rect 26780 11231 26838 11237
rect 26970 11228 26976 11240
rect 27028 11228 27034 11280
rect 28626 11228 28632 11280
rect 28684 11268 28690 11280
rect 29549 11271 29607 11277
rect 29549 11268 29561 11271
rect 28684 11240 29561 11268
rect 28684 11228 28690 11240
rect 29549 11237 29561 11240
rect 29595 11237 29607 11271
rect 29549 11231 29607 11237
rect 32401 11271 32459 11277
rect 32401 11237 32413 11271
rect 32447 11268 32459 11271
rect 33413 11271 33471 11277
rect 33413 11268 33425 11271
rect 32447 11240 33425 11268
rect 32447 11237 32459 11240
rect 32401 11231 32459 11237
rect 33413 11237 33425 11240
rect 33459 11268 33471 11271
rect 34422 11268 34428 11280
rect 33459 11240 34428 11268
rect 33459 11237 33471 11240
rect 33413 11231 33471 11237
rect 34422 11228 34428 11240
rect 34480 11228 34486 11280
rect 35161 11271 35219 11277
rect 35161 11237 35173 11271
rect 35207 11268 35219 11271
rect 35710 11268 35716 11280
rect 35207 11240 35716 11268
rect 35207 11237 35219 11240
rect 35161 11231 35219 11237
rect 35710 11228 35716 11240
rect 35768 11228 35774 11280
rect 24118 11209 24124 11212
rect 24112 11200 24124 11209
rect 22756 11172 24124 11200
rect 24112 11163 24124 11172
rect 24118 11160 24124 11163
rect 24176 11160 24182 11212
rect 24670 11160 24676 11212
rect 24728 11200 24734 11212
rect 27982 11200 27988 11212
rect 24728 11172 27988 11200
rect 24728 11160 24734 11172
rect 27982 11160 27988 11172
rect 28040 11160 28046 11212
rect 29178 11160 29184 11212
rect 29236 11200 29242 11212
rect 29365 11203 29423 11209
rect 29365 11200 29377 11203
rect 29236 11172 29377 11200
rect 29236 11160 29242 11172
rect 29365 11169 29377 11172
rect 29411 11169 29423 11203
rect 30926 11200 30932 11212
rect 30887 11172 30932 11200
rect 29365 11163 29423 11169
rect 30926 11160 30932 11172
rect 30984 11160 30990 11212
rect 34698 11160 34704 11212
rect 34756 11200 34762 11212
rect 35253 11203 35311 11209
rect 35253 11200 35265 11203
rect 34756 11172 35265 11200
rect 34756 11160 34762 11172
rect 35253 11169 35265 11172
rect 35299 11200 35311 11203
rect 35621 11203 35679 11209
rect 35621 11200 35633 11203
rect 35299 11172 35633 11200
rect 35299 11169 35311 11172
rect 35253 11163 35311 11169
rect 35621 11169 35633 11172
rect 35667 11169 35679 11203
rect 36170 11200 36176 11212
rect 36131 11172 36176 11200
rect 35621 11163 35679 11169
rect 36170 11160 36176 11172
rect 36228 11160 36234 11212
rect 2682 11092 2688 11144
rect 2740 11132 2746 11144
rect 2961 11135 3019 11141
rect 2740 11104 2785 11132
rect 2740 11092 2746 11104
rect 2961 11101 2973 11135
rect 3007 11132 3019 11135
rect 3697 11135 3755 11141
rect 3697 11132 3709 11135
rect 3007 11104 3709 11132
rect 3007 11101 3019 11104
rect 2961 11095 3019 11101
rect 3697 11101 3709 11104
rect 3743 11101 3755 11135
rect 3697 11095 3755 11101
rect 3878 11092 3884 11144
rect 3936 11132 3942 11144
rect 4338 11132 4344 11144
rect 3936 11104 4344 11132
rect 3936 11092 3942 11104
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11132 4675 11135
rect 4706 11132 4712 11144
rect 4663 11104 4712 11132
rect 4663 11101 4675 11104
rect 4617 11095 4675 11101
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 8573 11135 8631 11141
rect 8573 11101 8585 11135
rect 8619 11132 8631 11135
rect 9582 11132 9588 11144
rect 8619 11104 9588 11132
rect 8619 11101 8631 11104
rect 8573 11095 8631 11101
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 10318 11132 10324 11144
rect 10279 11104 10324 11132
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 12158 11092 12164 11144
rect 12216 11132 12222 11144
rect 12253 11135 12311 11141
rect 12253 11132 12265 11135
rect 12216 11104 12265 11132
rect 12216 11092 12222 11104
rect 12253 11101 12265 11104
rect 12299 11101 12311 11135
rect 16482 11132 16488 11144
rect 16443 11104 16488 11132
rect 12253 11095 12311 11101
rect 16482 11092 16488 11104
rect 16540 11092 16546 11144
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11101 16727 11135
rect 16669 11095 16727 11101
rect 5810 11064 5816 11076
rect 5771 11036 5816 11064
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 9766 11064 9772 11076
rect 9727 11036 9772 11064
rect 9766 11024 9772 11036
rect 9824 11024 9830 11076
rect 14921 11067 14979 11073
rect 14921 11033 14933 11067
rect 14967 11064 14979 11067
rect 15194 11064 15200 11076
rect 14967 11036 15200 11064
rect 14967 11033 14979 11036
rect 14921 11027 14979 11033
rect 15194 11024 15200 11036
rect 15252 11024 15258 11076
rect 16117 11067 16175 11073
rect 16117 11033 16129 11067
rect 16163 11064 16175 11067
rect 16206 11064 16212 11076
rect 16163 11036 16212 11064
rect 16163 11033 16175 11036
rect 16117 11027 16175 11033
rect 16206 11024 16212 11036
rect 16264 11024 16270 11076
rect 16684 11064 16712 11095
rect 17310 11092 17316 11144
rect 17368 11132 17374 11144
rect 17589 11135 17647 11141
rect 17589 11132 17601 11135
rect 17368 11104 17601 11132
rect 17368 11092 17374 11104
rect 17589 11101 17601 11104
rect 17635 11101 17647 11135
rect 17589 11095 17647 11101
rect 21266 11092 21272 11144
rect 21324 11132 21330 11144
rect 21361 11135 21419 11141
rect 21361 11132 21373 11135
rect 21324 11104 21373 11132
rect 21324 11092 21330 11104
rect 21361 11101 21373 11104
rect 21407 11101 21419 11135
rect 21361 11095 21419 11101
rect 23750 11092 23756 11144
rect 23808 11132 23814 11144
rect 23845 11135 23903 11141
rect 23845 11132 23857 11135
rect 23808 11104 23857 11132
rect 23808 11092 23814 11104
rect 23845 11101 23857 11104
rect 23891 11101 23903 11135
rect 23845 11095 23903 11101
rect 25314 11092 25320 11144
rect 25372 11132 25378 11144
rect 26510 11132 26516 11144
rect 25372 11104 26516 11132
rect 25372 11092 25378 11104
rect 26510 11092 26516 11104
rect 26568 11092 26574 11144
rect 29641 11135 29699 11141
rect 29641 11132 29653 11135
rect 28920 11104 29653 11132
rect 27890 11064 27896 11076
rect 16500 11036 17632 11064
rect 27851 11036 27896 11064
rect 2961 10999 3019 11005
rect 2961 10996 2973 10999
rect 2424 10968 2973 10996
rect 2961 10965 2973 10968
rect 3007 10965 3019 10999
rect 3142 10996 3148 11008
rect 3103 10968 3148 10996
rect 2961 10959 3019 10965
rect 3142 10956 3148 10968
rect 3200 10956 3206 11008
rect 3697 10999 3755 11005
rect 3697 10965 3709 10999
rect 3743 10996 3755 10999
rect 4157 10999 4215 11005
rect 4157 10996 4169 10999
rect 3743 10968 4169 10996
rect 3743 10965 3755 10968
rect 3697 10959 3755 10965
rect 4157 10965 4169 10968
rect 4203 10996 4215 10999
rect 5445 10999 5503 11005
rect 5445 10996 5457 10999
rect 4203 10968 5457 10996
rect 4203 10965 4215 10968
rect 4157 10959 4215 10965
rect 5445 10965 5457 10968
rect 5491 10965 5503 10999
rect 5445 10959 5503 10965
rect 6917 10999 6975 11005
rect 6917 10965 6929 10999
rect 6963 10996 6975 10999
rect 7190 10996 7196 11008
rect 6963 10968 7196 10996
rect 6963 10965 6975 10968
rect 6917 10959 6975 10965
rect 7190 10956 7196 10968
rect 7248 10956 7254 11008
rect 13630 10996 13636 11008
rect 13591 10968 13636 10996
rect 13630 10956 13636 10968
rect 13688 10956 13694 11008
rect 16390 10956 16396 11008
rect 16448 10996 16454 11008
rect 16500 10996 16528 11036
rect 16448 10968 16528 10996
rect 17604 10996 17632 11036
rect 27890 11024 27896 11036
rect 27948 11024 27954 11076
rect 18690 10996 18696 11008
rect 17604 10968 18696 10996
rect 16448 10956 16454 10968
rect 18690 10956 18696 10968
rect 18748 10996 18754 11008
rect 18969 10999 19027 11005
rect 18969 10996 18981 10999
rect 18748 10968 18981 10996
rect 18748 10956 18754 10968
rect 18969 10965 18981 10968
rect 19015 10965 19027 10999
rect 18969 10959 19027 10965
rect 20162 10956 20168 11008
rect 20220 10996 20226 11008
rect 22462 10996 22468 11008
rect 20220 10968 22468 10996
rect 20220 10956 20226 10968
rect 22462 10956 22468 10968
rect 22520 10956 22526 11008
rect 23290 10996 23296 11008
rect 23251 10968 23296 10996
rect 23290 10956 23296 10968
rect 23348 10956 23354 11008
rect 23753 10999 23811 11005
rect 23753 10965 23765 10999
rect 23799 10996 23811 10999
rect 23842 10996 23848 11008
rect 23799 10968 23848 10996
rect 23799 10965 23811 10968
rect 23753 10959 23811 10965
rect 23842 10956 23848 10968
rect 23900 10956 23906 11008
rect 28350 10956 28356 11008
rect 28408 10996 28414 11008
rect 28920 10996 28948 11104
rect 29641 11101 29653 11104
rect 29687 11101 29699 11135
rect 29641 11095 29699 11101
rect 32769 11135 32827 11141
rect 32769 11101 32781 11135
rect 32815 11132 32827 11135
rect 33042 11132 33048 11144
rect 32815 11104 33048 11132
rect 32815 11101 32827 11104
rect 32769 11095 32827 11101
rect 33042 11092 33048 11104
rect 33100 11092 33106 11144
rect 33318 11132 33324 11144
rect 33279 11104 33324 11132
rect 33318 11092 33324 11104
rect 33376 11092 33382 11144
rect 33502 11132 33508 11144
rect 33463 11104 33508 11132
rect 33502 11092 33508 11104
rect 33560 11092 33566 11144
rect 34517 11135 34575 11141
rect 34517 11101 34529 11135
rect 34563 11132 34575 11135
rect 35158 11132 35164 11144
rect 34563 11104 35164 11132
rect 34563 11101 34575 11104
rect 34517 11095 34575 11101
rect 35158 11092 35164 11104
rect 35216 11092 35222 11144
rect 28994 11024 29000 11076
rect 29052 11064 29058 11076
rect 29089 11067 29147 11073
rect 29089 11064 29101 11067
rect 29052 11036 29101 11064
rect 29052 11024 29058 11036
rect 29089 11033 29101 11036
rect 29135 11033 29147 11067
rect 30374 11064 30380 11076
rect 29089 11027 29147 11033
rect 30024 11036 30380 11064
rect 28408 10968 28948 10996
rect 28408 10956 28414 10968
rect 29362 10956 29368 11008
rect 29420 10996 29426 11008
rect 30024 11005 30052 11036
rect 30374 11024 30380 11036
rect 30432 11024 30438 11076
rect 32398 11024 32404 11076
rect 32456 11064 32462 11076
rect 32953 11067 33011 11073
rect 32953 11064 32965 11067
rect 32456 11036 32965 11064
rect 32456 11024 32462 11036
rect 32953 11033 32965 11036
rect 32999 11033 33011 11067
rect 32953 11027 33011 11033
rect 34701 11067 34759 11073
rect 34701 11033 34713 11067
rect 34747 11064 34759 11067
rect 36354 11064 36360 11076
rect 34747 11036 35940 11064
rect 36315 11036 36360 11064
rect 34747 11033 34759 11036
rect 34701 11027 34759 11033
rect 35912 11008 35940 11036
rect 36354 11024 36360 11036
rect 36412 11024 36418 11076
rect 30009 10999 30067 11005
rect 30009 10996 30021 10999
rect 29420 10968 30021 10996
rect 29420 10956 29426 10968
rect 30009 10965 30021 10968
rect 30055 10965 30067 10999
rect 33870 10996 33876 11008
rect 33831 10968 33876 10996
rect 30009 10959 30067 10965
rect 33870 10956 33876 10968
rect 33928 10956 33934 11008
rect 35894 10956 35900 11008
rect 35952 10956 35958 11008
rect 36817 10999 36875 11005
rect 36817 10965 36829 10999
rect 36863 10996 36875 10999
rect 36906 10996 36912 11008
rect 36863 10968 36912 10996
rect 36863 10965 36875 10968
rect 36817 10959 36875 10965
rect 36906 10956 36912 10968
rect 36964 10956 36970 11008
rect 1104 10906 38824 10928
rect 1104 10854 7648 10906
rect 7700 10854 7712 10906
rect 7764 10854 7776 10906
rect 7828 10854 7840 10906
rect 7892 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 34315 10906
rect 34367 10854 34379 10906
rect 34431 10854 34443 10906
rect 34495 10854 34507 10906
rect 34559 10854 38824 10906
rect 1104 10832 38824 10854
rect 2498 10792 2504 10804
rect 2459 10764 2504 10792
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 3602 10752 3608 10804
rect 3660 10792 3666 10804
rect 4065 10795 4123 10801
rect 4065 10792 4077 10795
rect 3660 10764 4077 10792
rect 3660 10752 3666 10764
rect 4065 10761 4077 10764
rect 4111 10761 4123 10795
rect 5718 10792 5724 10804
rect 5679 10764 5724 10792
rect 4065 10755 4123 10761
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 8757 10795 8815 10801
rect 8757 10761 8769 10795
rect 8803 10792 8815 10795
rect 9214 10792 9220 10804
rect 8803 10764 9220 10792
rect 8803 10761 8815 10764
rect 8757 10755 8815 10761
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 10318 10752 10324 10804
rect 10376 10792 10382 10804
rect 10597 10795 10655 10801
rect 10597 10792 10609 10795
rect 10376 10764 10609 10792
rect 10376 10752 10382 10764
rect 10597 10761 10609 10764
rect 10643 10792 10655 10795
rect 11241 10795 11299 10801
rect 11241 10792 11253 10795
rect 10643 10764 11253 10792
rect 10643 10761 10655 10764
rect 10597 10755 10655 10761
rect 11241 10761 11253 10764
rect 11287 10792 11299 10795
rect 11885 10795 11943 10801
rect 11885 10792 11897 10795
rect 11287 10764 11897 10792
rect 11287 10761 11299 10764
rect 11241 10755 11299 10761
rect 11885 10761 11897 10764
rect 11931 10792 11943 10795
rect 12342 10792 12348 10804
rect 11931 10764 12348 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 12526 10792 12532 10804
rect 12487 10764 12532 10792
rect 12526 10752 12532 10764
rect 12584 10752 12590 10804
rect 16117 10795 16175 10801
rect 16117 10761 16129 10795
rect 16163 10792 16175 10795
rect 16390 10792 16396 10804
rect 16163 10764 16396 10792
rect 16163 10761 16175 10764
rect 16117 10755 16175 10761
rect 16390 10752 16396 10764
rect 16448 10752 16454 10804
rect 16482 10752 16488 10804
rect 16540 10792 16546 10804
rect 17129 10795 17187 10801
rect 17129 10792 17141 10795
rect 16540 10764 17141 10792
rect 16540 10752 16546 10764
rect 17129 10761 17141 10764
rect 17175 10761 17187 10795
rect 17129 10755 17187 10761
rect 17862 10752 17868 10804
rect 17920 10792 17926 10804
rect 18233 10795 18291 10801
rect 18233 10792 18245 10795
rect 17920 10764 18245 10792
rect 17920 10752 17926 10764
rect 18233 10761 18245 10764
rect 18279 10761 18291 10795
rect 18690 10792 18696 10804
rect 18651 10764 18696 10792
rect 18233 10755 18291 10761
rect 18690 10752 18696 10764
rect 18748 10752 18754 10804
rect 21726 10752 21732 10804
rect 21784 10792 21790 10804
rect 21821 10795 21879 10801
rect 21821 10792 21833 10795
rect 21784 10764 21833 10792
rect 21784 10752 21790 10764
rect 21821 10761 21833 10764
rect 21867 10761 21879 10795
rect 21821 10755 21879 10761
rect 25958 10752 25964 10804
rect 26016 10792 26022 10804
rect 26142 10792 26148 10804
rect 26016 10764 26148 10792
rect 26016 10752 26022 10764
rect 26142 10752 26148 10764
rect 26200 10792 26206 10804
rect 26605 10795 26663 10801
rect 26605 10792 26617 10795
rect 26200 10764 26617 10792
rect 26200 10752 26206 10764
rect 26605 10761 26617 10764
rect 26651 10761 26663 10795
rect 30650 10792 30656 10804
rect 30611 10764 30656 10792
rect 26605 10755 26663 10761
rect 30650 10752 30656 10764
rect 30708 10752 30714 10804
rect 31665 10795 31723 10801
rect 31665 10761 31677 10795
rect 31711 10792 31723 10795
rect 33318 10792 33324 10804
rect 31711 10764 33324 10792
rect 31711 10761 31723 10764
rect 31665 10755 31723 10761
rect 33318 10752 33324 10764
rect 33376 10752 33382 10804
rect 34701 10795 34759 10801
rect 34701 10761 34713 10795
rect 34747 10792 34759 10795
rect 34790 10792 34796 10804
rect 34747 10764 34796 10792
rect 34747 10761 34759 10764
rect 34701 10755 34759 10761
rect 34790 10752 34796 10764
rect 34848 10792 34854 10804
rect 36538 10792 36544 10804
rect 34848 10764 35112 10792
rect 36499 10764 36544 10792
rect 34848 10752 34854 10764
rect 6914 10724 6920 10736
rect 6875 10696 6920 10724
rect 6914 10684 6920 10696
rect 6972 10684 6978 10736
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10616 1458 10668
rect 1949 10659 2007 10665
rect 1949 10625 1961 10659
rect 1995 10656 2007 10659
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 1995 10628 2881 10656
rect 1995 10625 2007 10628
rect 1949 10619 2007 10625
rect 2869 10625 2881 10628
rect 2915 10656 2927 10659
rect 3786 10656 3792 10668
rect 2915 10628 3792 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 3786 10616 3792 10628
rect 3844 10616 3850 10668
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 4525 10659 4583 10665
rect 4525 10656 4537 10659
rect 4396 10628 4537 10656
rect 4396 10616 4402 10628
rect 4525 10625 4537 10628
rect 4571 10656 4583 10659
rect 6178 10656 6184 10668
rect 4571 10628 6184 10656
rect 4571 10625 4583 10628
rect 4525 10619 4583 10625
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 12158 10616 12164 10668
rect 12216 10656 12222 10668
rect 13817 10659 13875 10665
rect 13817 10656 13829 10659
rect 12216 10628 13829 10656
rect 12216 10616 12222 10628
rect 13817 10625 13829 10628
rect 13863 10656 13875 10659
rect 14001 10659 14059 10665
rect 14001 10656 14013 10659
rect 13863 10628 14013 10656
rect 13863 10625 13875 10628
rect 13817 10619 13875 10625
rect 14001 10625 14013 10628
rect 14047 10625 14059 10659
rect 14001 10619 14059 10625
rect 4617 10591 4675 10597
rect 4617 10588 4629 10591
rect 3160 10560 4629 10588
rect 3160 10532 3188 10560
rect 4617 10557 4629 10560
rect 4663 10588 4675 10591
rect 4985 10591 5043 10597
rect 4985 10588 4997 10591
rect 4663 10560 4997 10588
rect 4663 10557 4675 10560
rect 4617 10551 4675 10557
rect 4985 10557 4997 10560
rect 5031 10557 5043 10591
rect 5537 10591 5595 10597
rect 5537 10588 5549 10591
rect 4985 10551 5043 10557
rect 5460 10560 5549 10588
rect 2317 10523 2375 10529
rect 2317 10489 2329 10523
rect 2363 10520 2375 10523
rect 2958 10520 2964 10532
rect 2363 10492 2964 10520
rect 2363 10489 2375 10492
rect 2317 10483 2375 10489
rect 2958 10480 2964 10492
rect 3016 10480 3022 10532
rect 3053 10523 3111 10529
rect 3053 10489 3065 10523
rect 3099 10520 3111 10523
rect 3142 10520 3148 10532
rect 3099 10492 3148 10520
rect 3099 10489 3111 10492
rect 3053 10483 3111 10489
rect 3142 10480 3148 10492
rect 3200 10480 3206 10532
rect 4525 10523 4583 10529
rect 4525 10520 4537 10523
rect 3436 10492 4537 10520
rect 3234 10412 3240 10464
rect 3292 10452 3298 10464
rect 3436 10461 3464 10492
rect 4525 10489 4537 10492
rect 4571 10489 4583 10523
rect 4525 10483 4583 10489
rect 5460 10464 5488 10560
rect 5537 10557 5549 10560
rect 5583 10557 5595 10591
rect 7469 10591 7527 10597
rect 7469 10588 7481 10591
rect 5537 10551 5595 10557
rect 6564 10560 7481 10588
rect 3421 10455 3479 10461
rect 3421 10452 3433 10455
rect 3292 10424 3433 10452
rect 3292 10412 3298 10424
rect 3421 10421 3433 10424
rect 3467 10421 3479 10455
rect 3421 10415 3479 10421
rect 3602 10412 3608 10464
rect 3660 10452 3666 10464
rect 3789 10455 3847 10461
rect 3789 10452 3801 10455
rect 3660 10424 3801 10452
rect 3660 10412 3666 10424
rect 3789 10421 3801 10424
rect 3835 10452 3847 10455
rect 4706 10452 4712 10464
rect 3835 10424 4712 10452
rect 3835 10421 3847 10424
rect 3789 10415 3847 10421
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 5442 10452 5448 10464
rect 5403 10424 5448 10452
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 6178 10452 6184 10464
rect 6139 10424 6184 10452
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 6362 10412 6368 10464
rect 6420 10452 6426 10464
rect 6564 10461 6592 10560
rect 7469 10557 7481 10560
rect 7515 10557 7527 10591
rect 7469 10551 7527 10557
rect 8941 10591 8999 10597
rect 8941 10557 8953 10591
rect 8987 10588 8999 10591
rect 9217 10591 9275 10597
rect 9217 10588 9229 10591
rect 8987 10560 9229 10588
rect 8987 10557 8999 10560
rect 8941 10551 8999 10557
rect 9217 10557 9229 10560
rect 9263 10557 9275 10591
rect 10042 10588 10048 10600
rect 9217 10551 9275 10557
rect 9416 10560 10048 10588
rect 7190 10520 7196 10532
rect 7151 10492 7196 10520
rect 7190 10480 7196 10492
rect 7248 10480 7254 10532
rect 8389 10523 8447 10529
rect 8389 10489 8401 10523
rect 8435 10520 8447 10523
rect 9416 10520 9444 10560
rect 10042 10548 10048 10560
rect 10100 10548 10106 10600
rect 12802 10588 12808 10600
rect 12763 10560 12808 10588
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 14016 10588 14044 10619
rect 16298 10616 16304 10668
rect 16356 10656 16362 10668
rect 16393 10659 16451 10665
rect 16393 10656 16405 10659
rect 16356 10628 16405 10656
rect 16356 10616 16362 10628
rect 16393 10625 16405 10628
rect 16439 10625 16451 10659
rect 16393 10619 16451 10625
rect 16669 10659 16727 10665
rect 16669 10625 16681 10659
rect 16715 10656 16727 10659
rect 17494 10656 17500 10668
rect 16715 10628 17500 10656
rect 16715 10625 16727 10628
rect 16669 10619 16727 10625
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 18708 10656 18736 10752
rect 23753 10727 23811 10733
rect 23753 10724 23765 10727
rect 22296 10696 23765 10724
rect 18708 10628 19380 10656
rect 14734 10588 14740 10600
rect 14016 10560 14740 10588
rect 14734 10548 14740 10560
rect 14792 10548 14798 10600
rect 19245 10591 19303 10597
rect 19245 10588 19257 10591
rect 19076 10560 19257 10588
rect 9490 10529 9496 10532
rect 8435 10492 9444 10520
rect 8435 10489 8447 10492
rect 8389 10483 8447 10489
rect 9484 10483 9496 10529
rect 9548 10520 9554 10532
rect 13078 10520 13084 10532
rect 9548 10492 9584 10520
rect 13039 10492 13084 10520
rect 9490 10480 9496 10483
rect 9548 10480 9554 10492
rect 13078 10480 13084 10492
rect 13136 10520 13142 10532
rect 13449 10523 13507 10529
rect 13449 10520 13461 10523
rect 13136 10492 13461 10520
rect 13136 10480 13142 10492
rect 13449 10489 13461 10492
rect 13495 10520 13507 10523
rect 13630 10520 13636 10532
rect 13495 10492 13636 10520
rect 13495 10489 13507 10492
rect 13449 10483 13507 10489
rect 13630 10480 13636 10492
rect 13688 10520 13694 10532
rect 14246 10523 14304 10529
rect 14246 10520 14258 10523
rect 13688 10492 14258 10520
rect 13688 10480 13694 10492
rect 14246 10489 14258 10492
rect 14292 10489 14304 10523
rect 14246 10483 14304 10489
rect 6549 10455 6607 10461
rect 6549 10452 6561 10455
rect 6420 10424 6561 10452
rect 6420 10412 6426 10424
rect 6549 10421 6561 10424
rect 6595 10421 6607 10455
rect 6549 10415 6607 10421
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 7377 10455 7435 10461
rect 7377 10452 7389 10455
rect 7064 10424 7389 10452
rect 7064 10412 7070 10424
rect 7377 10421 7389 10424
rect 7423 10421 7435 10455
rect 7377 10415 7435 10421
rect 8110 10412 8116 10464
rect 8168 10452 8174 10464
rect 8941 10455 8999 10461
rect 8941 10452 8953 10455
rect 8168 10424 8953 10452
rect 8168 10412 8174 10424
rect 8941 10421 8953 10424
rect 8987 10452 8999 10455
rect 9033 10455 9091 10461
rect 9033 10452 9045 10455
rect 8987 10424 9045 10452
rect 8987 10421 8999 10424
rect 8941 10415 8999 10421
rect 9033 10421 9045 10424
rect 9079 10421 9091 10455
rect 12158 10452 12164 10464
rect 12119 10424 12164 10452
rect 9033 10415 9091 10421
rect 12158 10412 12164 10424
rect 12216 10412 12222 10464
rect 12986 10452 12992 10464
rect 12947 10424 12992 10452
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 15378 10452 15384 10464
rect 15339 10424 15384 10452
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 17310 10412 17316 10464
rect 17368 10452 17374 10464
rect 19076 10461 19104 10560
rect 19245 10557 19257 10560
rect 19291 10557 19303 10591
rect 19352 10588 19380 10628
rect 22094 10616 22100 10668
rect 22152 10656 22158 10668
rect 22296 10665 22324 10696
rect 23753 10693 23765 10696
rect 23799 10693 23811 10727
rect 23753 10687 23811 10693
rect 26510 10684 26516 10736
rect 26568 10724 26574 10736
rect 27154 10724 27160 10736
rect 26568 10696 27160 10724
rect 26568 10684 26574 10696
rect 27154 10684 27160 10696
rect 27212 10684 27218 10736
rect 32306 10724 32312 10736
rect 32267 10696 32312 10724
rect 32306 10684 32312 10696
rect 32364 10684 32370 10736
rect 34977 10727 35035 10733
rect 34977 10693 34989 10727
rect 35023 10693 35035 10727
rect 34977 10687 35035 10693
rect 22281 10659 22339 10665
rect 22281 10656 22293 10659
rect 22152 10628 22293 10656
rect 22152 10616 22158 10628
rect 22281 10625 22293 10628
rect 22327 10625 22339 10659
rect 22281 10619 22339 10625
rect 22370 10616 22376 10668
rect 22428 10656 22434 10668
rect 22428 10628 22473 10656
rect 22428 10616 22434 10628
rect 22646 10616 22652 10668
rect 22704 10656 22710 10668
rect 22833 10659 22891 10665
rect 22833 10656 22845 10659
rect 22704 10628 22845 10656
rect 22704 10616 22710 10628
rect 22833 10625 22845 10628
rect 22879 10656 22891 10659
rect 23842 10656 23848 10668
rect 22879 10628 23848 10656
rect 22879 10625 22891 10628
rect 22833 10619 22891 10625
rect 23842 10616 23848 10628
rect 23900 10656 23906 10668
rect 24305 10659 24363 10665
rect 24305 10656 24317 10659
rect 23900 10628 24317 10656
rect 23900 10616 23906 10628
rect 24305 10625 24317 10628
rect 24351 10625 24363 10659
rect 24305 10619 24363 10625
rect 33134 10616 33140 10668
rect 33192 10656 33198 10668
rect 33873 10659 33931 10665
rect 33873 10656 33885 10659
rect 33192 10628 33885 10656
rect 33192 10616 33198 10628
rect 33873 10625 33885 10628
rect 33919 10656 33931 10659
rect 34698 10656 34704 10668
rect 33919 10628 34704 10656
rect 33919 10625 33931 10628
rect 33873 10619 33931 10625
rect 34698 10616 34704 10628
rect 34756 10616 34762 10668
rect 19501 10591 19559 10597
rect 19501 10588 19513 10591
rect 19352 10560 19513 10588
rect 19245 10551 19303 10557
rect 19501 10557 19513 10560
rect 19547 10557 19559 10591
rect 23290 10588 23296 10600
rect 19501 10551 19559 10557
rect 22296 10560 23296 10588
rect 22296 10532 22324 10560
rect 23290 10548 23296 10560
rect 23348 10548 23354 10600
rect 23477 10591 23535 10597
rect 23477 10557 23489 10591
rect 23523 10588 23535 10591
rect 23658 10588 23664 10600
rect 23523 10560 23664 10588
rect 23523 10557 23535 10560
rect 23477 10551 23535 10557
rect 23658 10548 23664 10560
rect 23716 10548 23722 10600
rect 23750 10548 23756 10600
rect 23808 10588 23814 10600
rect 24673 10591 24731 10597
rect 24673 10588 24685 10591
rect 23808 10560 24685 10588
rect 23808 10548 23814 10560
rect 24673 10557 24685 10560
rect 24719 10588 24731 10591
rect 25041 10591 25099 10597
rect 25041 10588 25053 10591
rect 24719 10560 25053 10588
rect 24719 10557 24731 10560
rect 24673 10551 24731 10557
rect 25041 10557 25053 10560
rect 25087 10588 25099 10591
rect 25130 10588 25136 10600
rect 25087 10560 25136 10588
rect 25087 10557 25099 10560
rect 25041 10551 25099 10557
rect 25130 10548 25136 10560
rect 25188 10588 25194 10600
rect 25225 10591 25283 10597
rect 25225 10588 25237 10591
rect 25188 10560 25237 10588
rect 25188 10548 25194 10560
rect 25225 10557 25237 10560
rect 25271 10588 25283 10591
rect 25314 10588 25320 10600
rect 25271 10560 25320 10588
rect 25271 10557 25283 10560
rect 25225 10551 25283 10557
rect 25314 10548 25320 10560
rect 25372 10548 25378 10600
rect 29273 10591 29331 10597
rect 29273 10557 29285 10591
rect 29319 10588 29331 10591
rect 29362 10588 29368 10600
rect 29319 10560 29368 10588
rect 29319 10557 29331 10560
rect 29273 10551 29331 10557
rect 29362 10548 29368 10560
rect 29420 10548 29426 10600
rect 32122 10588 32128 10600
rect 32083 10560 32128 10588
rect 32122 10548 32128 10560
rect 32180 10588 32186 10600
rect 32677 10591 32735 10597
rect 32677 10588 32689 10591
rect 32180 10560 32689 10588
rect 32180 10548 32186 10560
rect 32677 10557 32689 10560
rect 32723 10557 32735 10591
rect 32677 10551 32735 10557
rect 22278 10520 22284 10532
rect 22191 10492 22284 10520
rect 22278 10480 22284 10492
rect 22336 10480 22342 10532
rect 23676 10520 23704 10548
rect 24029 10523 24087 10529
rect 24029 10520 24041 10523
rect 23676 10492 24041 10520
rect 24029 10489 24041 10492
rect 24075 10489 24087 10523
rect 24029 10483 24087 10489
rect 25492 10523 25550 10529
rect 25492 10489 25504 10523
rect 25538 10520 25550 10523
rect 25682 10520 25688 10532
rect 25538 10492 25688 10520
rect 25538 10489 25550 10492
rect 25492 10483 25550 10489
rect 25682 10480 25688 10492
rect 25740 10480 25746 10532
rect 29086 10480 29092 10532
rect 29144 10520 29150 10532
rect 29518 10523 29576 10529
rect 29518 10520 29530 10523
rect 29144 10492 29530 10520
rect 29144 10480 29150 10492
rect 29518 10489 29530 10492
rect 29564 10489 29576 10523
rect 29518 10483 29576 10489
rect 31662 10480 31668 10532
rect 31720 10520 31726 10532
rect 33045 10523 33103 10529
rect 33045 10520 33057 10523
rect 31720 10492 33057 10520
rect 31720 10480 31726 10492
rect 33045 10489 33057 10492
rect 33091 10520 33103 10523
rect 33594 10520 33600 10532
rect 33091 10492 33600 10520
rect 33091 10489 33103 10492
rect 33045 10483 33103 10489
rect 33594 10480 33600 10492
rect 33652 10480 33658 10532
rect 34716 10520 34744 10616
rect 34992 10588 35020 10687
rect 35084 10656 35112 10764
rect 36538 10752 36544 10764
rect 36596 10752 36602 10804
rect 35345 10659 35403 10665
rect 35345 10656 35357 10659
rect 35084 10628 35357 10656
rect 35345 10625 35357 10628
rect 35391 10625 35403 10659
rect 35345 10619 35403 10625
rect 35894 10616 35900 10668
rect 35952 10656 35958 10668
rect 36909 10659 36967 10665
rect 36909 10656 36921 10659
rect 35952 10628 36921 10656
rect 35952 10616 35958 10628
rect 36909 10625 36921 10628
rect 36955 10656 36967 10659
rect 37090 10656 37096 10668
rect 36955 10628 37096 10656
rect 36955 10625 36967 10628
rect 36909 10619 36967 10625
rect 37090 10616 37096 10628
rect 37148 10616 37154 10668
rect 37461 10591 37519 10597
rect 37461 10588 37473 10591
rect 34992 10560 37473 10588
rect 35342 10520 35348 10532
rect 34716 10492 35348 10520
rect 35342 10480 35348 10492
rect 35400 10520 35406 10532
rect 37016 10529 37044 10560
rect 37461 10557 37473 10560
rect 37507 10557 37519 10591
rect 37461 10551 37519 10557
rect 35529 10523 35587 10529
rect 35529 10520 35541 10523
rect 35400 10492 35541 10520
rect 35400 10480 35406 10492
rect 35529 10489 35541 10492
rect 35575 10489 35587 10523
rect 35529 10483 35587 10489
rect 37001 10523 37059 10529
rect 37001 10489 37013 10523
rect 37047 10489 37059 10523
rect 37001 10483 37059 10489
rect 37093 10523 37151 10529
rect 37093 10489 37105 10523
rect 37139 10489 37151 10523
rect 37093 10483 37151 10489
rect 17589 10455 17647 10461
rect 17589 10452 17601 10455
rect 17368 10424 17601 10452
rect 17368 10412 17374 10424
rect 17589 10421 17601 10424
rect 17635 10452 17647 10455
rect 19061 10455 19119 10461
rect 19061 10452 19073 10455
rect 17635 10424 19073 10452
rect 17635 10421 17647 10424
rect 17589 10415 17647 10421
rect 19061 10421 19073 10424
rect 19107 10421 19119 10455
rect 19061 10415 19119 10421
rect 19518 10412 19524 10464
rect 19576 10452 19582 10464
rect 20625 10455 20683 10461
rect 20625 10452 20637 10455
rect 19576 10424 20637 10452
rect 19576 10412 19582 10424
rect 20625 10421 20637 10424
rect 20671 10452 20683 10455
rect 21174 10452 21180 10464
rect 20671 10424 21180 10452
rect 20671 10421 20683 10424
rect 20625 10415 20683 10421
rect 21174 10412 21180 10424
rect 21232 10412 21238 10464
rect 21266 10412 21272 10464
rect 21324 10452 21330 10464
rect 21361 10455 21419 10461
rect 21361 10452 21373 10455
rect 21324 10424 21373 10452
rect 21324 10412 21330 10424
rect 21361 10421 21373 10424
rect 21407 10421 21419 10455
rect 21361 10415 21419 10421
rect 23474 10412 23480 10464
rect 23532 10452 23538 10464
rect 24213 10455 24271 10461
rect 24213 10452 24225 10455
rect 23532 10424 24225 10452
rect 23532 10412 23538 10424
rect 24213 10421 24225 10424
rect 24259 10421 24271 10455
rect 28350 10452 28356 10464
rect 28311 10424 28356 10452
rect 24213 10415 24271 10421
rect 28350 10412 28356 10424
rect 28408 10412 28414 10464
rect 28626 10452 28632 10464
rect 28587 10424 28632 10452
rect 28626 10412 28632 10424
rect 28684 10412 28690 10464
rect 28997 10455 29055 10461
rect 28997 10421 29009 10455
rect 29043 10452 29055 10455
rect 29178 10452 29184 10464
rect 29043 10424 29184 10452
rect 29043 10421 29055 10424
rect 28997 10415 29055 10421
rect 29178 10412 29184 10424
rect 29236 10412 29242 10464
rect 30374 10412 30380 10464
rect 30432 10452 30438 10464
rect 30926 10452 30932 10464
rect 30432 10424 30932 10452
rect 30432 10412 30438 10424
rect 30926 10412 30932 10424
rect 30984 10452 30990 10464
rect 31205 10455 31263 10461
rect 31205 10452 31217 10455
rect 30984 10424 31217 10452
rect 30984 10412 30990 10424
rect 31205 10421 31217 10424
rect 31251 10421 31263 10455
rect 31205 10415 31263 10421
rect 32033 10455 32091 10461
rect 32033 10421 32045 10455
rect 32079 10452 32091 10455
rect 32950 10452 32956 10464
rect 32079 10424 32956 10452
rect 32079 10421 32091 10424
rect 32033 10415 32091 10421
rect 32950 10412 32956 10424
rect 33008 10412 33014 10464
rect 33318 10412 33324 10464
rect 33376 10452 33382 10464
rect 33781 10455 33839 10461
rect 33781 10452 33793 10455
rect 33376 10424 33793 10452
rect 33376 10412 33382 10424
rect 33781 10421 33793 10424
rect 33827 10452 33839 10455
rect 33870 10452 33876 10464
rect 33827 10424 33876 10452
rect 33827 10421 33839 10424
rect 33781 10415 33839 10421
rect 33870 10412 33876 10424
rect 33928 10412 33934 10464
rect 34330 10452 34336 10464
rect 34291 10424 34336 10452
rect 34330 10412 34336 10424
rect 34388 10412 34394 10464
rect 35434 10452 35440 10464
rect 35395 10424 35440 10452
rect 35434 10412 35440 10424
rect 35492 10412 35498 10464
rect 36170 10452 36176 10464
rect 36131 10424 36176 10452
rect 36170 10412 36176 10424
rect 36228 10412 36234 10464
rect 36906 10412 36912 10464
rect 36964 10452 36970 10464
rect 37108 10452 37136 10483
rect 36964 10424 37136 10452
rect 36964 10412 36970 10424
rect 1104 10362 38824 10384
rect 1104 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 27648 10362
rect 27700 10310 27712 10362
rect 27764 10310 27776 10362
rect 27828 10310 27840 10362
rect 27892 10310 38824 10362
rect 1104 10288 38824 10310
rect 2498 10248 2504 10260
rect 2459 10220 2504 10248
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 4338 10248 4344 10260
rect 4299 10220 4344 10248
rect 4338 10208 4344 10220
rect 4396 10208 4402 10260
rect 5902 10248 5908 10260
rect 5863 10220 5908 10248
rect 5902 10208 5908 10220
rect 5960 10208 5966 10260
rect 9674 10208 9680 10260
rect 9732 10208 9738 10260
rect 10226 10248 10232 10260
rect 10187 10220 10232 10248
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 11330 10208 11336 10260
rect 11388 10248 11394 10260
rect 12069 10251 12127 10257
rect 12069 10248 12081 10251
rect 11388 10220 12081 10248
rect 11388 10208 11394 10220
rect 12069 10217 12081 10220
rect 12115 10248 12127 10251
rect 12434 10248 12440 10260
rect 12115 10220 12440 10248
rect 12115 10217 12127 10220
rect 12069 10211 12127 10217
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 12986 10248 12992 10260
rect 12947 10220 12992 10248
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 16114 10248 16120 10260
rect 16075 10220 16120 10248
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 17773 10251 17831 10257
rect 17773 10217 17785 10251
rect 17819 10248 17831 10251
rect 17862 10248 17868 10260
rect 17819 10220 17868 10248
rect 17819 10217 17831 10220
rect 17773 10211 17831 10217
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 20717 10251 20775 10257
rect 20717 10217 20729 10251
rect 20763 10248 20775 10251
rect 22094 10248 22100 10260
rect 20763 10220 22100 10248
rect 20763 10217 20775 10220
rect 20717 10211 20775 10217
rect 22094 10208 22100 10220
rect 22152 10208 22158 10260
rect 22646 10248 22652 10260
rect 22607 10220 22652 10248
rect 22646 10208 22652 10220
rect 22704 10208 22710 10260
rect 24118 10248 24124 10260
rect 24079 10220 24124 10248
rect 24118 10208 24124 10220
rect 24176 10208 24182 10260
rect 25222 10248 25228 10260
rect 25183 10220 25228 10248
rect 25222 10208 25228 10220
rect 25280 10248 25286 10260
rect 26053 10251 26111 10257
rect 26053 10248 26065 10251
rect 25280 10220 26065 10248
rect 25280 10208 25286 10220
rect 26053 10217 26065 10220
rect 26099 10217 26111 10251
rect 26970 10248 26976 10260
rect 26931 10220 26976 10248
rect 26053 10211 26111 10217
rect 26970 10208 26976 10220
rect 27028 10208 27034 10260
rect 29825 10251 29883 10257
rect 29825 10217 29837 10251
rect 29871 10248 29883 10251
rect 31754 10248 31760 10260
rect 29871 10220 31760 10248
rect 29871 10217 29883 10220
rect 29825 10211 29883 10217
rect 31754 10208 31760 10220
rect 31812 10208 31818 10260
rect 36541 10251 36599 10257
rect 36541 10217 36553 10251
rect 36587 10248 36599 10251
rect 36906 10248 36912 10260
rect 36587 10220 36912 10248
rect 36587 10217 36599 10220
rect 36541 10211 36599 10217
rect 36906 10208 36912 10220
rect 36964 10208 36970 10260
rect 37090 10248 37096 10260
rect 37051 10220 37096 10248
rect 37090 10208 37096 10220
rect 37148 10208 37154 10260
rect 1857 10183 1915 10189
rect 1857 10149 1869 10183
rect 1903 10180 1915 10183
rect 2593 10183 2651 10189
rect 2593 10180 2605 10183
rect 1903 10152 2605 10180
rect 1903 10149 1915 10152
rect 1857 10143 1915 10149
rect 2593 10149 2605 10152
rect 2639 10180 2651 10183
rect 2682 10180 2688 10192
rect 2639 10152 2688 10180
rect 2639 10149 2651 10152
rect 2593 10143 2651 10149
rect 2682 10140 2688 10152
rect 2740 10180 2746 10192
rect 3421 10183 3479 10189
rect 3421 10180 3433 10183
rect 2740 10152 3433 10180
rect 2740 10140 2746 10152
rect 3421 10149 3433 10152
rect 3467 10180 3479 10183
rect 4522 10180 4528 10192
rect 3467 10152 4528 10180
rect 3467 10149 3479 10152
rect 3421 10143 3479 10149
rect 4522 10140 4528 10152
rect 4580 10180 4586 10192
rect 4770 10183 4828 10189
rect 4770 10180 4782 10183
rect 4580 10152 4782 10180
rect 4580 10140 4586 10152
rect 4770 10149 4782 10152
rect 4816 10149 4828 10183
rect 5920 10180 5948 10208
rect 7254 10183 7312 10189
rect 7254 10180 7266 10183
rect 5920 10152 7266 10180
rect 4770 10143 4828 10149
rect 7254 10149 7266 10152
rect 7300 10149 7312 10183
rect 7254 10143 7312 10149
rect 7009 10115 7067 10121
rect 7009 10081 7021 10115
rect 7055 10112 7067 10115
rect 7098 10112 7104 10124
rect 7055 10084 7104 10112
rect 7055 10081 7067 10084
rect 7009 10075 7067 10081
rect 7098 10072 7104 10084
rect 7156 10072 7162 10124
rect 9692 10112 9720 10208
rect 12621 10183 12679 10189
rect 12621 10149 12633 10183
rect 12667 10180 12679 10183
rect 13078 10180 13084 10192
rect 12667 10152 13084 10180
rect 12667 10149 12679 10152
rect 12621 10143 12679 10149
rect 13078 10140 13084 10152
rect 13136 10140 13142 10192
rect 13906 10140 13912 10192
rect 13964 10180 13970 10192
rect 14185 10183 14243 10189
rect 14185 10180 14197 10183
rect 13964 10152 14197 10180
rect 13964 10140 13970 10152
rect 14185 10149 14197 10152
rect 14231 10149 14243 10183
rect 14185 10143 14243 10149
rect 19334 10140 19340 10192
rect 19392 10180 19398 10192
rect 19797 10183 19855 10189
rect 19797 10180 19809 10183
rect 19392 10152 19809 10180
rect 19392 10140 19398 10152
rect 19797 10149 19809 10152
rect 19843 10149 19855 10183
rect 19797 10143 19855 10149
rect 21266 10140 21272 10192
rect 21324 10180 21330 10192
rect 21324 10152 21956 10180
rect 21324 10140 21330 10152
rect 21928 10124 21956 10152
rect 22002 10140 22008 10192
rect 22060 10180 22066 10192
rect 22186 10180 22192 10192
rect 22060 10152 22192 10180
rect 22060 10140 22066 10152
rect 22186 10140 22192 10152
rect 22244 10140 22250 10192
rect 25682 10180 25688 10192
rect 25643 10152 25688 10180
rect 25682 10140 25688 10152
rect 25740 10140 25746 10192
rect 27522 10140 27528 10192
rect 27580 10180 27586 10192
rect 32950 10189 32956 10192
rect 28261 10183 28319 10189
rect 28261 10180 28273 10183
rect 27580 10152 28273 10180
rect 27580 10140 27586 10152
rect 28261 10149 28273 10152
rect 28307 10180 28319 10183
rect 29347 10183 29405 10189
rect 29347 10180 29359 10183
rect 28307 10152 29359 10180
rect 28307 10149 28319 10152
rect 28261 10143 28319 10149
rect 29347 10149 29359 10152
rect 29393 10149 29405 10183
rect 29347 10143 29405 10149
rect 32585 10183 32643 10189
rect 32585 10149 32597 10183
rect 32631 10180 32643 10183
rect 32944 10180 32956 10189
rect 32631 10152 32956 10180
rect 32631 10149 32643 10152
rect 32585 10143 32643 10149
rect 32944 10143 32956 10152
rect 32950 10140 32956 10143
rect 33008 10140 33014 10192
rect 33042 10140 33048 10192
rect 33100 10140 33106 10192
rect 35342 10140 35348 10192
rect 35400 10189 35406 10192
rect 35400 10183 35464 10189
rect 35400 10149 35418 10183
rect 35452 10180 35464 10183
rect 35526 10180 35532 10192
rect 35452 10152 35532 10180
rect 35452 10149 35464 10152
rect 35400 10143 35464 10149
rect 35400 10140 35406 10143
rect 35526 10140 35532 10152
rect 35584 10140 35590 10192
rect 9950 10112 9956 10124
rect 9692 10084 9956 10112
rect 9950 10072 9956 10084
rect 10008 10112 10014 10124
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 10008 10084 10057 10112
rect 10008 10072 10014 10084
rect 10045 10081 10057 10084
rect 10091 10081 10103 10115
rect 10045 10075 10103 10081
rect 11425 10115 11483 10121
rect 11425 10081 11437 10115
rect 11471 10112 11483 10115
rect 11471 10084 12204 10112
rect 11471 10081 11483 10084
rect 11425 10075 11483 10081
rect 2406 10044 2412 10056
rect 2367 10016 2412 10044
rect 2406 10004 2412 10016
rect 2464 10004 2470 10056
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10044 9367 10047
rect 9490 10044 9496 10056
rect 9355 10016 9496 10044
rect 9355 10013 9367 10016
rect 9309 10007 9367 10013
rect 2038 9976 2044 9988
rect 1999 9948 2044 9976
rect 2038 9936 2044 9948
rect 2096 9936 2102 9988
rect 3053 9911 3111 9917
rect 3053 9877 3065 9911
rect 3099 9908 3111 9911
rect 3142 9908 3148 9920
rect 3099 9880 3148 9908
rect 3099 9877 3111 9880
rect 3053 9871 3111 9877
rect 3142 9868 3148 9880
rect 3200 9868 3206 9920
rect 3878 9908 3884 9920
rect 3839 9880 3884 9908
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 4540 9908 4568 10007
rect 9490 10004 9496 10016
rect 9548 10044 9554 10056
rect 10321 10047 10379 10053
rect 10321 10044 10333 10047
rect 9548 10016 10333 10044
rect 9548 10004 9554 10016
rect 10321 10013 10333 10016
rect 10367 10013 10379 10047
rect 12066 10044 12072 10056
rect 12027 10016 12072 10044
rect 10321 10007 10379 10013
rect 9769 9979 9827 9985
rect 9769 9945 9781 9979
rect 9815 9976 9827 9979
rect 10042 9976 10048 9988
rect 9815 9948 10048 9976
rect 9815 9945 9827 9948
rect 9769 9939 9827 9945
rect 10042 9936 10048 9948
rect 10100 9936 10106 9988
rect 4706 9908 4712 9920
rect 4540 9880 4712 9908
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 6454 9908 6460 9920
rect 6415 9880 6460 9908
rect 6454 9868 6460 9880
rect 6512 9868 6518 9920
rect 6917 9911 6975 9917
rect 6917 9877 6929 9911
rect 6963 9908 6975 9911
rect 7006 9908 7012 9920
rect 6963 9880 7012 9908
rect 6963 9877 6975 9880
rect 6917 9871 6975 9877
rect 7006 9868 7012 9880
rect 7064 9868 7070 9920
rect 8202 9868 8208 9920
rect 8260 9908 8266 9920
rect 8389 9911 8447 9917
rect 8389 9908 8401 9911
rect 8260 9880 8401 9908
rect 8260 9868 8266 9880
rect 8389 9877 8401 9880
rect 8435 9877 8447 9911
rect 10336 9908 10364 10007
rect 12066 10004 12072 10016
rect 12124 10004 12130 10056
rect 12176 10053 12204 10084
rect 12802 10072 12808 10124
rect 12860 10112 12866 10124
rect 13265 10115 13323 10121
rect 13265 10112 13277 10115
rect 12860 10084 13277 10112
rect 12860 10072 12866 10084
rect 13265 10081 13277 10084
rect 13311 10081 13323 10115
rect 13265 10075 13323 10081
rect 14090 10072 14096 10124
rect 14148 10112 14154 10124
rect 14277 10115 14335 10121
rect 14277 10112 14289 10115
rect 14148 10084 14289 10112
rect 14148 10072 14154 10084
rect 14277 10081 14289 10084
rect 14323 10112 14335 10115
rect 15102 10112 15108 10124
rect 14323 10084 15108 10112
rect 14323 10081 14335 10084
rect 14277 10075 14335 10081
rect 15102 10072 15108 10084
rect 15160 10112 15166 10124
rect 16649 10115 16707 10121
rect 16649 10112 16661 10115
rect 15160 10084 16661 10112
rect 15160 10072 15166 10084
rect 16649 10081 16661 10084
rect 16695 10112 16707 10115
rect 16942 10112 16948 10124
rect 16695 10084 16948 10112
rect 16695 10081 16707 10084
rect 16649 10075 16707 10081
rect 16942 10072 16948 10084
rect 17000 10112 17006 10124
rect 17586 10112 17592 10124
rect 17000 10084 17592 10112
rect 17000 10072 17006 10084
rect 17586 10072 17592 10084
rect 17644 10072 17650 10124
rect 21174 10112 21180 10124
rect 21087 10084 21180 10112
rect 21174 10072 21180 10084
rect 21232 10112 21238 10124
rect 21536 10115 21594 10121
rect 21536 10112 21548 10115
rect 21232 10084 21548 10112
rect 21232 10072 21238 10084
rect 21536 10081 21548 10084
rect 21582 10112 21594 10115
rect 21818 10112 21824 10124
rect 21582 10084 21824 10112
rect 21582 10081 21594 10084
rect 21536 10075 21594 10081
rect 21818 10072 21824 10084
rect 21876 10072 21882 10124
rect 21910 10072 21916 10124
rect 21968 10112 21974 10124
rect 23750 10112 23756 10124
rect 21968 10084 23756 10112
rect 21968 10072 21974 10084
rect 23750 10072 23756 10084
rect 23808 10072 23814 10124
rect 24946 10072 24952 10124
rect 25004 10112 25010 10124
rect 25041 10115 25099 10121
rect 25041 10112 25053 10115
rect 25004 10084 25053 10112
rect 25004 10072 25010 10084
rect 25041 10081 25053 10084
rect 25087 10081 25099 10115
rect 25314 10112 25320 10124
rect 25041 10075 25099 10081
rect 25148 10084 25320 10112
rect 12161 10047 12219 10053
rect 12161 10013 12173 10047
rect 12207 10044 12219 10047
rect 12342 10044 12348 10056
rect 12207 10016 12348 10044
rect 12207 10013 12219 10016
rect 12161 10007 12219 10013
rect 12342 10004 12348 10016
rect 12400 10004 12406 10056
rect 14182 10044 14188 10056
rect 14143 10016 14188 10044
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 15286 10004 15292 10056
rect 15344 10044 15350 10056
rect 16390 10044 16396 10056
rect 15344 10016 16396 10044
rect 15344 10004 15350 10016
rect 16390 10004 16396 10016
rect 16448 10004 16454 10056
rect 19153 10047 19211 10053
rect 19153 10013 19165 10047
rect 19199 10044 19211 10047
rect 19794 10044 19800 10056
rect 19199 10016 19800 10044
rect 19199 10013 19211 10016
rect 19153 10007 19211 10013
rect 19794 10004 19800 10016
rect 19852 10004 19858 10056
rect 19886 10004 19892 10056
rect 19944 10044 19950 10056
rect 19944 10016 21220 10044
rect 19944 10004 19950 10016
rect 11609 9979 11667 9985
rect 11609 9945 11621 9979
rect 11655 9976 11667 9979
rect 12986 9976 12992 9988
rect 11655 9948 12992 9976
rect 11655 9945 11667 9948
rect 11609 9939 11667 9945
rect 12986 9936 12992 9948
rect 13044 9936 13050 9988
rect 13538 9936 13544 9988
rect 13596 9976 13602 9988
rect 13725 9979 13783 9985
rect 13725 9976 13737 9979
rect 13596 9948 13737 9976
rect 13596 9936 13602 9948
rect 13725 9945 13737 9948
rect 13771 9945 13783 9979
rect 13725 9939 13783 9945
rect 19337 9979 19395 9985
rect 19337 9945 19349 9979
rect 19383 9976 19395 9979
rect 20622 9976 20628 9988
rect 19383 9948 20628 9976
rect 19383 9945 19395 9948
rect 19337 9939 19395 9945
rect 20622 9936 20628 9948
rect 20680 9936 20686 9988
rect 10873 9911 10931 9917
rect 10873 9908 10885 9911
rect 10336 9880 10885 9908
rect 8389 9871 8447 9877
rect 10873 9877 10885 9880
rect 10919 9908 10931 9911
rect 10962 9908 10968 9920
rect 10919 9880 10968 9908
rect 10919 9877 10931 9880
rect 10873 9871 10931 9877
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 18785 9911 18843 9917
rect 18785 9877 18797 9911
rect 18831 9908 18843 9911
rect 19518 9908 19524 9920
rect 18831 9880 19524 9908
rect 18831 9877 18843 9880
rect 18785 9871 18843 9877
rect 19518 9868 19524 9880
rect 19576 9868 19582 9920
rect 20349 9911 20407 9917
rect 20349 9877 20361 9911
rect 20395 9908 20407 9911
rect 20438 9908 20444 9920
rect 20395 9880 20444 9908
rect 20395 9877 20407 9880
rect 20349 9871 20407 9877
rect 20438 9868 20444 9880
rect 20496 9868 20502 9920
rect 21192 9908 21220 10016
rect 21266 10004 21272 10056
rect 21324 10044 21330 10056
rect 23474 10044 23480 10056
rect 21324 10016 21369 10044
rect 23435 10016 23480 10044
rect 21324 10004 21330 10016
rect 23474 10004 23480 10016
rect 23532 10004 23538 10056
rect 25148 10044 25176 10084
rect 25314 10072 25320 10084
rect 25372 10072 25378 10124
rect 32677 10115 32735 10121
rect 32677 10081 32689 10115
rect 32723 10112 32735 10115
rect 33060 10112 33088 10140
rect 32723 10084 33088 10112
rect 32723 10081 32735 10084
rect 32677 10075 32735 10081
rect 26510 10044 26516 10056
rect 24504 10016 25176 10044
rect 26471 10016 26516 10044
rect 24210 9936 24216 9988
rect 24268 9976 24274 9988
rect 24504 9985 24532 10016
rect 26510 10004 26516 10016
rect 26568 10004 26574 10056
rect 28166 10044 28172 10056
rect 28127 10016 28172 10044
rect 28166 10004 28172 10016
rect 28224 10004 28230 10056
rect 28350 10044 28356 10056
rect 28311 10016 28356 10044
rect 28350 10004 28356 10016
rect 28408 10004 28414 10056
rect 28810 10004 28816 10056
rect 28868 10044 28874 10056
rect 29730 10044 29736 10056
rect 28868 10016 29736 10044
rect 28868 10004 28874 10016
rect 29730 10004 29736 10016
rect 29788 10004 29794 10056
rect 29917 10047 29975 10053
rect 29917 10013 29929 10047
rect 29963 10013 29975 10047
rect 35158 10044 35164 10056
rect 35119 10016 35164 10044
rect 29917 10007 29975 10013
rect 24489 9979 24547 9985
rect 24489 9976 24501 9979
rect 24268 9948 24501 9976
rect 24268 9936 24274 9948
rect 24489 9945 24501 9948
rect 24535 9945 24547 9979
rect 24489 9939 24547 9945
rect 22646 9908 22652 9920
rect 21192 9880 22652 9908
rect 22646 9868 22652 9880
rect 22704 9868 22710 9920
rect 23845 9911 23903 9917
rect 23845 9877 23857 9911
rect 23891 9908 23903 9911
rect 24302 9908 24308 9920
rect 23891 9880 24308 9908
rect 23891 9877 23903 9880
rect 23845 9871 23903 9877
rect 24302 9868 24308 9880
rect 24360 9868 24366 9920
rect 24762 9908 24768 9920
rect 24723 9880 24768 9908
rect 24762 9868 24768 9880
rect 24820 9868 24826 9920
rect 27801 9911 27859 9917
rect 27801 9877 27813 9911
rect 27847 9908 27859 9911
rect 27982 9908 27988 9920
rect 27847 9880 27988 9908
rect 27847 9877 27859 9880
rect 27801 9871 27859 9877
rect 27982 9868 27988 9880
rect 28040 9868 28046 9920
rect 29178 9908 29184 9920
rect 29139 9880 29184 9908
rect 29178 9868 29184 9880
rect 29236 9908 29242 9920
rect 29932 9908 29960 10007
rect 35158 10004 35164 10016
rect 35216 10004 35222 10056
rect 29236 9880 29960 9908
rect 29236 9868 29242 9880
rect 30282 9868 30288 9920
rect 30340 9908 30346 9920
rect 30377 9911 30435 9917
rect 30377 9908 30389 9911
rect 30340 9880 30389 9908
rect 30340 9868 30346 9880
rect 30377 9877 30389 9880
rect 30423 9908 30435 9911
rect 33778 9908 33784 9920
rect 30423 9880 33784 9908
rect 30423 9877 30435 9880
rect 30377 9871 30435 9877
rect 33778 9868 33784 9880
rect 33836 9908 33842 9920
rect 34057 9911 34115 9917
rect 34057 9908 34069 9911
rect 33836 9880 34069 9908
rect 33836 9868 33842 9880
rect 34057 9877 34069 9880
rect 34103 9877 34115 9911
rect 34057 9871 34115 9877
rect 34977 9911 35035 9917
rect 34977 9877 34989 9911
rect 35023 9908 35035 9911
rect 35342 9908 35348 9920
rect 35023 9880 35348 9908
rect 35023 9877 35035 9880
rect 34977 9871 35035 9877
rect 35342 9868 35348 9880
rect 35400 9868 35406 9920
rect 1104 9818 38824 9840
rect 1104 9766 7648 9818
rect 7700 9766 7712 9818
rect 7764 9766 7776 9818
rect 7828 9766 7840 9818
rect 7892 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 34315 9818
rect 34367 9766 34379 9818
rect 34431 9766 34443 9818
rect 34495 9766 34507 9818
rect 34559 9766 38824 9818
rect 1104 9744 38824 9766
rect 4249 9707 4307 9713
rect 4249 9673 4261 9707
rect 4295 9704 4307 9707
rect 4522 9704 4528 9716
rect 4295 9676 4528 9704
rect 4295 9673 4307 9676
rect 4249 9667 4307 9673
rect 4522 9664 4528 9676
rect 4580 9704 4586 9716
rect 5169 9707 5227 9713
rect 5169 9704 5181 9707
rect 4580 9676 5181 9704
rect 4580 9664 4586 9676
rect 5169 9673 5181 9676
rect 5215 9673 5227 9707
rect 5169 9667 5227 9673
rect 5902 9664 5908 9716
rect 5960 9704 5966 9716
rect 6549 9707 6607 9713
rect 6549 9704 6561 9707
rect 5960 9676 6561 9704
rect 5960 9664 5966 9676
rect 6549 9673 6561 9676
rect 6595 9673 6607 9707
rect 6549 9667 6607 9673
rect 9950 9664 9956 9716
rect 10008 9704 10014 9716
rect 10045 9707 10103 9713
rect 10045 9704 10057 9707
rect 10008 9676 10057 9704
rect 10008 9664 10014 9676
rect 10045 9673 10057 9676
rect 10091 9673 10103 9707
rect 10045 9667 10103 9673
rect 14182 9664 14188 9716
rect 14240 9704 14246 9716
rect 14369 9707 14427 9713
rect 14369 9704 14381 9707
rect 14240 9676 14381 9704
rect 14240 9664 14246 9676
rect 14369 9673 14381 9676
rect 14415 9673 14427 9707
rect 14369 9667 14427 9673
rect 14734 9664 14740 9716
rect 14792 9704 14798 9716
rect 15105 9707 15163 9713
rect 15105 9704 15117 9707
rect 14792 9676 15117 9704
rect 14792 9664 14798 9676
rect 15105 9673 15117 9676
rect 15151 9704 15163 9707
rect 15286 9704 15292 9716
rect 15151 9676 15292 9704
rect 15151 9673 15163 9676
rect 15105 9667 15163 9673
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 16390 9664 16396 9716
rect 16448 9704 16454 9716
rect 17221 9707 17279 9713
rect 17221 9704 17233 9707
rect 16448 9676 17233 9704
rect 16448 9664 16454 9676
rect 17221 9673 17233 9676
rect 17267 9704 17279 9707
rect 17310 9704 17316 9716
rect 17267 9676 17316 9704
rect 17267 9673 17279 9676
rect 17221 9667 17279 9673
rect 17310 9664 17316 9676
rect 17368 9664 17374 9716
rect 17586 9704 17592 9716
rect 17547 9676 17592 9704
rect 17586 9664 17592 9676
rect 17644 9664 17650 9716
rect 19794 9664 19800 9716
rect 19852 9704 19858 9716
rect 19852 9676 20668 9704
rect 19852 9664 19858 9676
rect 5534 9636 5540 9648
rect 5495 9608 5540 9636
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 9769 9639 9827 9645
rect 9769 9605 9781 9639
rect 9815 9636 9827 9639
rect 10226 9636 10232 9648
rect 9815 9608 10232 9636
rect 9815 9605 9827 9608
rect 9769 9599 9827 9605
rect 10226 9596 10232 9608
rect 10284 9596 10290 9648
rect 10873 9639 10931 9645
rect 10873 9605 10885 9639
rect 10919 9636 10931 9639
rect 11974 9636 11980 9648
rect 10919 9608 11980 9636
rect 10919 9605 10931 9608
rect 10873 9599 10931 9605
rect 11974 9596 11980 9608
rect 12032 9596 12038 9648
rect 13814 9636 13820 9648
rect 13775 9608 13820 9636
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 14829 9639 14887 9645
rect 14829 9605 14841 9639
rect 14875 9636 14887 9639
rect 15010 9636 15016 9648
rect 14875 9608 15016 9636
rect 14875 9605 14887 9608
rect 14829 9599 14887 9605
rect 15010 9596 15016 9608
rect 15068 9596 15074 9648
rect 18782 9636 18788 9648
rect 18743 9608 18788 9636
rect 18782 9596 18788 9608
rect 18840 9596 18846 9648
rect 20346 9636 20352 9648
rect 20307 9608 20352 9636
rect 20346 9596 20352 9608
rect 20404 9596 20410 9648
rect 20640 9636 20668 9676
rect 21266 9664 21272 9716
rect 21324 9704 21330 9716
rect 25130 9704 25136 9716
rect 21324 9676 24992 9704
rect 25091 9676 25136 9704
rect 21324 9664 21330 9676
rect 21913 9639 21971 9645
rect 21913 9636 21925 9639
rect 20640 9608 21925 9636
rect 21913 9605 21925 9608
rect 21959 9605 21971 9639
rect 23842 9636 23848 9648
rect 23803 9608 23848 9636
rect 21913 9599 21971 9605
rect 23842 9596 23848 9608
rect 23900 9596 23906 9648
rect 1854 9568 1860 9580
rect 1815 9540 1860 9568
rect 1854 9528 1860 9540
rect 1912 9528 1918 9580
rect 2682 9528 2688 9580
rect 2740 9568 2746 9580
rect 2869 9571 2927 9577
rect 2869 9568 2881 9571
rect 2740 9540 2881 9568
rect 2740 9528 2746 9540
rect 2869 9537 2881 9540
rect 2915 9537 2927 9571
rect 7009 9571 7067 9577
rect 7009 9568 7021 9571
rect 2869 9531 2927 9537
rect 5276 9540 7021 9568
rect 1578 9500 1584 9512
rect 1539 9472 1584 9500
rect 1578 9460 1584 9472
rect 1636 9500 1642 9512
rect 2774 9500 2780 9512
rect 1636 9472 2780 9500
rect 1636 9460 1642 9472
rect 2774 9460 2780 9472
rect 2832 9460 2838 9512
rect 3136 9503 3194 9509
rect 3136 9500 3148 9503
rect 3068 9472 3148 9500
rect 2409 9435 2467 9441
rect 2409 9401 2421 9435
rect 2455 9432 2467 9435
rect 3068 9432 3096 9472
rect 3136 9469 3148 9472
rect 3182 9500 3194 9503
rect 3878 9500 3884 9512
rect 3182 9472 3884 9500
rect 3182 9469 3194 9472
rect 3136 9463 3194 9469
rect 3878 9460 3884 9472
rect 3936 9460 3942 9512
rect 4706 9460 4712 9512
rect 4764 9500 4770 9512
rect 4801 9503 4859 9509
rect 4801 9500 4813 9503
rect 4764 9472 4813 9500
rect 4764 9460 4770 9472
rect 4801 9469 4813 9472
rect 4847 9500 4859 9503
rect 5276 9500 5304 9540
rect 7009 9537 7021 9540
rect 7055 9568 7067 9571
rect 7098 9568 7104 9580
rect 7055 9540 7104 9568
rect 7055 9537 7067 9540
rect 7009 9531 7067 9537
rect 7098 9528 7104 9540
rect 7156 9568 7162 9580
rect 7469 9571 7527 9577
rect 7469 9568 7481 9571
rect 7156 9540 7481 9568
rect 7156 9528 7162 9540
rect 7469 9537 7481 9540
rect 7515 9568 7527 9571
rect 7653 9571 7711 9577
rect 7653 9568 7665 9571
rect 7515 9540 7665 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 7653 9537 7665 9540
rect 7699 9537 7711 9571
rect 7653 9531 7711 9537
rect 4847 9472 5304 9500
rect 5353 9503 5411 9509
rect 4847 9469 4859 9472
rect 4801 9463 4859 9469
rect 5353 9469 5365 9503
rect 5399 9500 5411 9503
rect 5399 9472 6040 9500
rect 5399 9469 5411 9472
rect 5353 9463 5411 9469
rect 2455 9404 3096 9432
rect 2455 9401 2467 9404
rect 2409 9395 2467 9401
rect 6012 9376 6040 9472
rect 7668 9432 7696 9531
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 11422 9568 11428 9580
rect 11112 9540 11428 9568
rect 11112 9528 11118 9540
rect 11422 9528 11428 9540
rect 11480 9528 11486 9580
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9568 11943 9571
rect 15028 9568 15056 9596
rect 19337 9571 19395 9577
rect 11931 9540 12572 9568
rect 15028 9540 15424 9568
rect 11931 9537 11943 9540
rect 11885 9531 11943 9537
rect 7920 9503 7978 9509
rect 7920 9469 7932 9503
rect 7966 9500 7978 9503
rect 8202 9500 8208 9512
rect 7966 9472 8208 9500
rect 7966 9469 7978 9472
rect 7920 9463 7978 9469
rect 8202 9460 8208 9472
rect 8260 9460 8266 9512
rect 11238 9460 11244 9512
rect 11296 9500 11302 9512
rect 12158 9500 12164 9512
rect 11296 9472 12164 9500
rect 11296 9460 11302 9472
rect 12158 9460 12164 9472
rect 12216 9500 12222 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 12216 9472 12449 9500
rect 12216 9460 12222 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 8110 9432 8116 9444
rect 7668 9404 8116 9432
rect 8110 9392 8116 9404
rect 8168 9392 8174 9444
rect 11146 9432 11152 9444
rect 11059 9404 11152 9432
rect 11146 9392 11152 9404
rect 11204 9392 11210 9444
rect 12544 9432 12572 9540
rect 15102 9460 15108 9512
rect 15160 9500 15166 9512
rect 15286 9500 15292 9512
rect 15160 9472 15292 9500
rect 15160 9460 15166 9472
rect 15286 9460 15292 9472
rect 15344 9460 15350 9512
rect 15396 9500 15424 9540
rect 19337 9537 19349 9571
rect 19383 9568 19395 9571
rect 19518 9568 19524 9580
rect 19383 9540 19524 9568
rect 19383 9537 19395 9540
rect 19337 9531 19395 9537
rect 19518 9528 19524 9540
rect 19576 9528 19582 9580
rect 19797 9571 19855 9577
rect 19797 9537 19809 9571
rect 19843 9568 19855 9571
rect 19886 9568 19892 9580
rect 19843 9540 19892 9568
rect 19843 9537 19855 9540
rect 19797 9531 19855 9537
rect 19886 9528 19892 9540
rect 19944 9528 19950 9580
rect 20070 9568 20076 9580
rect 20031 9540 20076 9568
rect 20070 9528 20076 9540
rect 20128 9528 20134 9580
rect 22186 9528 22192 9580
rect 22244 9568 22250 9580
rect 22465 9571 22523 9577
rect 22465 9568 22477 9571
rect 22244 9540 22477 9568
rect 22244 9528 22250 9540
rect 22465 9537 22477 9540
rect 22511 9537 22523 9571
rect 22465 9531 22523 9537
rect 23477 9571 23535 9577
rect 23477 9537 23489 9571
rect 23523 9568 23535 9571
rect 24305 9571 24363 9577
rect 24305 9568 24317 9571
rect 23523 9540 24317 9568
rect 23523 9537 23535 9540
rect 23477 9531 23535 9537
rect 24305 9537 24317 9540
rect 24351 9568 24363 9571
rect 24670 9568 24676 9580
rect 24351 9540 24676 9568
rect 24351 9537 24363 9540
rect 24305 9531 24363 9537
rect 24670 9528 24676 9540
rect 24728 9528 24734 9580
rect 24964 9568 24992 9676
rect 25130 9664 25136 9676
rect 25188 9664 25194 9716
rect 25314 9664 25320 9716
rect 25372 9704 25378 9716
rect 25372 9676 26280 9704
rect 25372 9664 25378 9676
rect 26252 9636 26280 9676
rect 27154 9664 27160 9716
rect 27212 9704 27218 9716
rect 27212 9676 27660 9704
rect 27212 9664 27218 9676
rect 26697 9639 26755 9645
rect 26697 9636 26709 9639
rect 26252 9608 26709 9636
rect 26697 9605 26709 9608
rect 26743 9605 26755 9639
rect 26697 9599 26755 9605
rect 27433 9639 27491 9645
rect 27433 9605 27445 9639
rect 27479 9636 27491 9639
rect 27522 9636 27528 9648
rect 27479 9608 27528 9636
rect 27479 9605 27491 9608
rect 27433 9599 27491 9605
rect 27522 9596 27528 9608
rect 27580 9596 27586 9648
rect 27632 9636 27660 9676
rect 28534 9664 28540 9716
rect 28592 9704 28598 9716
rect 33045 9707 33103 9713
rect 33045 9704 33057 9707
rect 28592 9676 33057 9704
rect 28592 9664 28598 9676
rect 33045 9673 33057 9676
rect 33091 9673 33103 9707
rect 35158 9704 35164 9716
rect 33045 9667 33103 9673
rect 34440 9676 35164 9704
rect 28629 9639 28687 9645
rect 28629 9636 28641 9639
rect 27632 9608 28641 9636
rect 28629 9605 28641 9608
rect 28675 9636 28687 9639
rect 29362 9636 29368 9648
rect 28675 9608 29368 9636
rect 28675 9605 28687 9608
rect 28629 9599 28687 9605
rect 29362 9596 29368 9608
rect 29420 9636 29426 9648
rect 33060 9636 33088 9667
rect 33321 9639 33379 9645
rect 29420 9608 29592 9636
rect 33060 9608 33272 9636
rect 29420 9596 29426 9608
rect 24964 9540 25452 9568
rect 15545 9503 15603 9509
rect 15545 9500 15557 9503
rect 15396 9472 15557 9500
rect 15545 9469 15557 9472
rect 15591 9500 15603 9503
rect 16758 9500 16764 9512
rect 15591 9472 16764 9500
rect 15591 9469 15603 9472
rect 15545 9463 15603 9469
rect 16758 9460 16764 9472
rect 16816 9460 16822 9512
rect 20438 9460 20444 9512
rect 20496 9500 20502 9512
rect 20901 9503 20959 9509
rect 20901 9500 20913 9503
rect 20496 9472 20913 9500
rect 20496 9460 20502 9472
rect 20901 9469 20913 9472
rect 20947 9469 20959 9503
rect 22002 9500 22008 9512
rect 20901 9463 20959 9469
rect 21192 9472 22008 9500
rect 12710 9441 12716 9444
rect 12704 9432 12716 9441
rect 12544 9404 12716 9432
rect 12704 9395 12716 9404
rect 12710 9392 12716 9395
rect 12768 9392 12774 9444
rect 18874 9392 18880 9444
rect 18932 9432 18938 9444
rect 19061 9435 19119 9441
rect 19061 9432 19073 9435
rect 18932 9404 19073 9432
rect 18932 9392 18938 9404
rect 19061 9401 19073 9404
rect 19107 9401 19119 9435
rect 19061 9395 19119 9401
rect 20625 9435 20683 9441
rect 20625 9401 20637 9435
rect 20671 9432 20683 9435
rect 20714 9432 20720 9444
rect 20671 9404 20720 9432
rect 20671 9401 20683 9404
rect 20625 9395 20683 9401
rect 20714 9392 20720 9404
rect 20772 9392 20778 9444
rect 21192 9432 21220 9472
rect 22002 9460 22008 9472
rect 22060 9460 22066 9512
rect 23109 9503 23167 9509
rect 23109 9469 23121 9503
rect 23155 9500 23167 9503
rect 24397 9503 24455 9509
rect 24397 9500 24409 9503
rect 23155 9472 24409 9500
rect 23155 9469 23167 9472
rect 23109 9463 23167 9469
rect 24397 9469 24409 9472
rect 24443 9500 24455 9503
rect 25222 9500 25228 9512
rect 24443 9472 25228 9500
rect 24443 9469 24455 9472
rect 24397 9463 24455 9469
rect 25222 9460 25228 9472
rect 25280 9460 25286 9512
rect 25317 9503 25375 9509
rect 25317 9469 25329 9503
rect 25363 9469 25375 9503
rect 25317 9463 25375 9469
rect 22189 9435 22247 9441
rect 22189 9432 22201 9435
rect 20824 9404 21220 9432
rect 21284 9404 22201 9432
rect 2682 9364 2688 9376
rect 2643 9336 2688 9364
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 5994 9364 6000 9376
rect 5955 9336 6000 9364
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 9030 9364 9036 9376
rect 8991 9336 9036 9364
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 10594 9364 10600 9376
rect 10555 9336 10600 9364
rect 10594 9324 10600 9336
rect 10652 9364 10658 9376
rect 11164 9364 11192 9392
rect 10652 9336 11192 9364
rect 11333 9367 11391 9373
rect 10652 9324 10658 9336
rect 11333 9333 11345 9367
rect 11379 9364 11391 9367
rect 11422 9364 11428 9376
rect 11379 9336 11428 9364
rect 11379 9333 11391 9336
rect 11333 9327 11391 9333
rect 11422 9324 11428 9336
rect 11480 9324 11486 9376
rect 16666 9364 16672 9376
rect 16627 9336 16672 9364
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 18322 9324 18328 9376
rect 18380 9364 18386 9376
rect 18509 9367 18567 9373
rect 18509 9364 18521 9367
rect 18380 9336 18521 9364
rect 18380 9324 18386 9336
rect 18509 9333 18521 9336
rect 18555 9364 18567 9367
rect 19245 9367 19303 9373
rect 19245 9364 19257 9367
rect 18555 9336 19257 9364
rect 18555 9333 18567 9336
rect 18509 9327 18567 9333
rect 19245 9333 19257 9336
rect 19291 9364 19303 9367
rect 19426 9364 19432 9376
rect 19291 9336 19432 9364
rect 19291 9333 19303 9336
rect 19245 9327 19303 9333
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 20070 9324 20076 9376
rect 20128 9364 20134 9376
rect 20824 9373 20852 9404
rect 21284 9376 21312 9404
rect 22189 9401 22201 9404
rect 22235 9432 22247 9435
rect 23474 9432 23480 9444
rect 22235 9404 23480 9432
rect 22235 9401 22247 9404
rect 22189 9395 22247 9401
rect 23474 9392 23480 9404
rect 23532 9392 23538 9444
rect 24302 9432 24308 9444
rect 24263 9404 24308 9432
rect 24302 9392 24308 9404
rect 24360 9392 24366 9444
rect 25130 9392 25136 9444
rect 25188 9432 25194 9444
rect 25332 9432 25360 9463
rect 25188 9404 25360 9432
rect 25188 9392 25194 9404
rect 20809 9367 20867 9373
rect 20809 9364 20821 9367
rect 20128 9336 20821 9364
rect 20128 9324 20134 9336
rect 20809 9333 20821 9336
rect 20855 9333 20867 9367
rect 21266 9364 21272 9376
rect 21227 9336 21272 9364
rect 20809 9327 20867 9333
rect 21266 9324 21272 9336
rect 21324 9324 21330 9376
rect 21726 9364 21732 9376
rect 21639 9336 21732 9364
rect 21726 9324 21732 9336
rect 21784 9364 21790 9376
rect 22370 9364 22376 9376
rect 21784 9336 22376 9364
rect 21784 9324 21790 9336
rect 22370 9324 22376 9336
rect 22428 9324 22434 9376
rect 24857 9367 24915 9373
rect 24857 9333 24869 9367
rect 24903 9364 24915 9367
rect 24946 9364 24952 9376
rect 24903 9336 24952 9364
rect 24903 9333 24915 9336
rect 24857 9327 24915 9333
rect 24946 9324 24952 9336
rect 25004 9324 25010 9376
rect 25424 9364 25452 9540
rect 28902 9528 28908 9580
rect 28960 9568 28966 9580
rect 29089 9571 29147 9577
rect 29089 9568 29101 9571
rect 28960 9540 29101 9568
rect 28960 9528 28966 9540
rect 29089 9537 29101 9540
rect 29135 9568 29147 9571
rect 29270 9568 29276 9580
rect 29135 9540 29276 9568
rect 29135 9537 29147 9540
rect 29089 9531 29147 9537
rect 29270 9528 29276 9540
rect 29328 9528 29334 9580
rect 29564 9577 29592 9608
rect 29549 9571 29607 9577
rect 29549 9537 29561 9571
rect 29595 9537 29607 9571
rect 29549 9531 29607 9537
rect 32033 9571 32091 9577
rect 32033 9537 32045 9571
rect 32079 9568 32091 9571
rect 33042 9568 33048 9580
rect 32079 9540 33048 9568
rect 32079 9537 32091 9540
rect 32033 9531 32091 9537
rect 33042 9528 33048 9540
rect 33100 9528 33106 9580
rect 25590 9509 25596 9512
rect 25584 9500 25596 9509
rect 25503 9472 25596 9500
rect 25584 9463 25596 9472
rect 25648 9500 25654 9512
rect 26142 9500 26148 9512
rect 25648 9472 26148 9500
rect 25590 9460 25596 9463
rect 25648 9460 25654 9472
rect 26142 9460 26148 9472
rect 26200 9460 26206 9512
rect 29816 9503 29874 9509
rect 29816 9469 29828 9503
rect 29862 9500 29874 9503
rect 30282 9500 30288 9512
rect 29862 9472 30288 9500
rect 29862 9469 29874 9472
rect 29816 9463 29874 9469
rect 30282 9460 30288 9472
rect 30340 9460 30346 9512
rect 32122 9500 32128 9512
rect 32035 9472 32128 9500
rect 32122 9460 32128 9472
rect 32180 9500 32186 9512
rect 32180 9472 32812 9500
rect 32180 9460 32186 9472
rect 26602 9392 26608 9444
rect 26660 9432 26666 9444
rect 28077 9435 28135 9441
rect 28077 9432 28089 9435
rect 26660 9404 28089 9432
rect 26660 9392 26666 9404
rect 28077 9401 28089 9404
rect 28123 9432 28135 9435
rect 28350 9432 28356 9444
rect 28123 9404 28356 9432
rect 28123 9401 28135 9404
rect 28077 9395 28135 9401
rect 28350 9392 28356 9404
rect 28408 9432 28414 9444
rect 29086 9432 29092 9444
rect 28408 9404 29092 9432
rect 28408 9392 28414 9404
rect 29086 9392 29092 9404
rect 29144 9392 29150 9444
rect 32784 9376 32812 9472
rect 27709 9367 27767 9373
rect 27709 9364 27721 9367
rect 25424 9336 27721 9364
rect 27709 9333 27721 9336
rect 27755 9364 27767 9367
rect 28166 9364 28172 9376
rect 27755 9336 28172 9364
rect 27755 9333 27767 9336
rect 27709 9327 27767 9333
rect 28166 9324 28172 9336
rect 28224 9324 28230 9376
rect 29178 9324 29184 9376
rect 29236 9364 29242 9376
rect 30929 9367 30987 9373
rect 30929 9364 30941 9367
rect 29236 9336 30941 9364
rect 29236 9324 29242 9336
rect 30929 9333 30941 9336
rect 30975 9333 30987 9367
rect 32306 9364 32312 9376
rect 32267 9336 32312 9364
rect 30929 9327 30987 9333
rect 32306 9324 32312 9336
rect 32364 9324 32370 9376
rect 32766 9364 32772 9376
rect 32727 9336 32772 9364
rect 32766 9324 32772 9336
rect 32824 9324 32830 9376
rect 33244 9364 33272 9608
rect 33321 9605 33333 9639
rect 33367 9605 33379 9639
rect 33321 9599 33379 9605
rect 33336 9500 33364 9599
rect 33962 9596 33968 9648
rect 34020 9636 34026 9648
rect 34440 9636 34468 9676
rect 35158 9664 35164 9676
rect 35216 9704 35222 9716
rect 35216 9676 35940 9704
rect 35216 9664 35222 9676
rect 34020 9608 34468 9636
rect 34020 9596 34026 9608
rect 34606 9596 34612 9648
rect 34664 9636 34670 9648
rect 35912 9645 35940 9676
rect 34977 9639 35035 9645
rect 34977 9636 34989 9639
rect 34664 9608 34989 9636
rect 34664 9596 34670 9608
rect 34977 9605 34989 9608
rect 35023 9605 35035 9639
rect 34977 9599 35035 9605
rect 35897 9639 35955 9645
rect 35897 9605 35909 9639
rect 35943 9605 35955 9639
rect 35897 9599 35955 9605
rect 33778 9528 33784 9580
rect 33836 9568 33842 9580
rect 37550 9568 37556 9580
rect 33836 9540 36492 9568
rect 37511 9540 37556 9568
rect 33836 9528 33842 9540
rect 33336 9472 35480 9500
rect 35452 9444 35480 9472
rect 35526 9460 35532 9512
rect 35584 9500 35590 9512
rect 36464 9509 36492 9540
rect 37550 9528 37556 9540
rect 37608 9528 37614 9580
rect 36265 9503 36323 9509
rect 36265 9500 36277 9503
rect 35584 9472 36277 9500
rect 35584 9460 35590 9472
rect 36265 9469 36277 9472
rect 36311 9469 36323 9503
rect 36265 9463 36323 9469
rect 36449 9503 36507 9509
rect 36449 9469 36461 9503
rect 36495 9500 36507 9503
rect 37001 9503 37059 9509
rect 37001 9500 37013 9503
rect 36495 9472 37013 9500
rect 36495 9469 36507 9472
rect 36449 9463 36507 9469
rect 37001 9469 37013 9472
rect 37047 9469 37059 9503
rect 37001 9463 37059 9469
rect 33502 9392 33508 9444
rect 33560 9432 33566 9444
rect 33597 9435 33655 9441
rect 33597 9432 33609 9435
rect 33560 9404 33609 9432
rect 33560 9392 33566 9404
rect 33597 9401 33609 9404
rect 33643 9401 33655 9435
rect 33870 9432 33876 9444
rect 33831 9404 33876 9432
rect 33597 9395 33655 9401
rect 33870 9392 33876 9404
rect 33928 9392 33934 9444
rect 35250 9432 35256 9444
rect 35163 9404 35256 9432
rect 35250 9392 35256 9404
rect 35308 9392 35314 9444
rect 35434 9432 35440 9444
rect 35347 9404 35440 9432
rect 35434 9392 35440 9404
rect 35492 9392 35498 9444
rect 33778 9364 33784 9376
rect 33244 9336 33784 9364
rect 33778 9324 33784 9336
rect 33836 9324 33842 9376
rect 34333 9367 34391 9373
rect 34333 9333 34345 9367
rect 34379 9364 34391 9367
rect 34422 9364 34428 9376
rect 34379 9336 34428 9364
rect 34379 9333 34391 9336
rect 34333 9327 34391 9333
rect 34422 9324 34428 9336
rect 34480 9324 34486 9376
rect 34606 9364 34612 9376
rect 34567 9336 34612 9364
rect 34606 9324 34612 9336
rect 34664 9364 34670 9376
rect 35268 9364 35296 9392
rect 34664 9336 35296 9364
rect 36633 9367 36691 9373
rect 34664 9324 34670 9336
rect 36633 9333 36645 9367
rect 36679 9364 36691 9367
rect 36906 9364 36912 9376
rect 36679 9336 36912 9364
rect 36679 9333 36691 9336
rect 36633 9327 36691 9333
rect 36906 9324 36912 9336
rect 36964 9324 36970 9376
rect 1104 9274 38824 9296
rect 1104 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 27648 9274
rect 27700 9222 27712 9274
rect 27764 9222 27776 9274
rect 27828 9222 27840 9274
rect 27892 9222 38824 9274
rect 1104 9200 38824 9222
rect 3970 9120 3976 9172
rect 4028 9160 4034 9172
rect 4249 9163 4307 9169
rect 4249 9160 4261 9163
rect 4028 9132 4261 9160
rect 4028 9120 4034 9132
rect 4249 9129 4261 9132
rect 4295 9129 4307 9163
rect 4614 9160 4620 9172
rect 4575 9132 4620 9160
rect 4249 9123 4307 9129
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 4982 9160 4988 9172
rect 4943 9132 4988 9160
rect 4982 9120 4988 9132
rect 5040 9120 5046 9172
rect 8202 9160 8208 9172
rect 7760 9132 8208 9160
rect 1949 9095 2007 9101
rect 1949 9061 1961 9095
rect 1995 9092 2007 9095
rect 3053 9095 3111 9101
rect 3053 9092 3065 9095
rect 1995 9064 3065 9092
rect 1995 9061 2007 9064
rect 1949 9055 2007 9061
rect 3053 9061 3065 9064
rect 3099 9061 3111 9095
rect 6086 9092 6092 9104
rect 6047 9064 6092 9092
rect 3053 9055 3111 9061
rect 6086 9052 6092 9064
rect 6144 9052 6150 9104
rect 7282 9052 7288 9104
rect 7340 9092 7346 9104
rect 7466 9092 7472 9104
rect 7340 9064 7472 9092
rect 7340 9052 7346 9064
rect 7466 9052 7472 9064
rect 7524 9092 7530 9104
rect 7760 9101 7788 9132
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 9490 9160 9496 9172
rect 9451 9132 9496 9160
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 11330 9160 11336 9172
rect 11291 9132 11336 9160
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 14090 9160 14096 9172
rect 14051 9132 14096 9160
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 17586 9120 17592 9172
rect 17644 9160 17650 9172
rect 17865 9163 17923 9169
rect 17865 9160 17877 9163
rect 17644 9132 17877 9160
rect 17644 9120 17650 9132
rect 17865 9129 17877 9132
rect 17911 9129 17923 9163
rect 17865 9123 17923 9129
rect 19153 9163 19211 9169
rect 19153 9129 19165 9163
rect 19199 9160 19211 9163
rect 19334 9160 19340 9172
rect 19199 9132 19340 9160
rect 19199 9129 19211 9132
rect 19153 9123 19211 9129
rect 19334 9120 19340 9132
rect 19392 9120 19398 9172
rect 20346 9120 20352 9172
rect 20404 9160 20410 9172
rect 20625 9163 20683 9169
rect 20625 9160 20637 9163
rect 20404 9132 20637 9160
rect 20404 9120 20410 9132
rect 20625 9129 20637 9132
rect 20671 9160 20683 9163
rect 20671 9132 21312 9160
rect 20671 9129 20683 9132
rect 20625 9123 20683 9129
rect 7653 9095 7711 9101
rect 7653 9092 7665 9095
rect 7524 9064 7665 9092
rect 7524 9052 7530 9064
rect 7653 9061 7665 9064
rect 7699 9061 7711 9095
rect 7653 9055 7711 9061
rect 7745 9095 7803 9101
rect 7745 9061 7757 9095
rect 7791 9061 7803 9095
rect 7745 9055 7803 9061
rect 10229 9095 10287 9101
rect 10229 9061 10241 9095
rect 10275 9092 10287 9095
rect 10962 9092 10968 9104
rect 10275 9064 10968 9092
rect 10275 9061 10287 9064
rect 10229 9055 10287 9061
rect 10962 9052 10968 9064
rect 11020 9052 11026 9104
rect 11422 9052 11428 9104
rect 11480 9052 11486 9104
rect 11698 9101 11704 9104
rect 11681 9095 11704 9101
rect 11681 9061 11693 9095
rect 11681 9055 11704 9061
rect 11698 9052 11704 9055
rect 11756 9052 11762 9104
rect 19794 9092 19800 9104
rect 19755 9064 19800 9092
rect 19794 9052 19800 9064
rect 19852 9052 19858 9104
rect 21284 9101 21312 9132
rect 22186 9120 22192 9172
rect 22244 9160 22250 9172
rect 22281 9163 22339 9169
rect 22281 9160 22293 9163
rect 22244 9132 22293 9160
rect 22244 9120 22250 9132
rect 22281 9129 22293 9132
rect 22327 9129 22339 9163
rect 25590 9160 25596 9172
rect 25551 9132 25596 9160
rect 22281 9123 22339 9129
rect 25590 9120 25596 9132
rect 25648 9120 25654 9172
rect 27154 9160 27160 9172
rect 27115 9132 27160 9160
rect 27154 9120 27160 9132
rect 27212 9120 27218 9172
rect 27709 9163 27767 9169
rect 27709 9129 27721 9163
rect 27755 9160 27767 9163
rect 27982 9160 27988 9172
rect 27755 9132 27988 9160
rect 27755 9129 27767 9132
rect 27709 9123 27767 9129
rect 27982 9120 27988 9132
rect 28040 9120 28046 9172
rect 30926 9160 30932 9172
rect 30887 9132 30932 9160
rect 30926 9120 30932 9132
rect 30984 9120 30990 9172
rect 35434 9120 35440 9172
rect 35492 9160 35498 9172
rect 36449 9163 36507 9169
rect 36449 9160 36461 9163
rect 35492 9132 36461 9160
rect 35492 9120 35498 9132
rect 36449 9129 36461 9132
rect 36495 9129 36507 9163
rect 36449 9123 36507 9129
rect 21269 9095 21327 9101
rect 21269 9061 21281 9095
rect 21315 9061 21327 9095
rect 21269 9055 21327 9061
rect 21453 9095 21511 9101
rect 21453 9061 21465 9095
rect 21499 9061 21511 9095
rect 21453 9055 21511 9061
rect 3513 9027 3571 9033
rect 3513 9024 3525 9027
rect 1964 8996 3525 9024
rect 1964 8968 1992 8996
rect 3513 8993 3525 8996
rect 3559 8993 3571 9027
rect 3513 8987 3571 8993
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 9024 4123 9027
rect 4614 9024 4620 9036
rect 4111 8996 4620 9024
rect 4111 8993 4123 8996
rect 4065 8987 4123 8993
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 5445 9027 5503 9033
rect 5445 8993 5457 9027
rect 5491 9024 5503 9027
rect 6181 9027 6239 9033
rect 6181 9024 6193 9027
rect 5491 8996 6193 9024
rect 5491 8993 5503 8996
rect 5445 8987 5503 8993
rect 6181 8993 6193 8996
rect 6227 9024 6239 9027
rect 6730 9024 6736 9036
rect 6227 8996 6736 9024
rect 6227 8993 6239 8996
rect 6181 8987 6239 8993
rect 6730 8984 6736 8996
rect 6788 9024 6794 9036
rect 6917 9027 6975 9033
rect 6917 9024 6929 9027
rect 6788 8996 6929 9024
rect 6788 8984 6794 8996
rect 6917 8993 6929 8996
rect 6963 9024 6975 9027
rect 8573 9027 8631 9033
rect 8573 9024 8585 9027
rect 6963 8996 8585 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 8573 8993 8585 8996
rect 8619 9024 8631 9027
rect 9030 9024 9036 9036
rect 8619 8996 9036 9024
rect 8619 8993 8631 8996
rect 8573 8987 8631 8993
rect 9030 8984 9036 8996
rect 9088 9024 9094 9036
rect 10321 9027 10379 9033
rect 10321 9024 10333 9027
rect 9088 8996 10333 9024
rect 9088 8984 9094 8996
rect 10321 8993 10333 8996
rect 10367 8993 10379 9027
rect 10321 8987 10379 8993
rect 10410 8984 10416 9036
rect 10468 9024 10474 9036
rect 10873 9027 10931 9033
rect 10873 9024 10885 9027
rect 10468 8996 10885 9024
rect 10468 8984 10474 8996
rect 10873 8993 10885 8996
rect 10919 9024 10931 9027
rect 11440 9024 11468 9052
rect 10919 8996 11468 9024
rect 16752 9027 16810 9033
rect 10919 8993 10931 8996
rect 10873 8987 10931 8993
rect 16752 8993 16764 9027
rect 16798 9024 16810 9027
rect 17126 9024 17132 9036
rect 16798 8996 17132 9024
rect 16798 8993 16810 8996
rect 16752 8987 16810 8993
rect 17126 8984 17132 8996
rect 17184 8984 17190 9036
rect 19426 8984 19432 9036
rect 19484 9024 19490 9036
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 19484 8996 19625 9024
rect 19484 8984 19490 8996
rect 19613 8993 19625 8996
rect 19659 9024 19671 9027
rect 19978 9024 19984 9036
rect 19659 8996 19984 9024
rect 19659 8993 19671 8996
rect 19613 8987 19671 8993
rect 19978 8984 19984 8996
rect 20036 8984 20042 9036
rect 21468 9024 21496 9055
rect 21634 9052 21640 9104
rect 21692 9092 21698 9104
rect 22833 9095 22891 9101
rect 21692 9064 22324 9092
rect 21692 9052 21698 9064
rect 20824 8996 21496 9024
rect 21545 9027 21603 9033
rect 1946 8956 1952 8968
rect 1907 8928 1952 8956
rect 1946 8916 1952 8928
rect 2004 8916 2010 8968
rect 2041 8959 2099 8965
rect 2041 8925 2053 8959
rect 2087 8956 2099 8959
rect 2406 8956 2412 8968
rect 2087 8928 2412 8956
rect 2087 8925 2099 8928
rect 2041 8919 2099 8925
rect 2406 8916 2412 8928
rect 2464 8916 2470 8968
rect 2682 8916 2688 8968
rect 2740 8956 2746 8968
rect 4706 8956 4712 8968
rect 2740 8928 4712 8956
rect 2740 8916 2746 8928
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 6086 8956 6092 8968
rect 6047 8928 6092 8956
rect 6086 8916 6092 8928
rect 6144 8916 6150 8968
rect 6546 8916 6552 8968
rect 6604 8956 6610 8968
rect 7650 8956 7656 8968
rect 6604 8928 7656 8956
rect 6604 8916 6610 8928
rect 7650 8916 7656 8928
rect 7708 8916 7714 8968
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8956 10287 8959
rect 10502 8956 10508 8968
rect 10275 8928 10508 8956
rect 10275 8925 10287 8928
rect 10229 8919 10287 8925
rect 10502 8916 10508 8928
rect 10560 8916 10566 8968
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 11425 8959 11483 8965
rect 11425 8956 11437 8959
rect 11296 8928 11437 8956
rect 11296 8916 11302 8928
rect 11425 8925 11437 8928
rect 11471 8925 11483 8959
rect 11425 8919 11483 8925
rect 15102 8916 15108 8968
rect 15160 8956 15166 8968
rect 16485 8959 16543 8965
rect 16485 8956 16497 8959
rect 15160 8928 16497 8956
rect 15160 8916 15166 8928
rect 16485 8925 16497 8928
rect 16531 8925 16543 8959
rect 16485 8919 16543 8925
rect 19889 8959 19947 8965
rect 19889 8925 19901 8959
rect 19935 8956 19947 8959
rect 20346 8956 20352 8968
rect 19935 8928 20352 8956
rect 19935 8925 19947 8928
rect 19889 8919 19947 8925
rect 20346 8916 20352 8928
rect 20404 8916 20410 8968
rect 20824 8900 20852 8996
rect 21545 8993 21557 9027
rect 21591 9024 21603 9027
rect 22186 9024 22192 9036
rect 21591 8996 22192 9024
rect 21591 8993 21603 8996
rect 21545 8987 21603 8993
rect 22186 8984 22192 8996
rect 22244 8984 22250 9036
rect 22296 9024 22324 9064
rect 22833 9061 22845 9095
rect 22879 9092 22891 9095
rect 23477 9095 23535 9101
rect 23477 9092 23489 9095
rect 22879 9064 23489 9092
rect 22879 9061 22891 9064
rect 22833 9055 22891 9061
rect 23477 9061 23489 9064
rect 23523 9092 23535 9095
rect 24563 9095 24621 9101
rect 24563 9092 24575 9095
rect 23523 9064 24575 9092
rect 23523 9061 23535 9064
rect 23477 9055 23535 9061
rect 24563 9061 24575 9064
rect 24609 9061 24621 9095
rect 24563 9055 24621 9061
rect 24854 9052 24860 9104
rect 24912 9092 24918 9104
rect 25041 9095 25099 9101
rect 25041 9092 25053 9095
rect 24912 9064 25053 9092
rect 24912 9052 24918 9064
rect 25041 9061 25053 9064
rect 25087 9061 25099 9095
rect 25041 9055 25099 9061
rect 25222 9052 25228 9104
rect 25280 9092 25286 9104
rect 26053 9095 26111 9101
rect 26053 9092 26065 9095
rect 25280 9064 26065 9092
rect 25280 9052 25286 9064
rect 26053 9061 26065 9064
rect 26099 9092 26111 9095
rect 26602 9092 26608 9104
rect 26099 9064 26608 9092
rect 26099 9061 26111 9064
rect 26053 9055 26111 9061
rect 26602 9052 26608 9064
rect 26660 9052 26666 9104
rect 27172 9092 27200 9120
rect 28077 9095 28135 9101
rect 28077 9092 28089 9095
rect 27172 9064 28089 9092
rect 28077 9061 28089 9064
rect 28123 9061 28135 9095
rect 28077 9055 28135 9061
rect 31846 9052 31852 9104
rect 31904 9092 31910 9104
rect 33137 9095 33195 9101
rect 33137 9092 33149 9095
rect 31904 9064 33149 9092
rect 31904 9052 31910 9064
rect 33137 9061 33149 9064
rect 33183 9061 33195 9095
rect 33137 9055 33195 9061
rect 23293 9027 23351 9033
rect 23293 9024 23305 9027
rect 22296 8996 23305 9024
rect 23293 8993 23305 8996
rect 23339 8993 23351 9027
rect 23293 8987 23351 8993
rect 26142 8984 26148 9036
rect 26200 9024 26206 9036
rect 26973 9027 27031 9033
rect 26973 9024 26985 9027
rect 26200 8996 26985 9024
rect 26200 8984 26206 8996
rect 26973 8993 26985 8996
rect 27019 9024 27031 9027
rect 28353 9027 28411 9033
rect 28353 9024 28365 9027
rect 27019 8996 28365 9024
rect 27019 8993 27031 8996
rect 26973 8987 27031 8993
rect 28353 8993 28365 8996
rect 28399 8993 28411 9027
rect 28353 8987 28411 8993
rect 28718 8984 28724 9036
rect 28776 9024 28782 9036
rect 29178 9024 29184 9036
rect 28776 8996 29184 9024
rect 28776 8984 28782 8996
rect 29178 8984 29184 8996
rect 29236 9024 29242 9036
rect 29805 9027 29863 9033
rect 29805 9024 29817 9027
rect 29236 8996 29817 9024
rect 29236 8984 29242 8996
rect 29805 8993 29817 8996
rect 29851 8993 29863 9027
rect 29805 8987 29863 8993
rect 32493 9027 32551 9033
rect 32493 8993 32505 9027
rect 32539 9024 32551 9027
rect 32950 9024 32956 9036
rect 32539 8996 32956 9024
rect 32539 8993 32551 8996
rect 32493 8987 32551 8993
rect 32950 8984 32956 8996
rect 33008 8984 33014 9036
rect 33870 8984 33876 9036
rect 33928 9024 33934 9036
rect 34422 9033 34428 9036
rect 34416 9024 34428 9033
rect 33928 8996 34428 9024
rect 33928 8984 33934 8996
rect 34416 8987 34428 8996
rect 34480 9024 34486 9036
rect 35894 9024 35900 9036
rect 34480 8996 35900 9024
rect 34422 8984 34428 8987
rect 34480 8984 34486 8996
rect 35894 8984 35900 8996
rect 35952 8984 35958 9036
rect 23566 8956 23572 8968
rect 23527 8928 23572 8956
rect 23566 8916 23572 8928
rect 23624 8916 23630 8968
rect 24302 8916 24308 8968
rect 24360 8956 24366 8968
rect 24949 8959 25007 8965
rect 24949 8956 24961 8959
rect 24360 8928 24961 8956
rect 24360 8916 24366 8928
rect 24949 8925 24961 8928
rect 24995 8925 25007 8959
rect 25130 8956 25136 8968
rect 25091 8928 25136 8956
rect 24949 8919 25007 8925
rect 25130 8916 25136 8928
rect 25188 8916 25194 8968
rect 27246 8956 27252 8968
rect 27207 8928 27252 8956
rect 27246 8916 27252 8928
rect 27304 8916 27310 8968
rect 29362 8916 29368 8968
rect 29420 8956 29426 8968
rect 29546 8956 29552 8968
rect 29420 8928 29552 8956
rect 29420 8916 29426 8928
rect 29546 8916 29552 8928
rect 29604 8916 29610 8968
rect 33226 8956 33232 8968
rect 33187 8928 33232 8956
rect 33226 8916 33232 8928
rect 33284 8916 33290 8968
rect 33962 8916 33968 8968
rect 34020 8956 34026 8968
rect 34149 8959 34207 8965
rect 34149 8956 34161 8959
rect 34020 8928 34161 8956
rect 34020 8916 34026 8928
rect 34149 8925 34161 8928
rect 34195 8925 34207 8959
rect 36630 8956 36636 8968
rect 36591 8928 36636 8956
rect 34149 8919 34207 8925
rect 36630 8916 36636 8928
rect 36688 8916 36694 8968
rect 1486 8888 1492 8900
rect 1447 8860 1492 8888
rect 1486 8848 1492 8860
rect 1544 8848 1550 8900
rect 2869 8891 2927 8897
rect 2869 8857 2881 8891
rect 2915 8888 2927 8891
rect 3142 8888 3148 8900
rect 2915 8860 3148 8888
rect 2915 8857 2927 8860
rect 2869 8851 2927 8857
rect 3142 8848 3148 8860
rect 3200 8848 3206 8900
rect 5629 8891 5687 8897
rect 5629 8857 5641 8891
rect 5675 8888 5687 8891
rect 5718 8888 5724 8900
rect 5675 8860 5724 8888
rect 5675 8857 5687 8860
rect 5629 8851 5687 8857
rect 5718 8848 5724 8860
rect 5776 8888 5782 8900
rect 6454 8888 6460 8900
rect 5776 8860 6460 8888
rect 5776 8848 5782 8860
rect 6454 8848 6460 8860
rect 6512 8848 6518 8900
rect 19337 8891 19395 8897
rect 19337 8857 19349 8891
rect 19383 8888 19395 8891
rect 20806 8888 20812 8900
rect 19383 8860 20812 8888
rect 19383 8857 19395 8860
rect 19337 8851 19395 8857
rect 20806 8848 20812 8860
rect 20864 8848 20870 8900
rect 23014 8888 23020 8900
rect 22975 8860 23020 8888
rect 23014 8848 23020 8860
rect 23072 8848 23078 8900
rect 35526 8888 35532 8900
rect 35487 8860 35532 8888
rect 35526 8848 35532 8860
rect 35584 8888 35590 8900
rect 36081 8891 36139 8897
rect 36081 8888 36093 8891
rect 35584 8860 36093 8888
rect 35584 8848 35590 8860
rect 36081 8857 36093 8860
rect 36127 8857 36139 8891
rect 36081 8851 36139 8857
rect 1302 8780 1308 8832
rect 1360 8820 1366 8832
rect 2958 8820 2964 8832
rect 1360 8792 2964 8820
rect 1360 8780 1366 8792
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 3053 8823 3111 8829
rect 3053 8789 3065 8823
rect 3099 8820 3111 8823
rect 3237 8823 3295 8829
rect 3237 8820 3249 8823
rect 3099 8792 3249 8820
rect 3099 8789 3111 8792
rect 3053 8783 3111 8789
rect 3237 8789 3249 8792
rect 3283 8820 3295 8823
rect 4338 8820 4344 8832
rect 3283 8792 4344 8820
rect 3283 8789 3295 8792
rect 3237 8783 3295 8789
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 6641 8823 6699 8829
rect 6641 8789 6653 8823
rect 6687 8820 6699 8823
rect 7193 8823 7251 8829
rect 7193 8820 7205 8823
rect 6687 8792 7205 8820
rect 6687 8789 6699 8792
rect 6641 8783 6699 8789
rect 7193 8789 7205 8792
rect 7239 8820 7251 8823
rect 7466 8820 7472 8832
rect 7239 8792 7472 8820
rect 7239 8789 7251 8792
rect 7193 8783 7251 8789
rect 7466 8780 7472 8792
rect 7524 8780 7530 8832
rect 9766 8820 9772 8832
rect 9727 8792 9772 8820
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 12158 8780 12164 8832
rect 12216 8820 12222 8832
rect 12805 8823 12863 8829
rect 12805 8820 12817 8823
rect 12216 8792 12817 8820
rect 12216 8780 12222 8792
rect 12805 8789 12817 8792
rect 12851 8789 12863 8823
rect 12805 8783 12863 8789
rect 13725 8823 13783 8829
rect 13725 8789 13737 8823
rect 13771 8820 13783 8823
rect 13814 8820 13820 8832
rect 13771 8792 13820 8820
rect 13771 8789 13783 8792
rect 13725 8783 13783 8789
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 18785 8823 18843 8829
rect 18785 8789 18797 8823
rect 18831 8820 18843 8823
rect 18874 8820 18880 8832
rect 18831 8792 18880 8820
rect 18831 8789 18843 8792
rect 18785 8783 18843 8789
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 20349 8823 20407 8829
rect 20349 8789 20361 8823
rect 20395 8820 20407 8823
rect 20714 8820 20720 8832
rect 20395 8792 20720 8820
rect 20395 8789 20407 8792
rect 20349 8783 20407 8789
rect 20714 8780 20720 8792
rect 20772 8780 20778 8832
rect 20993 8823 21051 8829
rect 20993 8789 21005 8823
rect 21039 8820 21051 8823
rect 21634 8820 21640 8832
rect 21039 8792 21640 8820
rect 21039 8789 21051 8792
rect 20993 8783 21051 8789
rect 21634 8780 21640 8792
rect 21692 8780 21698 8832
rect 21910 8820 21916 8832
rect 21871 8792 21916 8820
rect 21910 8780 21916 8792
rect 21968 8780 21974 8832
rect 24210 8820 24216 8832
rect 24171 8792 24216 8820
rect 24210 8780 24216 8792
rect 24268 8780 24274 8832
rect 26694 8820 26700 8832
rect 26655 8792 26700 8820
rect 26694 8780 26700 8792
rect 26752 8780 26758 8832
rect 28902 8820 28908 8832
rect 28863 8792 28908 8820
rect 28902 8780 28908 8792
rect 28960 8780 28966 8832
rect 29365 8823 29423 8829
rect 29365 8789 29377 8823
rect 29411 8820 29423 8823
rect 29730 8820 29736 8832
rect 29411 8792 29736 8820
rect 29411 8789 29423 8792
rect 29365 8783 29423 8789
rect 29730 8780 29736 8792
rect 29788 8780 29794 8832
rect 32677 8823 32735 8829
rect 32677 8789 32689 8823
rect 32723 8820 32735 8823
rect 33134 8820 33140 8832
rect 32723 8792 33140 8820
rect 32723 8789 32735 8792
rect 32677 8783 32735 8789
rect 33134 8780 33140 8792
rect 33192 8780 33198 8832
rect 33502 8780 33508 8832
rect 33560 8820 33566 8832
rect 33597 8823 33655 8829
rect 33597 8820 33609 8823
rect 33560 8792 33609 8820
rect 33560 8780 33566 8792
rect 33597 8789 33609 8792
rect 33643 8789 33655 8823
rect 34054 8820 34060 8832
rect 34015 8792 34060 8820
rect 33597 8783 33655 8789
rect 34054 8780 34060 8792
rect 34112 8780 34118 8832
rect 1104 8730 38824 8752
rect 1104 8678 7648 8730
rect 7700 8678 7712 8730
rect 7764 8678 7776 8730
rect 7828 8678 7840 8730
rect 7892 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 34315 8730
rect 34367 8678 34379 8730
rect 34431 8678 34443 8730
rect 34495 8678 34507 8730
rect 34559 8678 38824 8730
rect 1104 8656 38824 8678
rect 2041 8619 2099 8625
rect 2041 8585 2053 8619
rect 2087 8616 2099 8619
rect 2087 8588 3832 8616
rect 2087 8585 2099 8588
rect 2041 8579 2099 8585
rect 1578 8548 1584 8560
rect 1539 8520 1584 8548
rect 1578 8508 1584 8520
rect 1636 8508 1642 8560
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 2056 8412 2084 8579
rect 3804 8548 3832 8588
rect 3878 8576 3884 8628
rect 3936 8616 3942 8628
rect 3973 8619 4031 8625
rect 3973 8616 3985 8619
rect 3936 8588 3985 8616
rect 3936 8576 3942 8588
rect 3973 8585 3985 8588
rect 4019 8585 4031 8619
rect 4614 8616 4620 8628
rect 4575 8588 4620 8616
rect 3973 8579 4031 8585
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 5074 8616 5080 8628
rect 4987 8588 5080 8616
rect 5074 8576 5080 8588
rect 5132 8616 5138 8628
rect 6178 8616 6184 8628
rect 5132 8588 6184 8616
rect 5132 8576 5138 8588
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 6273 8619 6331 8625
rect 6273 8585 6285 8619
rect 6319 8616 6331 8619
rect 6546 8616 6552 8628
rect 6319 8588 6552 8616
rect 6319 8585 6331 8588
rect 6273 8579 6331 8585
rect 5258 8548 5264 8560
rect 3804 8520 5120 8548
rect 5219 8520 5264 8548
rect 5092 8480 5120 8520
rect 5258 8508 5264 8520
rect 5316 8508 5322 8560
rect 6288 8548 6316 8579
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 7006 8616 7012 8628
rect 6967 8588 7012 8616
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 8389 8619 8447 8625
rect 8389 8616 8401 8619
rect 8168 8588 8401 8616
rect 8168 8576 8174 8588
rect 8389 8585 8401 8588
rect 8435 8585 8447 8619
rect 10962 8616 10968 8628
rect 10923 8588 10968 8616
rect 8389 8579 8447 8585
rect 5368 8520 6316 8548
rect 5368 8480 5396 8520
rect 7282 8508 7288 8560
rect 7340 8548 7346 8560
rect 7929 8551 7987 8557
rect 7929 8548 7941 8551
rect 7340 8520 7941 8548
rect 7340 8508 7346 8520
rect 7929 8517 7941 8520
rect 7975 8517 7987 8551
rect 7929 8511 7987 8517
rect 5718 8480 5724 8492
rect 5092 8452 5396 8480
rect 5679 8452 5724 8480
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8480 6699 8483
rect 7469 8483 7527 8489
rect 7469 8480 7481 8483
rect 6687 8452 7481 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 7469 8449 7481 8452
rect 7515 8480 7527 8483
rect 8018 8480 8024 8492
rect 7515 8452 8024 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 8018 8440 8024 8452
rect 8076 8440 8082 8492
rect 8404 8480 8432 8579
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11238 8576 11244 8628
rect 11296 8616 11302 8628
rect 11425 8619 11483 8625
rect 11425 8616 11437 8619
rect 11296 8588 11437 8616
rect 11296 8576 11302 8588
rect 11425 8585 11437 8588
rect 11471 8616 11483 8619
rect 11514 8616 11520 8628
rect 11471 8588 11520 8616
rect 11471 8585 11483 8588
rect 11425 8579 11483 8585
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 12066 8576 12072 8628
rect 12124 8616 12130 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 12124 8588 12173 8616
rect 12124 8576 12130 8588
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 12161 8579 12219 8585
rect 13909 8619 13967 8625
rect 13909 8585 13921 8619
rect 13955 8616 13967 8619
rect 14918 8616 14924 8628
rect 13955 8588 14924 8616
rect 13955 8585 13967 8588
rect 13909 8579 13967 8585
rect 14918 8576 14924 8588
rect 14976 8576 14982 8628
rect 16758 8616 16764 8628
rect 16719 8588 16764 8616
rect 16758 8576 16764 8588
rect 16816 8576 16822 8628
rect 18598 8576 18604 8628
rect 18656 8616 18662 8628
rect 18693 8619 18751 8625
rect 18693 8616 18705 8619
rect 18656 8588 18705 8616
rect 18656 8576 18662 8588
rect 18693 8585 18705 8588
rect 18739 8585 18751 8619
rect 19058 8616 19064 8628
rect 19019 8588 19064 8616
rect 18693 8579 18751 8585
rect 19058 8576 19064 8588
rect 19116 8576 19122 8628
rect 19334 8616 19340 8628
rect 19295 8588 19340 8616
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 23477 8619 23535 8625
rect 23477 8585 23489 8619
rect 23523 8616 23535 8619
rect 24302 8616 24308 8628
rect 23523 8588 24308 8616
rect 23523 8585 23535 8588
rect 23477 8579 23535 8585
rect 24302 8576 24308 8588
rect 24360 8576 24366 8628
rect 24578 8576 24584 8628
rect 24636 8616 24642 8628
rect 25130 8616 25136 8628
rect 24636 8588 25136 8616
rect 24636 8576 24642 8588
rect 25130 8576 25136 8588
rect 25188 8616 25194 8628
rect 25225 8619 25283 8625
rect 25225 8616 25237 8619
rect 25188 8588 25237 8616
rect 25188 8576 25194 8588
rect 25225 8585 25237 8588
rect 25271 8585 25283 8619
rect 26142 8616 26148 8628
rect 26103 8588 26148 8616
rect 25225 8579 25283 8585
rect 26142 8576 26148 8588
rect 26200 8576 26206 8628
rect 27709 8619 27767 8625
rect 27709 8585 27721 8619
rect 27755 8616 27767 8619
rect 28902 8616 28908 8628
rect 27755 8588 28908 8616
rect 27755 8585 27767 8588
rect 27709 8579 27767 8585
rect 28902 8576 28908 8588
rect 28960 8576 28966 8628
rect 29546 8576 29552 8628
rect 29604 8616 29610 8628
rect 30285 8619 30343 8625
rect 30285 8616 30297 8619
rect 29604 8588 30297 8616
rect 29604 8576 29610 8588
rect 30285 8585 30297 8588
rect 30331 8585 30343 8619
rect 30285 8579 30343 8585
rect 33689 8619 33747 8625
rect 33689 8585 33701 8619
rect 33735 8616 33747 8619
rect 33870 8616 33876 8628
rect 33735 8588 33876 8616
rect 33735 8585 33747 8588
rect 33689 8579 33747 8585
rect 9950 8548 9956 8560
rect 9911 8520 9956 8548
rect 9950 8508 9956 8520
rect 10008 8548 10014 8560
rect 11698 8548 11704 8560
rect 10008 8520 11704 8548
rect 10008 8508 10014 8520
rect 11698 8508 11704 8520
rect 11756 8548 11762 8560
rect 11793 8551 11851 8557
rect 11793 8548 11805 8551
rect 11756 8520 11805 8548
rect 11756 8508 11762 8520
rect 11793 8517 11805 8520
rect 11839 8517 11851 8551
rect 28718 8548 28724 8560
rect 28679 8520 28724 8548
rect 11793 8511 11851 8517
rect 28718 8508 28724 8520
rect 28776 8508 28782 8560
rect 29362 8548 29368 8560
rect 29323 8520 29368 8548
rect 29362 8508 29368 8520
rect 29420 8508 29426 8560
rect 30300 8548 30328 8579
rect 33870 8576 33876 8588
rect 33928 8576 33934 8628
rect 35894 8616 35900 8628
rect 35855 8588 35900 8616
rect 35894 8576 35900 8588
rect 35952 8576 35958 8628
rect 30300 8520 32260 8548
rect 8573 8483 8631 8489
rect 8573 8480 8585 8483
rect 8404 8452 8585 8480
rect 8573 8449 8585 8452
rect 8619 8449 8631 8483
rect 8573 8443 8631 8449
rect 13357 8483 13415 8489
rect 13357 8449 13369 8483
rect 13403 8480 13415 8483
rect 14458 8480 14464 8492
rect 13403 8452 14464 8480
rect 13403 8449 13415 8452
rect 13357 8443 13415 8449
rect 2593 8415 2651 8421
rect 2593 8412 2605 8415
rect 1443 8384 2084 8412
rect 2424 8384 2605 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 1854 8236 1860 8288
rect 1912 8276 1918 8288
rect 2424 8285 2452 8384
rect 2593 8381 2605 8384
rect 2639 8412 2651 8415
rect 2682 8412 2688 8424
rect 2639 8384 2688 8412
rect 2639 8381 2651 8384
rect 2593 8375 2651 8381
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 7558 8412 7564 8424
rect 6788 8384 7564 8412
rect 6788 8372 6794 8384
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 8588 8412 8616 8443
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 15102 8440 15108 8492
rect 15160 8480 15166 8492
rect 15381 8483 15439 8489
rect 15381 8480 15393 8483
rect 15160 8452 15393 8480
rect 15160 8440 15166 8452
rect 15381 8449 15393 8452
rect 15427 8449 15439 8483
rect 15381 8443 15439 8449
rect 19518 8440 19524 8492
rect 19576 8480 19582 8492
rect 19889 8483 19947 8489
rect 19889 8480 19901 8483
rect 19576 8452 19901 8480
rect 19576 8440 19582 8452
rect 19889 8449 19901 8452
rect 19935 8480 19947 8483
rect 19978 8480 19984 8492
rect 19935 8452 19984 8480
rect 19935 8449 19947 8452
rect 19889 8443 19947 8449
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 24210 8440 24216 8492
rect 24268 8480 24274 8492
rect 24857 8483 24915 8489
rect 24857 8480 24869 8483
rect 24268 8452 24869 8480
rect 24268 8440 24274 8452
rect 24857 8449 24869 8452
rect 24903 8449 24915 8483
rect 26510 8480 26516 8492
rect 26471 8452 26516 8480
rect 24857 8443 24915 8449
rect 26510 8440 26516 8452
rect 26568 8440 26574 8492
rect 26602 8440 26608 8492
rect 26660 8480 26666 8492
rect 26697 8483 26755 8489
rect 26697 8480 26709 8483
rect 26660 8452 26709 8480
rect 26660 8440 26666 8452
rect 26697 8449 26709 8452
rect 26743 8449 26755 8483
rect 28166 8480 28172 8492
rect 28079 8452 28172 8480
rect 26697 8443 26755 8449
rect 28166 8440 28172 8452
rect 28224 8480 28230 8492
rect 28810 8480 28816 8492
rect 28224 8452 28816 8480
rect 28224 8440 28230 8452
rect 28810 8440 28816 8452
rect 28868 8440 28874 8492
rect 29089 8483 29147 8489
rect 29089 8449 29101 8483
rect 29135 8480 29147 8483
rect 29178 8480 29184 8492
rect 29135 8452 29184 8480
rect 29135 8449 29147 8452
rect 29089 8443 29147 8449
rect 29178 8440 29184 8452
rect 29236 8480 29242 8492
rect 29917 8483 29975 8489
rect 29917 8480 29929 8483
rect 29236 8452 29929 8480
rect 29236 8440 29242 8452
rect 29917 8449 29929 8452
rect 29963 8449 29975 8483
rect 31294 8480 31300 8492
rect 31255 8452 31300 8480
rect 29917 8443 29975 8449
rect 31294 8440 31300 8452
rect 31352 8440 31358 8492
rect 11238 8412 11244 8424
rect 8588 8384 11244 8412
rect 11238 8372 11244 8384
rect 11296 8372 11302 8424
rect 13725 8415 13783 8421
rect 13725 8381 13737 8415
rect 13771 8412 13783 8415
rect 13771 8384 14412 8412
rect 13771 8381 13783 8384
rect 13725 8375 13783 8381
rect 2860 8347 2918 8353
rect 2860 8313 2872 8347
rect 2906 8344 2918 8347
rect 3142 8344 3148 8356
rect 2906 8316 3148 8344
rect 2906 8313 2918 8316
rect 2860 8307 2918 8313
rect 3142 8304 3148 8316
rect 3200 8304 3206 8356
rect 5442 8304 5448 8356
rect 5500 8344 5506 8356
rect 5718 8344 5724 8356
rect 5500 8316 5724 8344
rect 5500 8304 5506 8316
rect 5718 8304 5724 8316
rect 5776 8304 5782 8356
rect 5813 8347 5871 8353
rect 5813 8313 5825 8347
rect 5859 8344 5871 8347
rect 6362 8344 6368 8356
rect 5859 8316 6368 8344
rect 5859 8313 5871 8316
rect 5813 8307 5871 8313
rect 2409 8279 2467 8285
rect 2409 8276 2421 8279
rect 1912 8248 2421 8276
rect 1912 8236 1918 8248
rect 2409 8245 2421 8248
rect 2455 8245 2467 8279
rect 2409 8239 2467 8245
rect 5166 8236 5172 8288
rect 5224 8276 5230 8288
rect 5828 8276 5856 8307
rect 6362 8304 6368 8316
rect 6420 8304 6426 8356
rect 7576 8344 7604 8372
rect 8818 8347 8876 8353
rect 8818 8344 8830 8347
rect 7576 8316 8830 8344
rect 8818 8313 8830 8316
rect 8864 8344 8876 8347
rect 9398 8344 9404 8356
rect 8864 8316 9404 8344
rect 8864 8313 8876 8316
rect 8818 8307 8876 8313
rect 9398 8304 9404 8316
rect 9456 8304 9462 8356
rect 10502 8344 10508 8356
rect 10463 8316 10508 8344
rect 10502 8304 10508 8316
rect 10560 8304 10566 8356
rect 14182 8344 14188 8356
rect 14143 8316 14188 8344
rect 14182 8304 14188 8316
rect 14240 8304 14246 8356
rect 14384 8353 14412 8384
rect 15194 8372 15200 8424
rect 15252 8372 15258 8424
rect 19058 8372 19064 8424
rect 19116 8412 19122 8424
rect 20809 8415 20867 8421
rect 19116 8384 19840 8412
rect 19116 8372 19122 8384
rect 14369 8347 14427 8353
rect 14369 8313 14381 8347
rect 14415 8344 14427 8347
rect 14642 8344 14648 8356
rect 14415 8316 14648 8344
rect 14415 8313 14427 8316
rect 14369 8307 14427 8313
rect 14642 8304 14648 8316
rect 14700 8304 14706 8356
rect 14921 8347 14979 8353
rect 14921 8313 14933 8347
rect 14967 8344 14979 8347
rect 15212 8344 15240 8372
rect 15654 8353 15660 8356
rect 15648 8344 15660 8353
rect 14967 8316 15660 8344
rect 14967 8313 14979 8316
rect 14921 8307 14979 8313
rect 15648 8307 15660 8316
rect 15654 8304 15660 8307
rect 15712 8304 15718 8356
rect 18046 8344 18052 8356
rect 18007 8316 18052 8344
rect 18046 8304 18052 8316
rect 18104 8304 18110 8356
rect 18598 8304 18604 8356
rect 18656 8344 18662 8356
rect 19812 8353 19840 8384
rect 20809 8381 20821 8415
rect 20855 8412 20867 8415
rect 20898 8412 20904 8424
rect 20855 8384 20904 8412
rect 20855 8381 20867 8384
rect 20809 8375 20867 8381
rect 20898 8372 20904 8384
rect 20956 8372 20962 8424
rect 26142 8372 26148 8424
rect 26200 8412 26206 8424
rect 26528 8412 26556 8440
rect 26200 8384 26556 8412
rect 27157 8415 27215 8421
rect 26200 8372 26206 8384
rect 27157 8381 27169 8415
rect 27203 8412 27215 8415
rect 27246 8412 27252 8424
rect 27203 8384 27252 8412
rect 27203 8381 27215 8384
rect 27157 8375 27215 8381
rect 27246 8372 27252 8384
rect 27304 8412 27310 8424
rect 27525 8415 27583 8421
rect 27525 8412 27537 8415
rect 27304 8384 27537 8412
rect 27304 8372 27310 8384
rect 27525 8381 27537 8384
rect 27571 8412 27583 8415
rect 27571 8384 28304 8412
rect 27571 8381 27583 8384
rect 27525 8375 27583 8381
rect 28276 8356 28304 8384
rect 28902 8372 28908 8424
rect 28960 8412 28966 8424
rect 32232 8421 32260 8520
rect 34146 8508 34152 8560
rect 34204 8548 34210 8560
rect 34977 8551 35035 8557
rect 34977 8548 34989 8551
rect 34204 8520 34989 8548
rect 34204 8508 34210 8520
rect 34977 8517 34989 8520
rect 35023 8517 35035 8551
rect 34977 8511 35035 8517
rect 34054 8440 34060 8492
rect 34112 8480 34118 8492
rect 35437 8483 35495 8489
rect 35437 8480 35449 8483
rect 34112 8452 35449 8480
rect 34112 8440 34118 8452
rect 35437 8449 35449 8452
rect 35483 8480 35495 8483
rect 35802 8480 35808 8492
rect 35483 8452 35808 8480
rect 35483 8449 35495 8452
rect 35437 8443 35495 8449
rect 35802 8440 35808 8452
rect 35860 8440 35866 8492
rect 36725 8483 36783 8489
rect 36725 8449 36737 8483
rect 36771 8480 36783 8483
rect 36814 8480 36820 8492
rect 36771 8452 36820 8480
rect 36771 8449 36783 8452
rect 36725 8443 36783 8449
rect 36814 8440 36820 8452
rect 36872 8440 36878 8492
rect 31021 8415 31079 8421
rect 31021 8412 31033 8415
rect 28960 8384 29868 8412
rect 28960 8372 28966 8384
rect 19613 8347 19671 8353
rect 19613 8344 19625 8347
rect 18656 8316 19625 8344
rect 18656 8304 18662 8316
rect 19613 8313 19625 8316
rect 19659 8313 19671 8347
rect 19613 8307 19671 8313
rect 19797 8347 19855 8353
rect 19797 8313 19809 8347
rect 19843 8313 19855 8347
rect 20346 8344 20352 8356
rect 20259 8316 20352 8344
rect 19797 8307 19855 8313
rect 20346 8304 20352 8316
rect 20404 8344 20410 8356
rect 21076 8347 21134 8353
rect 21076 8344 21088 8347
rect 20404 8316 21088 8344
rect 20404 8304 20410 8316
rect 21076 8313 21088 8316
rect 21122 8344 21134 8347
rect 21450 8344 21456 8356
rect 21122 8316 21456 8344
rect 21122 8313 21134 8316
rect 21076 8307 21134 8313
rect 21450 8304 21456 8316
rect 21508 8304 21514 8356
rect 23934 8304 23940 8356
rect 23992 8344 23998 8356
rect 24029 8347 24087 8353
rect 24029 8344 24041 8347
rect 23992 8316 24041 8344
rect 23992 8304 23998 8316
rect 24029 8313 24041 8316
rect 24075 8344 24087 8347
rect 24581 8347 24639 8353
rect 24581 8344 24593 8347
rect 24075 8316 24593 8344
rect 24075 8313 24087 8316
rect 24029 8307 24087 8313
rect 24581 8313 24593 8316
rect 24627 8344 24639 8347
rect 25961 8347 26019 8353
rect 24627 8316 25912 8344
rect 24627 8313 24639 8316
rect 24581 8307 24639 8313
rect 7466 8276 7472 8288
rect 5224 8248 5856 8276
rect 7427 8248 7472 8276
rect 5224 8236 5230 8248
rect 7466 8236 7472 8248
rect 7524 8236 7530 8288
rect 12713 8279 12771 8285
rect 12713 8245 12725 8279
rect 12759 8276 12771 8279
rect 12894 8276 12900 8288
rect 12759 8248 12900 8276
rect 12759 8245 12771 8248
rect 12713 8239 12771 8245
rect 12894 8236 12900 8248
rect 12952 8236 12958 8288
rect 15102 8236 15108 8288
rect 15160 8276 15166 8288
rect 15197 8279 15255 8285
rect 15197 8276 15209 8279
rect 15160 8248 15209 8276
rect 15160 8236 15166 8248
rect 15197 8245 15209 8248
rect 15243 8245 15255 8279
rect 17310 8276 17316 8288
rect 17271 8248 17316 8276
rect 15197 8239 15255 8245
rect 17310 8236 17316 8248
rect 17368 8236 17374 8288
rect 20717 8279 20775 8285
rect 20717 8245 20729 8279
rect 20763 8276 20775 8279
rect 20898 8276 20904 8288
rect 20763 8248 20904 8276
rect 20763 8245 20775 8248
rect 20717 8239 20775 8245
rect 20898 8236 20904 8248
rect 20956 8236 20962 8288
rect 22186 8276 22192 8288
rect 22147 8248 22192 8276
rect 22186 8236 22192 8248
rect 22244 8236 22250 8288
rect 22922 8276 22928 8288
rect 22883 8248 22928 8276
rect 22922 8236 22928 8248
rect 22980 8236 22986 8288
rect 23474 8236 23480 8288
rect 23532 8276 23538 8288
rect 24302 8276 24308 8288
rect 23532 8248 24308 8276
rect 23532 8236 23538 8248
rect 24302 8236 24308 8248
rect 24360 8276 24366 8288
rect 24765 8279 24823 8285
rect 24765 8276 24777 8279
rect 24360 8248 24777 8276
rect 24360 8236 24366 8248
rect 24765 8245 24777 8248
rect 24811 8245 24823 8279
rect 25884 8276 25912 8316
rect 25961 8313 25973 8347
rect 26007 8344 26019 8347
rect 26418 8344 26424 8356
rect 26007 8316 26424 8344
rect 26007 8313 26019 8316
rect 25961 8307 26019 8313
rect 26418 8304 26424 8316
rect 26476 8344 26482 8356
rect 26605 8347 26663 8353
rect 26605 8344 26617 8347
rect 26476 8316 26617 8344
rect 26476 8304 26482 8316
rect 26605 8313 26617 8316
rect 26651 8344 26663 8347
rect 27062 8344 27068 8356
rect 26651 8316 27068 8344
rect 26651 8313 26663 8316
rect 26605 8307 26663 8313
rect 27062 8304 27068 8316
rect 27120 8304 27126 8356
rect 28074 8304 28080 8356
rect 28132 8344 28138 8356
rect 28169 8347 28227 8353
rect 28169 8344 28181 8347
rect 28132 8316 28181 8344
rect 28132 8304 28138 8316
rect 28169 8313 28181 8316
rect 28215 8313 28227 8347
rect 28169 8307 28227 8313
rect 28258 8304 28264 8356
rect 28316 8344 28322 8356
rect 28316 8316 28361 8344
rect 28316 8304 28322 8316
rect 29546 8304 29552 8356
rect 29604 8344 29610 8356
rect 29840 8353 29868 8384
rect 30944 8384 31033 8412
rect 29641 8347 29699 8353
rect 29641 8344 29653 8347
rect 29604 8316 29653 8344
rect 29604 8304 29610 8316
rect 29641 8313 29653 8316
rect 29687 8313 29699 8347
rect 29641 8307 29699 8313
rect 29825 8347 29883 8353
rect 29825 8313 29837 8347
rect 29871 8313 29883 8347
rect 29825 8307 29883 8313
rect 30944 8288 30972 8384
rect 31021 8381 31033 8384
rect 31067 8381 31079 8415
rect 31021 8375 31079 8381
rect 32217 8415 32275 8421
rect 32217 8381 32229 8415
rect 32263 8412 32275 8415
rect 32309 8415 32367 8421
rect 32309 8412 32321 8415
rect 32263 8384 32321 8412
rect 32263 8381 32275 8384
rect 32217 8375 32275 8381
rect 32309 8381 32321 8384
rect 32355 8412 32367 8415
rect 33042 8412 33048 8424
rect 32355 8384 33048 8412
rect 32355 8381 32367 8384
rect 32309 8375 32367 8381
rect 33042 8372 33048 8384
rect 33100 8412 33106 8424
rect 33962 8412 33968 8424
rect 33100 8384 33968 8412
rect 33100 8372 33106 8384
rect 33962 8372 33968 8384
rect 34020 8412 34026 8424
rect 34333 8415 34391 8421
rect 34333 8412 34345 8415
rect 34020 8384 34345 8412
rect 34020 8372 34026 8384
rect 34333 8381 34345 8384
rect 34379 8412 34391 8415
rect 34422 8412 34428 8424
rect 34379 8384 34428 8412
rect 34379 8381 34391 8384
rect 34333 8375 34391 8381
rect 34422 8372 34428 8384
rect 34480 8372 34486 8424
rect 36265 8415 36323 8421
rect 36265 8412 36277 8415
rect 35452 8384 36277 8412
rect 35452 8356 35480 8384
rect 36265 8381 36277 8384
rect 36311 8381 36323 8415
rect 36446 8412 36452 8424
rect 36407 8384 36452 8412
rect 36265 8375 36323 8381
rect 36446 8372 36452 8384
rect 36504 8412 36510 8424
rect 37185 8415 37243 8421
rect 37185 8412 37197 8415
rect 36504 8384 37197 8412
rect 36504 8372 36510 8384
rect 37185 8381 37197 8384
rect 37231 8381 37243 8415
rect 37185 8375 37243 8381
rect 31846 8344 31852 8356
rect 31807 8316 31852 8344
rect 31846 8304 31852 8316
rect 31904 8304 31910 8356
rect 32582 8353 32588 8356
rect 32576 8344 32588 8353
rect 32543 8316 32588 8344
rect 32576 8307 32588 8316
rect 32582 8304 32588 8307
rect 32640 8304 32646 8356
rect 33226 8304 33232 8356
rect 33284 8344 33290 8356
rect 34701 8347 34759 8353
rect 34701 8344 34713 8347
rect 33284 8316 34713 8344
rect 33284 8304 33290 8316
rect 34701 8313 34713 8316
rect 34747 8344 34759 8347
rect 35434 8344 35440 8356
rect 34747 8316 35296 8344
rect 35347 8316 35440 8344
rect 34747 8313 34759 8316
rect 34701 8307 34759 8313
rect 26694 8276 26700 8288
rect 25884 8248 26700 8276
rect 24765 8239 24823 8245
rect 26694 8236 26700 8248
rect 26752 8276 26758 8288
rect 28350 8276 28356 8288
rect 26752 8248 28356 8276
rect 26752 8236 26758 8248
rect 28350 8236 28356 8248
rect 28408 8236 28414 8288
rect 30926 8276 30932 8288
rect 30887 8248 30932 8276
rect 30926 8236 30932 8248
rect 30984 8236 30990 8288
rect 35268 8276 35296 8316
rect 35434 8304 35440 8316
rect 35492 8304 35498 8356
rect 35529 8347 35587 8353
rect 35529 8313 35541 8347
rect 35575 8313 35587 8347
rect 35529 8307 35587 8313
rect 35544 8276 35572 8307
rect 35268 8248 35572 8276
rect 1104 8186 38824 8208
rect 1104 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 27648 8186
rect 27700 8134 27712 8186
rect 27764 8134 27776 8186
rect 27828 8134 27840 8186
rect 27892 8134 38824 8186
rect 1104 8112 38824 8134
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 2832 8044 3801 8072
rect 2832 8032 2838 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 4246 8072 4252 8084
rect 4207 8044 4252 8072
rect 3789 8035 3847 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4893 8075 4951 8081
rect 4893 8041 4905 8075
rect 4939 8072 4951 8075
rect 5442 8072 5448 8084
rect 4939 8044 5448 8072
rect 4939 8041 4951 8044
rect 4893 8035 4951 8041
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 6086 8032 6092 8084
rect 6144 8072 6150 8084
rect 6365 8075 6423 8081
rect 6365 8072 6377 8075
rect 6144 8044 6377 8072
rect 6144 8032 6150 8044
rect 6365 8041 6377 8044
rect 6411 8072 6423 8075
rect 8021 8075 8079 8081
rect 6411 8044 7880 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 2958 8004 2964 8016
rect 2919 7976 2964 8004
rect 2958 7964 2964 7976
rect 3016 7964 3022 8016
rect 5166 8004 5172 8016
rect 5127 7976 5172 8004
rect 5166 7964 5172 7976
rect 5224 7964 5230 8016
rect 5905 8007 5963 8013
rect 5905 7973 5917 8007
rect 5951 7973 5963 8007
rect 6730 8004 6736 8016
rect 6691 7976 6736 8004
rect 5905 7967 5963 7973
rect 2406 7896 2412 7948
rect 2464 7936 2470 7948
rect 3421 7939 3479 7945
rect 3421 7936 3433 7939
rect 2464 7908 3433 7936
rect 2464 7896 2470 7908
rect 3421 7905 3433 7908
rect 3467 7905 3479 7939
rect 4062 7936 4068 7948
rect 4023 7908 4068 7936
rect 3421 7899 3479 7905
rect 4062 7896 4068 7908
rect 4120 7896 4126 7948
rect 5920 7936 5948 7967
rect 6730 7964 6736 7976
rect 6788 7964 6794 8016
rect 7006 7964 7012 8016
rect 7064 8004 7070 8016
rect 7469 8007 7527 8013
rect 7469 8004 7481 8007
rect 7064 7976 7481 8004
rect 7064 7964 7070 7976
rect 7469 7973 7481 7976
rect 7515 8004 7527 8007
rect 7742 8004 7748 8016
rect 7515 7976 7748 8004
rect 7515 7973 7527 7976
rect 7469 7967 7527 7973
rect 7742 7964 7748 7976
rect 7800 7964 7806 8016
rect 7852 8004 7880 8044
rect 8021 8041 8033 8075
rect 8067 8072 8079 8075
rect 8202 8072 8208 8084
rect 8067 8044 8208 8072
rect 8067 8041 8079 8044
rect 8021 8035 8079 8041
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 9398 8072 9404 8084
rect 9359 8044 9404 8072
rect 9398 8032 9404 8044
rect 9456 8032 9462 8084
rect 10226 8072 10232 8084
rect 10187 8044 10232 8072
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 15654 8032 15660 8084
rect 15712 8072 15718 8084
rect 16301 8075 16359 8081
rect 16301 8072 16313 8075
rect 15712 8044 16313 8072
rect 15712 8032 15718 8044
rect 16301 8041 16313 8044
rect 16347 8041 16359 8075
rect 17126 8072 17132 8084
rect 17087 8044 17132 8072
rect 16301 8035 16359 8041
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 18690 8072 18696 8084
rect 18651 8044 18696 8072
rect 18690 8032 18696 8044
rect 18748 8032 18754 8084
rect 19978 8072 19984 8084
rect 19939 8044 19984 8072
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 20714 8032 20720 8084
rect 20772 8072 20778 8084
rect 20901 8075 20959 8081
rect 20901 8072 20913 8075
rect 20772 8044 20913 8072
rect 20772 8032 20778 8044
rect 20901 8041 20913 8044
rect 20947 8041 20959 8075
rect 21450 8072 21456 8084
rect 21411 8044 21456 8072
rect 20901 8035 20959 8041
rect 21450 8032 21456 8044
rect 21508 8032 21514 8084
rect 21634 8032 21640 8084
rect 21692 8072 21698 8084
rect 22097 8075 22155 8081
rect 22097 8072 22109 8075
rect 21692 8044 22109 8072
rect 21692 8032 21698 8044
rect 22097 8041 22109 8044
rect 22143 8041 22155 8075
rect 22097 8035 22155 8041
rect 24673 8075 24731 8081
rect 24673 8041 24685 8075
rect 24719 8072 24731 8075
rect 24762 8072 24768 8084
rect 24719 8044 24768 8072
rect 24719 8041 24731 8044
rect 24673 8035 24731 8041
rect 24762 8032 24768 8044
rect 24820 8032 24826 8084
rect 26142 8072 26148 8084
rect 26103 8044 26148 8072
rect 26142 8032 26148 8044
rect 26200 8032 26206 8084
rect 27985 8075 28043 8081
rect 27985 8041 27997 8075
rect 28031 8072 28043 8075
rect 28166 8072 28172 8084
rect 28031 8044 28172 8072
rect 28031 8041 28043 8044
rect 27985 8035 28043 8041
rect 28166 8032 28172 8044
rect 28224 8032 28230 8084
rect 30650 8072 30656 8084
rect 30611 8044 30656 8072
rect 30650 8032 30656 8044
rect 30708 8032 30714 8084
rect 34882 8072 34888 8084
rect 34843 8044 34888 8072
rect 34882 8032 34888 8044
rect 34940 8032 34946 8084
rect 35066 8032 35072 8084
rect 35124 8072 35130 8084
rect 36446 8072 36452 8084
rect 35124 8044 36452 8072
rect 35124 8032 35130 8044
rect 36446 8032 36452 8044
rect 36504 8032 36510 8084
rect 36630 8032 36636 8084
rect 36688 8072 36694 8084
rect 36817 8075 36875 8081
rect 36817 8072 36829 8075
rect 36688 8044 36829 8072
rect 36688 8032 36694 8044
rect 36817 8041 36829 8044
rect 36863 8041 36875 8075
rect 36817 8035 36875 8041
rect 8481 8007 8539 8013
rect 8481 8004 8493 8007
rect 7852 7976 8493 8004
rect 8481 7973 8493 7976
rect 8527 7973 8539 8007
rect 11762 8007 11820 8013
rect 11762 8004 11774 8007
rect 8481 7967 8539 7973
rect 11256 7976 11774 8004
rect 6914 7936 6920 7948
rect 5920 7908 6920 7936
rect 6914 7896 6920 7908
rect 6972 7936 6978 7948
rect 8297 7939 8355 7945
rect 8297 7936 8309 7939
rect 6972 7908 8309 7936
rect 6972 7896 6978 7908
rect 8297 7905 8309 7908
rect 8343 7905 8355 7939
rect 8297 7899 8355 7905
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7868 1455 7871
rect 2225 7871 2283 7877
rect 2225 7868 2237 7871
rect 1443 7840 2237 7868
rect 1443 7837 1455 7840
rect 1397 7831 1455 7837
rect 2225 7837 2237 7840
rect 2271 7868 2283 7871
rect 2869 7871 2927 7877
rect 2869 7868 2881 7871
rect 2271 7840 2881 7868
rect 2271 7837 2283 7840
rect 2225 7831 2283 7837
rect 2869 7837 2881 7840
rect 2915 7837 2927 7871
rect 3050 7868 3056 7880
rect 3011 7840 3056 7868
rect 2869 7831 2927 7837
rect 3050 7828 3056 7840
rect 3108 7828 3114 7880
rect 5258 7828 5264 7880
rect 5316 7868 5322 7880
rect 5902 7868 5908 7880
rect 5316 7840 5908 7868
rect 5316 7828 5322 7840
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 5997 7871 6055 7877
rect 5997 7837 6009 7871
rect 6043 7868 6055 7871
rect 6178 7868 6184 7880
rect 6043 7840 6184 7868
rect 6043 7837 6055 7840
rect 5997 7831 6055 7837
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7837 7435 7871
rect 7558 7868 7564 7880
rect 7519 7840 7564 7868
rect 7377 7831 7435 7837
rect 5350 7760 5356 7812
rect 5408 7800 5414 7812
rect 5445 7803 5503 7809
rect 5445 7800 5457 7803
rect 5408 7772 5457 7800
rect 5408 7760 5414 7772
rect 5445 7769 5457 7772
rect 5491 7769 5503 7803
rect 5445 7763 5503 7769
rect 7009 7803 7067 7809
rect 7009 7769 7021 7803
rect 7055 7800 7067 7803
rect 7190 7800 7196 7812
rect 7055 7772 7196 7800
rect 7055 7769 7067 7772
rect 7009 7763 7067 7769
rect 7190 7760 7196 7772
rect 7248 7760 7254 7812
rect 7392 7800 7420 7831
rect 7558 7828 7564 7840
rect 7616 7828 7622 7880
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7868 10379 7871
rect 10778 7868 10784 7880
rect 10367 7840 10784 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 7466 7800 7472 7812
rect 7379 7772 7472 7800
rect 7466 7760 7472 7772
rect 7524 7800 7530 7812
rect 7650 7800 7656 7812
rect 7524 7772 7656 7800
rect 7524 7760 7530 7772
rect 7650 7760 7656 7772
rect 7708 7760 7714 7812
rect 10244 7800 10272 7831
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 11256 7800 11284 7976
rect 11762 7973 11774 7976
rect 11808 8004 11820 8007
rect 12158 8004 12164 8016
rect 11808 7976 12164 8004
rect 11808 7973 11820 7976
rect 11762 7967 11820 7973
rect 12158 7964 12164 7976
rect 12216 7964 12222 8016
rect 19705 8007 19763 8013
rect 19705 7973 19717 8007
rect 19751 8004 19763 8007
rect 19794 8004 19800 8016
rect 19751 7976 19800 8004
rect 19751 7973 19763 7976
rect 19705 7967 19763 7973
rect 19794 7964 19800 7976
rect 19852 8004 19858 8016
rect 25038 8004 25044 8016
rect 19852 7976 25044 8004
rect 19852 7964 19858 7976
rect 25038 7964 25044 7976
rect 25096 7964 25102 8016
rect 25314 8004 25320 8016
rect 25275 7976 25320 8004
rect 25314 7964 25320 7976
rect 25372 7964 25378 8016
rect 27065 8007 27123 8013
rect 27065 7973 27077 8007
rect 27111 7973 27123 8007
rect 27065 7967 27123 7973
rect 28988 8007 29046 8013
rect 28988 7973 29000 8007
rect 29034 8004 29046 8007
rect 29086 8004 29092 8016
rect 29034 7976 29092 8004
rect 29034 7973 29046 7976
rect 28988 7967 29046 7973
rect 11514 7936 11520 7948
rect 11475 7908 11520 7936
rect 11514 7896 11520 7908
rect 11572 7896 11578 7948
rect 15657 7939 15715 7945
rect 15657 7905 15669 7939
rect 15703 7936 15715 7939
rect 16393 7939 16451 7945
rect 16393 7936 16405 7939
rect 15703 7908 16405 7936
rect 15703 7905 15715 7908
rect 15657 7899 15715 7905
rect 16393 7905 16405 7908
rect 16439 7936 16451 7939
rect 16758 7936 16764 7948
rect 16439 7908 16764 7936
rect 16439 7905 16451 7908
rect 16393 7899 16451 7905
rect 16758 7896 16764 7908
rect 16816 7896 16822 7948
rect 17586 7945 17592 7948
rect 17580 7936 17592 7945
rect 17547 7908 17592 7936
rect 17580 7899 17592 7908
rect 17586 7896 17592 7899
rect 17644 7896 17650 7948
rect 20717 7939 20775 7945
rect 20717 7905 20729 7939
rect 20763 7936 20775 7939
rect 20806 7936 20812 7948
rect 20763 7908 20812 7936
rect 20763 7905 20775 7908
rect 20717 7899 20775 7905
rect 20806 7896 20812 7908
rect 20864 7896 20870 7948
rect 21821 7939 21879 7945
rect 21821 7905 21833 7939
rect 21867 7936 21879 7939
rect 22186 7936 22192 7948
rect 21867 7908 22192 7936
rect 21867 7905 21879 7908
rect 21821 7899 21879 7905
rect 22186 7896 22192 7908
rect 22244 7936 22250 7948
rect 22548 7939 22606 7945
rect 22548 7936 22560 7939
rect 22244 7908 22560 7936
rect 22244 7896 22250 7908
rect 22548 7905 22560 7908
rect 22594 7936 22606 7939
rect 23474 7936 23480 7948
rect 22594 7908 23480 7936
rect 22594 7905 22606 7908
rect 22548 7899 22606 7905
rect 23474 7896 23480 7908
rect 23532 7896 23538 7948
rect 24946 7896 24952 7948
rect 25004 7936 25010 7948
rect 25133 7939 25191 7945
rect 25133 7936 25145 7939
rect 25004 7908 25145 7936
rect 25004 7896 25010 7908
rect 25133 7905 25145 7908
rect 25179 7905 25191 7939
rect 25133 7899 25191 7905
rect 16298 7868 16304 7880
rect 16259 7840 16304 7868
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 17310 7868 17316 7880
rect 17271 7840 17316 7868
rect 17310 7828 17316 7840
rect 17368 7828 17374 7880
rect 21910 7828 21916 7880
rect 21968 7868 21974 7880
rect 22094 7868 22100 7880
rect 21968 7840 22100 7868
rect 21968 7828 21974 7840
rect 22094 7828 22100 7840
rect 22152 7868 22158 7880
rect 22281 7871 22339 7877
rect 22281 7868 22293 7871
rect 22152 7840 22293 7868
rect 22152 7828 22158 7840
rect 22281 7837 22293 7840
rect 22327 7837 22339 7871
rect 25406 7868 25412 7880
rect 25367 7840 25412 7868
rect 22281 7831 22339 7837
rect 25406 7828 25412 7840
rect 25464 7828 25470 7880
rect 26970 7868 26976 7880
rect 26931 7840 26976 7868
rect 26970 7828 26976 7840
rect 27028 7828 27034 7880
rect 11330 7800 11336 7812
rect 10244 7772 10364 7800
rect 11256 7772 11336 7800
rect 10336 7744 10364 7772
rect 11330 7760 11336 7772
rect 11388 7760 11394 7812
rect 24857 7803 24915 7809
rect 24857 7769 24869 7803
rect 24903 7800 24915 7803
rect 27080 7800 27108 7967
rect 29086 7964 29092 7976
rect 29144 7964 29150 8016
rect 33226 8013 33232 8016
rect 32769 8007 32827 8013
rect 32769 7973 32781 8007
rect 32815 8004 32827 8007
rect 33220 8004 33232 8013
rect 32815 7976 33232 8004
rect 32815 7973 32827 7976
rect 32769 7967 32827 7973
rect 33220 7967 33232 7976
rect 33226 7964 33232 7967
rect 33284 7964 33290 8016
rect 35986 8004 35992 8016
rect 35947 7976 35992 8004
rect 35986 7964 35992 7976
rect 36044 7964 36050 8016
rect 36078 7964 36084 8016
rect 36136 7964 36142 8016
rect 28718 7936 28724 7948
rect 28631 7908 28724 7936
rect 28718 7896 28724 7908
rect 28776 7936 28782 7948
rect 29454 7936 29460 7948
rect 28776 7908 29460 7936
rect 28776 7896 28782 7908
rect 29454 7896 29460 7908
rect 29512 7896 29518 7948
rect 32953 7939 33011 7945
rect 32953 7905 32965 7939
rect 32999 7936 33011 7939
rect 33042 7936 33048 7948
rect 32999 7908 33048 7936
rect 32999 7905 33011 7908
rect 32953 7899 33011 7905
rect 33042 7896 33048 7908
rect 33100 7896 33106 7948
rect 36096 7936 36124 7964
rect 36004 7908 36124 7936
rect 27157 7871 27215 7877
rect 27157 7837 27169 7871
rect 27203 7868 27215 7871
rect 28074 7868 28080 7880
rect 27203 7840 28080 7868
rect 27203 7837 27215 7840
rect 27157 7831 27215 7837
rect 28074 7828 28080 7840
rect 28132 7828 28138 7880
rect 36004 7877 36032 7908
rect 35989 7871 36047 7877
rect 35989 7837 36001 7871
rect 36035 7837 36047 7871
rect 35989 7831 36047 7837
rect 36081 7871 36139 7877
rect 36081 7837 36093 7871
rect 36127 7837 36139 7871
rect 36081 7831 36139 7837
rect 27525 7803 27583 7809
rect 27525 7800 27537 7803
rect 24903 7772 27537 7800
rect 24903 7769 24915 7772
rect 24857 7763 24915 7769
rect 27525 7769 27537 7772
rect 27571 7769 27583 7803
rect 27525 7763 27583 7769
rect 32401 7803 32459 7809
rect 32401 7769 32413 7803
rect 32447 7800 32459 7803
rect 32582 7800 32588 7812
rect 32447 7772 32588 7800
rect 32447 7769 32459 7772
rect 32401 7763 32459 7769
rect 32582 7760 32588 7772
rect 32640 7800 32646 7812
rect 32640 7772 32996 7800
rect 32640 7760 32646 7772
rect 1854 7732 1860 7744
rect 1815 7704 1860 7732
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 2314 7692 2320 7744
rect 2372 7732 2378 7744
rect 2501 7735 2559 7741
rect 2501 7732 2513 7735
rect 2372 7704 2513 7732
rect 2372 7692 2378 7704
rect 2501 7701 2513 7704
rect 2547 7701 2559 7735
rect 9766 7732 9772 7744
rect 9727 7704 9772 7732
rect 2501 7695 2559 7701
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 10318 7692 10324 7744
rect 10376 7692 10382 7744
rect 10781 7735 10839 7741
rect 10781 7701 10793 7735
rect 10827 7732 10839 7735
rect 11146 7732 11152 7744
rect 10827 7704 11152 7732
rect 10827 7701 10839 7704
rect 10781 7695 10839 7701
rect 11146 7692 11152 7704
rect 11204 7692 11210 7744
rect 12894 7732 12900 7744
rect 12855 7704 12900 7732
rect 12894 7692 12900 7704
rect 12952 7692 12958 7744
rect 13909 7735 13967 7741
rect 13909 7701 13921 7735
rect 13955 7732 13967 7735
rect 14182 7732 14188 7744
rect 13955 7704 14188 7732
rect 13955 7701 13967 7704
rect 13909 7695 13967 7701
rect 14182 7692 14188 7704
rect 14240 7732 14246 7744
rect 14734 7732 14740 7744
rect 14240 7704 14740 7732
rect 14240 7692 14246 7704
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 15838 7732 15844 7744
rect 15799 7704 15844 7732
rect 15838 7692 15844 7704
rect 15896 7692 15902 7744
rect 19334 7732 19340 7744
rect 19295 7704 19340 7732
rect 19334 7692 19340 7704
rect 19392 7692 19398 7744
rect 22922 7692 22928 7744
rect 22980 7732 22986 7744
rect 23566 7732 23572 7744
rect 22980 7704 23572 7732
rect 22980 7692 22986 7704
rect 23566 7692 23572 7704
rect 23624 7732 23630 7744
rect 23661 7735 23719 7741
rect 23661 7732 23673 7735
rect 23624 7704 23673 7732
rect 23624 7692 23630 7704
rect 23661 7701 23673 7704
rect 23707 7701 23719 7735
rect 24302 7732 24308 7744
rect 24263 7704 24308 7732
rect 23661 7695 23719 7701
rect 24302 7692 24308 7704
rect 24360 7692 24366 7744
rect 26234 7692 26240 7744
rect 26292 7732 26298 7744
rect 26605 7735 26663 7741
rect 26605 7732 26617 7735
rect 26292 7704 26617 7732
rect 26292 7692 26298 7704
rect 26605 7701 26617 7704
rect 26651 7701 26663 7735
rect 26605 7695 26663 7701
rect 28258 7692 28264 7744
rect 28316 7732 28322 7744
rect 28629 7735 28687 7741
rect 28629 7732 28641 7735
rect 28316 7704 28641 7732
rect 28316 7692 28322 7704
rect 28629 7701 28641 7704
rect 28675 7732 28687 7735
rect 30098 7732 30104 7744
rect 28675 7704 30104 7732
rect 28675 7701 28687 7704
rect 28629 7695 28687 7701
rect 30098 7692 30104 7704
rect 30156 7692 30162 7744
rect 32968 7732 32996 7772
rect 35434 7760 35440 7812
rect 35492 7800 35498 7812
rect 35529 7803 35587 7809
rect 35529 7800 35541 7803
rect 35492 7772 35541 7800
rect 35492 7760 35498 7772
rect 35529 7769 35541 7772
rect 35575 7769 35587 7803
rect 35529 7763 35587 7769
rect 33594 7732 33600 7744
rect 32968 7704 33600 7732
rect 33594 7692 33600 7704
rect 33652 7732 33658 7744
rect 34333 7735 34391 7741
rect 34333 7732 34345 7735
rect 33652 7704 34345 7732
rect 33652 7692 33658 7704
rect 34333 7701 34345 7704
rect 34379 7701 34391 7735
rect 35250 7732 35256 7744
rect 35211 7704 35256 7732
rect 34333 7695 34391 7701
rect 35250 7692 35256 7704
rect 35308 7732 35314 7744
rect 36096 7732 36124 7831
rect 36538 7732 36544 7744
rect 35308 7704 36544 7732
rect 35308 7692 35314 7704
rect 36538 7692 36544 7704
rect 36596 7692 36602 7744
rect 1104 7642 38824 7664
rect 1104 7590 7648 7642
rect 7700 7590 7712 7642
rect 7764 7590 7776 7642
rect 7828 7590 7840 7642
rect 7892 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 34315 7642
rect 34367 7590 34379 7642
rect 34431 7590 34443 7642
rect 34495 7590 34507 7642
rect 34559 7590 38824 7642
rect 1104 7568 38824 7590
rect 3142 7528 3148 7540
rect 3103 7500 3148 7528
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 4157 7531 4215 7537
rect 4157 7528 4169 7531
rect 4120 7500 4169 7528
rect 4120 7488 4126 7500
rect 4157 7497 4169 7500
rect 4203 7528 4215 7531
rect 6178 7528 6184 7540
rect 4203 7500 6040 7528
rect 6139 7500 6184 7528
rect 4203 7497 4215 7500
rect 4157 7491 4215 7497
rect 6012 7460 6040 7500
rect 6178 7488 6184 7500
rect 6236 7488 6242 7540
rect 6914 7488 6920 7540
rect 6972 7528 6978 7540
rect 7101 7531 7159 7537
rect 7101 7528 7113 7531
rect 6972 7500 7113 7528
rect 6972 7488 6978 7500
rect 7101 7497 7113 7500
rect 7147 7528 7159 7531
rect 7466 7528 7472 7540
rect 7147 7500 7472 7528
rect 7147 7497 7159 7500
rect 7101 7491 7159 7497
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 10137 7531 10195 7537
rect 10137 7497 10149 7531
rect 10183 7528 10195 7531
rect 10226 7528 10232 7540
rect 10183 7500 10232 7528
rect 10183 7497 10195 7500
rect 10137 7491 10195 7497
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 13814 7488 13820 7540
rect 13872 7528 13878 7540
rect 15105 7531 15163 7537
rect 15105 7528 15117 7531
rect 13872 7500 15117 7528
rect 13872 7488 13878 7500
rect 15105 7497 15117 7500
rect 15151 7528 15163 7531
rect 16298 7528 16304 7540
rect 15151 7500 16304 7528
rect 15151 7497 15163 7500
rect 15105 7491 15163 7497
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 20806 7488 20812 7540
rect 20864 7528 20870 7540
rect 20901 7531 20959 7537
rect 20901 7528 20913 7531
rect 20864 7500 20913 7528
rect 20864 7488 20870 7500
rect 20901 7497 20913 7500
rect 20947 7497 20959 7531
rect 23474 7528 23480 7540
rect 23387 7500 23480 7528
rect 20901 7491 20959 7497
rect 6641 7463 6699 7469
rect 6641 7460 6653 7463
rect 6012 7432 6653 7460
rect 6641 7429 6653 7432
rect 6687 7460 6699 7463
rect 7006 7460 7012 7472
rect 6687 7432 7012 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 7006 7420 7012 7432
rect 7064 7460 7070 7472
rect 7374 7460 7380 7472
rect 7064 7432 7380 7460
rect 7064 7420 7070 7432
rect 7374 7420 7380 7432
rect 7432 7420 7438 7472
rect 10686 7460 10692 7472
rect 10647 7432 10692 7460
rect 10686 7420 10692 7432
rect 10744 7420 10750 7472
rect 11514 7420 11520 7472
rect 11572 7460 11578 7472
rect 11609 7463 11667 7469
rect 11609 7460 11621 7463
rect 11572 7432 11621 7460
rect 11572 7420 11578 7432
rect 11609 7429 11621 7432
rect 11655 7460 11667 7463
rect 12161 7463 12219 7469
rect 12161 7460 12173 7463
rect 11655 7432 12173 7460
rect 11655 7429 11667 7432
rect 11609 7423 11667 7429
rect 12161 7429 12173 7432
rect 12207 7429 12219 7463
rect 12161 7423 12219 7429
rect 1765 7327 1823 7333
rect 1765 7324 1777 7327
rect 1596 7296 1777 7324
rect 1486 7148 1492 7200
rect 1544 7188 1550 7200
rect 1596 7188 1624 7296
rect 1765 7293 1777 7296
rect 1811 7324 1823 7327
rect 1854 7324 1860 7336
rect 1811 7296 1860 7324
rect 1811 7293 1823 7296
rect 1765 7287 1823 7293
rect 1854 7284 1860 7296
rect 1912 7284 1918 7336
rect 2032 7327 2090 7333
rect 2032 7293 2044 7327
rect 2078 7324 2090 7327
rect 2406 7324 2412 7336
rect 2078 7296 2412 7324
rect 2078 7293 2090 7296
rect 2032 7287 2090 7293
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 4249 7327 4307 7333
rect 4249 7293 4261 7327
rect 4295 7293 4307 7327
rect 4249 7287 4307 7293
rect 1673 7259 1731 7265
rect 1673 7225 1685 7259
rect 1719 7256 1731 7259
rect 2958 7256 2964 7268
rect 1719 7228 2964 7256
rect 1719 7225 1731 7228
rect 1673 7219 1731 7225
rect 2958 7216 2964 7228
rect 3016 7256 3022 7268
rect 3970 7256 3976 7268
rect 3016 7228 3976 7256
rect 3016 7216 3022 7228
rect 3970 7216 3976 7228
rect 4028 7216 4034 7268
rect 3789 7191 3847 7197
rect 3789 7188 3801 7191
rect 1544 7160 3801 7188
rect 1544 7148 1550 7160
rect 3789 7157 3801 7160
rect 3835 7188 3847 7191
rect 3878 7188 3884 7200
rect 3835 7160 3884 7188
rect 3835 7157 3847 7160
rect 3789 7151 3847 7157
rect 3878 7148 3884 7160
rect 3936 7188 3942 7200
rect 4264 7188 4292 7287
rect 6730 7284 6736 7336
rect 6788 7324 6794 7336
rect 7469 7327 7527 7333
rect 7469 7324 7481 7327
rect 6788 7296 7481 7324
rect 6788 7284 6794 7296
rect 7469 7293 7481 7296
rect 7515 7324 7527 7327
rect 8110 7324 8116 7336
rect 7515 7296 8116 7324
rect 7515 7293 7527 7296
rect 7469 7287 7527 7293
rect 8110 7284 8116 7296
rect 8168 7284 8174 7336
rect 10778 7284 10784 7336
rect 10836 7324 10842 7336
rect 11241 7327 11299 7333
rect 11241 7324 11253 7327
rect 10836 7296 11253 7324
rect 10836 7284 10842 7296
rect 11241 7293 11253 7296
rect 11287 7293 11299 7327
rect 12176 7324 12204 7423
rect 15654 7420 15660 7472
rect 15712 7460 15718 7472
rect 15749 7463 15807 7469
rect 15749 7460 15761 7463
rect 15712 7432 15761 7460
rect 15712 7420 15718 7432
rect 15749 7429 15761 7432
rect 15795 7429 15807 7463
rect 16206 7460 16212 7472
rect 16167 7432 16212 7460
rect 15749 7423 15807 7429
rect 16206 7420 16212 7432
rect 16264 7420 16270 7472
rect 17129 7463 17187 7469
rect 17129 7460 17141 7463
rect 16592 7432 17141 7460
rect 16592 7404 16620 7432
rect 17129 7429 17141 7432
rect 17175 7460 17187 7463
rect 17218 7460 17224 7472
rect 17175 7432 17224 7460
rect 17175 7429 17187 7432
rect 17129 7423 17187 7429
rect 17218 7420 17224 7432
rect 17276 7420 17282 7472
rect 19610 7460 19616 7472
rect 19571 7432 19616 7460
rect 19610 7420 19616 7432
rect 19668 7420 19674 7472
rect 16574 7392 16580 7404
rect 16535 7364 16580 7392
rect 16574 7352 16580 7364
rect 16632 7352 16638 7404
rect 16758 7392 16764 7404
rect 16719 7364 16764 7392
rect 16758 7352 16764 7364
rect 16816 7352 16822 7404
rect 19426 7392 19432 7404
rect 19339 7364 19432 7392
rect 19426 7352 19432 7364
rect 19484 7392 19490 7404
rect 20073 7395 20131 7401
rect 20073 7392 20085 7395
rect 19484 7364 20085 7392
rect 19484 7352 19490 7364
rect 20073 7361 20085 7364
rect 20119 7392 20131 7395
rect 20622 7392 20628 7404
rect 20119 7364 20628 7392
rect 20119 7361 20131 7364
rect 20073 7355 20131 7361
rect 20622 7352 20628 7364
rect 20680 7352 20686 7404
rect 20916 7392 20944 7491
rect 23474 7488 23480 7500
rect 23532 7528 23538 7540
rect 24578 7528 24584 7540
rect 23532 7500 24584 7528
rect 23532 7488 23538 7500
rect 24578 7488 24584 7500
rect 24636 7488 24642 7540
rect 25958 7528 25964 7540
rect 25871 7500 25964 7528
rect 25958 7488 25964 7500
rect 26016 7528 26022 7540
rect 28074 7528 28080 7540
rect 26016 7500 28080 7528
rect 26016 7488 26022 7500
rect 28074 7488 28080 7500
rect 28132 7488 28138 7540
rect 28718 7528 28724 7540
rect 28679 7500 28724 7528
rect 28718 7488 28724 7500
rect 28776 7528 28782 7540
rect 28997 7531 29055 7537
rect 28997 7528 29009 7531
rect 28776 7500 29009 7528
rect 28776 7488 28782 7500
rect 28997 7497 29009 7500
rect 29043 7497 29055 7531
rect 28997 7491 29055 7497
rect 32217 7531 32275 7537
rect 32217 7497 32229 7531
rect 32263 7528 32275 7531
rect 33042 7528 33048 7540
rect 32263 7500 33048 7528
rect 32263 7497 32275 7500
rect 32217 7491 32275 7497
rect 27154 7460 27160 7472
rect 27115 7432 27160 7460
rect 27154 7420 27160 7432
rect 27212 7420 27218 7472
rect 29012 7404 29040 7491
rect 32324 7404 32352 7500
rect 33042 7488 33048 7500
rect 33100 7488 33106 7540
rect 33226 7488 33232 7540
rect 33284 7528 33290 7540
rect 33689 7531 33747 7537
rect 33689 7528 33701 7531
rect 33284 7500 33701 7528
rect 33284 7488 33290 7500
rect 33689 7497 33701 7500
rect 33735 7528 33747 7531
rect 33778 7528 33784 7540
rect 33735 7500 33784 7528
rect 33735 7497 33747 7500
rect 33689 7491 33747 7497
rect 33778 7488 33784 7500
rect 33836 7488 33842 7540
rect 35894 7488 35900 7540
rect 35952 7528 35958 7540
rect 36541 7531 36599 7537
rect 36541 7528 36553 7531
rect 35952 7500 36553 7528
rect 35952 7488 35958 7500
rect 36541 7497 36553 7500
rect 36587 7497 36599 7531
rect 36541 7491 36599 7497
rect 34974 7460 34980 7472
rect 34935 7432 34980 7460
rect 34974 7420 34980 7432
rect 35032 7420 35038 7472
rect 35989 7463 36047 7469
rect 35989 7429 36001 7463
rect 36035 7460 36047 7463
rect 36078 7460 36084 7472
rect 36035 7432 36084 7460
rect 36035 7429 36047 7432
rect 35989 7423 36047 7429
rect 36078 7420 36084 7432
rect 36136 7420 36142 7472
rect 21082 7392 21088 7404
rect 20916 7364 21088 7392
rect 21082 7352 21088 7364
rect 21140 7352 21146 7404
rect 28994 7392 29000 7404
rect 28907 7364 29000 7392
rect 28994 7352 29000 7364
rect 29052 7392 29058 7404
rect 29273 7395 29331 7401
rect 29273 7392 29285 7395
rect 29052 7364 29285 7392
rect 29052 7352 29058 7364
rect 29273 7361 29285 7364
rect 29319 7361 29331 7395
rect 32306 7392 32312 7404
rect 32219 7364 32312 7392
rect 29273 7355 29331 7361
rect 32306 7352 32312 7364
rect 32364 7352 32370 7404
rect 36538 7352 36544 7404
rect 36596 7392 36602 7404
rect 37093 7395 37151 7401
rect 37093 7392 37105 7395
rect 36596 7364 37105 7392
rect 36596 7352 36602 7364
rect 37093 7361 37105 7364
rect 37139 7361 37151 7395
rect 37093 7355 37151 7361
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 12176 7296 12449 7324
rect 11241 7287 11299 7293
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 15470 7324 15476 7336
rect 15383 7296 15476 7324
rect 12437 7287 12495 7293
rect 4516 7259 4574 7265
rect 4516 7225 4528 7259
rect 4562 7256 4574 7259
rect 4706 7256 4712 7268
rect 4562 7228 4712 7256
rect 4562 7225 4574 7228
rect 4516 7219 4574 7225
rect 4706 7216 4712 7228
rect 4764 7216 4770 7268
rect 7742 7265 7748 7268
rect 7736 7256 7748 7265
rect 7703 7228 7748 7256
rect 7736 7219 7748 7228
rect 7742 7216 7748 7219
rect 7800 7216 7806 7268
rect 10962 7256 10968 7268
rect 10875 7228 10968 7256
rect 10962 7216 10968 7228
rect 11020 7216 11026 7268
rect 11146 7256 11152 7268
rect 11107 7228 11152 7256
rect 11146 7216 11152 7228
rect 11204 7216 11210 7268
rect 5626 7188 5632 7200
rect 3936 7160 4292 7188
rect 5587 7160 5632 7188
rect 3936 7148 3942 7160
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 8849 7191 8907 7197
rect 8849 7157 8861 7191
rect 8895 7188 8907 7191
rect 9582 7188 9588 7200
rect 8895 7160 9588 7188
rect 8895 7157 8907 7160
rect 8849 7151 8907 7157
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 9769 7191 9827 7197
rect 9769 7157 9781 7191
rect 9815 7188 9827 7191
rect 10318 7188 10324 7200
rect 9815 7160 10324 7188
rect 9815 7157 9827 7160
rect 9769 7151 9827 7157
rect 10318 7148 10324 7160
rect 10376 7148 10382 7200
rect 10410 7148 10416 7200
rect 10468 7188 10474 7200
rect 10980 7188 11008 7216
rect 10468 7160 11008 7188
rect 11256 7188 11284 7287
rect 15470 7284 15476 7296
rect 15528 7324 15534 7336
rect 19061 7327 19119 7333
rect 15528 7296 16712 7324
rect 15528 7284 15534 7296
rect 16684 7268 16712 7296
rect 19061 7293 19073 7327
rect 19107 7324 19119 7327
rect 24578 7324 24584 7336
rect 19107 7296 20208 7324
rect 24539 7296 24584 7324
rect 19107 7293 19119 7296
rect 19061 7287 19119 7293
rect 20180 7268 20208 7296
rect 24578 7284 24584 7296
rect 24636 7284 24642 7336
rect 24670 7284 24676 7336
rect 24728 7324 24734 7336
rect 24848 7327 24906 7333
rect 24848 7324 24860 7327
rect 24728 7296 24860 7324
rect 24728 7284 24734 7296
rect 24848 7293 24860 7296
rect 24894 7324 24906 7327
rect 25406 7324 25412 7336
rect 24894 7296 25412 7324
rect 24894 7293 24906 7296
rect 24848 7287 24906 7293
rect 25406 7284 25412 7296
rect 25464 7284 25470 7336
rect 29540 7327 29598 7333
rect 29540 7293 29552 7327
rect 29586 7324 29598 7327
rect 30098 7324 30104 7336
rect 29586 7296 30104 7324
rect 29586 7293 29598 7296
rect 29540 7287 29598 7293
rect 30098 7284 30104 7296
rect 30156 7284 30162 7336
rect 34882 7284 34888 7336
rect 34940 7324 34946 7336
rect 35253 7327 35311 7333
rect 35253 7324 35265 7327
rect 34940 7296 35265 7324
rect 34940 7284 34946 7296
rect 35253 7293 35265 7296
rect 35299 7324 35311 7327
rect 35342 7324 35348 7336
rect 35299 7296 35348 7324
rect 35299 7293 35311 7296
rect 35253 7287 35311 7293
rect 35342 7284 35348 7296
rect 35400 7284 35406 7336
rect 36630 7284 36636 7336
rect 36688 7324 36694 7336
rect 36817 7327 36875 7333
rect 36817 7324 36829 7327
rect 36688 7296 36829 7324
rect 36688 7284 36694 7296
rect 36817 7293 36829 7296
rect 36863 7293 36875 7327
rect 36817 7287 36875 7293
rect 11974 7216 11980 7268
rect 12032 7256 12038 7268
rect 12682 7259 12740 7265
rect 12682 7256 12694 7259
rect 12032 7228 12694 7256
rect 12032 7216 12038 7228
rect 12682 7225 12694 7228
rect 12728 7256 12740 7259
rect 12894 7256 12900 7268
rect 12728 7228 12900 7256
rect 12728 7225 12740 7228
rect 12682 7219 12740 7225
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 16666 7256 16672 7268
rect 16627 7228 16672 7256
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 18693 7259 18751 7265
rect 18693 7225 18705 7259
rect 18739 7256 18751 7259
rect 20162 7256 20168 7268
rect 18739 7228 19840 7256
rect 20123 7228 20168 7256
rect 18739 7225 18751 7228
rect 18693 7219 18751 7225
rect 13817 7191 13875 7197
rect 13817 7188 13829 7191
rect 11256 7160 13829 7188
rect 10468 7148 10474 7160
rect 13817 7157 13829 7160
rect 13863 7157 13875 7191
rect 13817 7151 13875 7157
rect 17310 7148 17316 7200
rect 17368 7188 17374 7200
rect 17589 7191 17647 7197
rect 17589 7188 17601 7191
rect 17368 7160 17601 7188
rect 17368 7148 17374 7160
rect 17589 7157 17601 7160
rect 17635 7188 17647 7191
rect 18230 7188 18236 7200
rect 17635 7160 18236 7188
rect 17635 7157 17647 7160
rect 17589 7151 17647 7157
rect 18230 7148 18236 7160
rect 18288 7148 18294 7200
rect 19812 7188 19840 7228
rect 20162 7216 20168 7228
rect 20220 7216 20226 7268
rect 21174 7216 21180 7268
rect 21232 7256 21238 7268
rect 21330 7259 21388 7265
rect 21330 7256 21342 7259
rect 21232 7228 21342 7256
rect 21232 7216 21238 7228
rect 21330 7225 21342 7228
rect 21376 7256 21388 7259
rect 22922 7256 22928 7268
rect 21376 7228 22928 7256
rect 21376 7225 21388 7228
rect 21330 7219 21388 7225
rect 22922 7216 22928 7228
rect 22980 7216 22986 7268
rect 24121 7259 24179 7265
rect 24121 7225 24133 7259
rect 24167 7256 24179 7259
rect 24688 7256 24716 7284
rect 24167 7228 24716 7256
rect 26605 7259 26663 7265
rect 24167 7225 24179 7228
rect 24121 7219 24179 7225
rect 26605 7225 26617 7259
rect 26651 7256 26663 7259
rect 27246 7256 27252 7268
rect 26651 7228 27252 7256
rect 26651 7225 26663 7228
rect 26605 7219 26663 7225
rect 27246 7216 27252 7228
rect 27304 7256 27310 7268
rect 27433 7259 27491 7265
rect 27433 7256 27445 7259
rect 27304 7228 27445 7256
rect 27304 7216 27310 7228
rect 27433 7225 27445 7228
rect 27479 7225 27491 7259
rect 27433 7219 27491 7225
rect 27709 7259 27767 7265
rect 27709 7225 27721 7259
rect 27755 7256 27767 7259
rect 27982 7256 27988 7268
rect 27755 7228 27988 7256
rect 27755 7225 27767 7228
rect 27709 7219 27767 7225
rect 27982 7216 27988 7228
rect 28040 7216 28046 7268
rect 31849 7259 31907 7265
rect 31849 7225 31861 7259
rect 31895 7256 31907 7259
rect 32554 7259 32612 7265
rect 32554 7256 32566 7259
rect 31895 7228 32566 7256
rect 31895 7225 31907 7228
rect 31849 7219 31907 7225
rect 32554 7225 32566 7228
rect 32600 7256 32612 7259
rect 33042 7256 33048 7268
rect 32600 7228 33048 7256
rect 32600 7225 32612 7228
rect 32554 7219 32612 7225
rect 33042 7216 33048 7228
rect 33100 7216 33106 7268
rect 35526 7256 35532 7268
rect 35487 7228 35532 7256
rect 35526 7216 35532 7228
rect 35584 7216 35590 7268
rect 36446 7216 36452 7268
rect 36504 7256 36510 7268
rect 36998 7256 37004 7268
rect 36504 7228 37004 7256
rect 36504 7216 36510 7228
rect 36998 7216 37004 7228
rect 37056 7216 37062 7268
rect 20073 7191 20131 7197
rect 20073 7188 20085 7191
rect 19812 7160 20085 7188
rect 20073 7157 20085 7160
rect 20119 7188 20131 7191
rect 20622 7188 20628 7200
rect 20119 7160 20628 7188
rect 20119 7157 20131 7160
rect 20073 7151 20131 7157
rect 20622 7148 20628 7160
rect 20680 7148 20686 7200
rect 22462 7188 22468 7200
rect 22423 7160 22468 7188
rect 22462 7148 22468 7160
rect 22520 7148 22526 7200
rect 23106 7188 23112 7200
rect 23019 7160 23112 7188
rect 23106 7148 23112 7160
rect 23164 7188 23170 7200
rect 24489 7191 24547 7197
rect 24489 7188 24501 7191
rect 23164 7160 24501 7188
rect 23164 7148 23170 7160
rect 24489 7157 24501 7160
rect 24535 7188 24547 7191
rect 24578 7188 24584 7200
rect 24535 7160 24584 7188
rect 24535 7157 24547 7160
rect 24489 7151 24547 7157
rect 24578 7148 24584 7160
rect 24636 7188 24642 7200
rect 24762 7188 24768 7200
rect 24636 7160 24768 7188
rect 24636 7148 24642 7160
rect 24762 7148 24768 7160
rect 24820 7148 24826 7200
rect 26878 7188 26884 7200
rect 26839 7160 26884 7188
rect 26878 7148 26884 7160
rect 26936 7188 26942 7200
rect 27617 7191 27675 7197
rect 27617 7188 27629 7191
rect 26936 7160 27629 7188
rect 26936 7148 26942 7160
rect 27617 7157 27629 7160
rect 27663 7157 27675 7191
rect 30650 7188 30656 7200
rect 30611 7160 30656 7188
rect 27617 7151 27675 7157
rect 30650 7148 30656 7160
rect 30708 7148 30714 7200
rect 33686 7148 33692 7200
rect 33744 7188 33750 7200
rect 33962 7188 33968 7200
rect 33744 7160 33968 7188
rect 33744 7148 33750 7160
rect 33962 7148 33968 7160
rect 34020 7148 34026 7200
rect 34330 7188 34336 7200
rect 34291 7160 34336 7188
rect 34330 7148 34336 7160
rect 34388 7148 34394 7200
rect 34698 7188 34704 7200
rect 34611 7160 34704 7188
rect 34698 7148 34704 7160
rect 34756 7188 34762 7200
rect 35437 7191 35495 7197
rect 35437 7188 35449 7191
rect 34756 7160 35449 7188
rect 34756 7148 34762 7160
rect 35437 7157 35449 7160
rect 35483 7157 35495 7191
rect 35437 7151 35495 7157
rect 35986 7148 35992 7200
rect 36044 7188 36050 7200
rect 36357 7191 36415 7197
rect 36357 7188 36369 7191
rect 36044 7160 36369 7188
rect 36044 7148 36050 7160
rect 36357 7157 36369 7160
rect 36403 7188 36415 7191
rect 36630 7188 36636 7200
rect 36403 7160 36636 7188
rect 36403 7157 36415 7160
rect 36357 7151 36415 7157
rect 36630 7148 36636 7160
rect 36688 7148 36694 7200
rect 1104 7098 38824 7120
rect 1104 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 27648 7098
rect 27700 7046 27712 7098
rect 27764 7046 27776 7098
rect 27828 7046 27840 7098
rect 27892 7046 38824 7098
rect 1104 7024 38824 7046
rect 2406 6944 2412 6996
rect 2464 6984 2470 6996
rect 2869 6987 2927 6993
rect 2869 6984 2881 6987
rect 2464 6956 2881 6984
rect 2464 6944 2470 6956
rect 2869 6953 2881 6956
rect 2915 6953 2927 6987
rect 2869 6947 2927 6953
rect 3050 6944 3056 6996
rect 3108 6984 3114 6996
rect 3789 6987 3847 6993
rect 3789 6984 3801 6987
rect 3108 6956 3801 6984
rect 3108 6944 3114 6956
rect 3789 6953 3801 6956
rect 3835 6953 3847 6987
rect 6730 6984 6736 6996
rect 6691 6956 6736 6984
rect 3789 6947 3847 6953
rect 6730 6944 6736 6956
rect 6788 6984 6794 6996
rect 7929 6987 7987 6993
rect 7929 6984 7941 6987
rect 6788 6956 7941 6984
rect 6788 6944 6794 6956
rect 7929 6953 7941 6956
rect 7975 6953 7987 6987
rect 7929 6947 7987 6953
rect 10134 6944 10140 6996
rect 10192 6984 10198 6996
rect 10229 6987 10287 6993
rect 10229 6984 10241 6987
rect 10192 6956 10241 6984
rect 10192 6944 10198 6956
rect 10229 6953 10241 6956
rect 10275 6984 10287 6987
rect 10686 6984 10692 6996
rect 10275 6956 10692 6984
rect 10275 6953 10287 6956
rect 10229 6947 10287 6953
rect 10686 6944 10692 6956
rect 10744 6944 10750 6996
rect 11790 6944 11796 6996
rect 11848 6984 11854 6996
rect 11885 6987 11943 6993
rect 11885 6984 11897 6987
rect 11848 6956 11897 6984
rect 11848 6944 11854 6956
rect 11885 6953 11897 6956
rect 11931 6953 11943 6987
rect 11885 6947 11943 6953
rect 16758 6944 16764 6996
rect 16816 6984 16822 6996
rect 17129 6987 17187 6993
rect 17129 6984 17141 6987
rect 16816 6956 17141 6984
rect 16816 6944 16822 6956
rect 17129 6953 17141 6956
rect 17175 6984 17187 6987
rect 17402 6984 17408 6996
rect 17175 6956 17408 6984
rect 17175 6953 17187 6956
rect 17129 6947 17187 6953
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 21174 6984 21180 6996
rect 21135 6956 21180 6984
rect 21174 6944 21180 6956
rect 21232 6944 21238 6996
rect 23661 6987 23719 6993
rect 23661 6953 23673 6987
rect 23707 6984 23719 6987
rect 23934 6984 23940 6996
rect 23707 6956 23940 6984
rect 23707 6953 23719 6956
rect 23661 6947 23719 6953
rect 23934 6944 23940 6956
rect 23992 6984 23998 6996
rect 24670 6984 24676 6996
rect 23992 6956 24676 6984
rect 23992 6944 23998 6956
rect 24670 6944 24676 6956
rect 24728 6944 24734 6996
rect 25958 6984 25964 6996
rect 25919 6956 25964 6984
rect 25958 6944 25964 6956
rect 26016 6944 26022 6996
rect 27065 6987 27123 6993
rect 27065 6953 27077 6987
rect 27111 6953 27123 6987
rect 27065 6947 27123 6953
rect 3326 6876 3332 6928
rect 3384 6916 3390 6928
rect 3970 6916 3976 6928
rect 3384 6888 3976 6916
rect 3384 6876 3390 6888
rect 3970 6876 3976 6888
rect 4028 6876 4034 6928
rect 5905 6919 5963 6925
rect 5905 6885 5917 6919
rect 5951 6916 5963 6919
rect 6270 6916 6276 6928
rect 5951 6888 6276 6916
rect 5951 6885 5963 6888
rect 5905 6879 5963 6885
rect 6270 6876 6276 6888
rect 6328 6876 6334 6928
rect 7006 6876 7012 6928
rect 7064 6916 7070 6928
rect 7285 6919 7343 6925
rect 7285 6916 7297 6919
rect 7064 6888 7297 6916
rect 7064 6876 7070 6888
rect 7285 6885 7297 6888
rect 7331 6885 7343 6919
rect 7285 6879 7343 6885
rect 7469 6919 7527 6925
rect 7469 6885 7481 6919
rect 7515 6916 7527 6919
rect 7558 6916 7564 6928
rect 7515 6888 7564 6916
rect 7515 6885 7527 6888
rect 7469 6879 7527 6885
rect 7558 6876 7564 6888
rect 7616 6876 7622 6928
rect 9766 6876 9772 6928
rect 9824 6916 9830 6928
rect 10045 6919 10103 6925
rect 10045 6916 10057 6919
rect 9824 6888 10057 6916
rect 9824 6876 9830 6888
rect 10045 6885 10057 6888
rect 10091 6885 10103 6919
rect 10045 6879 10103 6885
rect 13449 6919 13507 6925
rect 13449 6885 13461 6919
rect 13495 6885 13507 6919
rect 13449 6879 13507 6885
rect 1486 6848 1492 6860
rect 1447 6820 1492 6848
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 1762 6857 1768 6860
rect 1756 6848 1768 6857
rect 1723 6820 1768 6848
rect 1756 6811 1768 6820
rect 1762 6808 1768 6811
rect 1820 6808 1826 6860
rect 3786 6808 3792 6860
rect 3844 6848 3850 6860
rect 4065 6851 4123 6857
rect 4065 6848 4077 6851
rect 3844 6820 4077 6848
rect 3844 6808 3850 6820
rect 4065 6817 4077 6820
rect 4111 6817 4123 6851
rect 4065 6811 4123 6817
rect 5074 6808 5080 6860
rect 5132 6848 5138 6860
rect 5721 6851 5779 6857
rect 5721 6848 5733 6851
rect 5132 6820 5733 6848
rect 5132 6808 5138 6820
rect 5721 6817 5733 6820
rect 5767 6848 5779 6851
rect 8481 6851 8539 6857
rect 8481 6848 8493 6851
rect 5767 6820 8493 6848
rect 5767 6817 5779 6820
rect 5721 6811 5779 6817
rect 8481 6817 8493 6820
rect 8527 6817 8539 6851
rect 8938 6848 8944 6860
rect 8899 6820 8944 6848
rect 8481 6811 8539 6817
rect 8938 6808 8944 6820
rect 8996 6808 9002 6860
rect 10689 6851 10747 6857
rect 10689 6848 10701 6851
rect 9416 6820 10701 6848
rect 4706 6780 4712 6792
rect 4619 6752 4712 6780
rect 4706 6740 4712 6752
rect 4764 6780 4770 6792
rect 5261 6783 5319 6789
rect 5261 6780 5273 6783
rect 4764 6752 5273 6780
rect 4764 6740 4770 6752
rect 5261 6749 5273 6752
rect 5307 6780 5319 6783
rect 5810 6780 5816 6792
rect 5307 6752 5816 6780
rect 5307 6749 5319 6752
rect 5261 6743 5319 6749
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 5902 6740 5908 6792
rect 5960 6780 5966 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 5960 6752 6009 6780
rect 5960 6740 5966 6752
rect 5997 6749 6009 6752
rect 6043 6780 6055 6783
rect 6365 6783 6423 6789
rect 6365 6780 6377 6783
rect 6043 6752 6377 6780
rect 6043 6749 6055 6752
rect 5997 6743 6055 6749
rect 6365 6749 6377 6752
rect 6411 6780 6423 6783
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 6411 6752 7573 6780
rect 6411 6749 6423 6752
rect 6365 6743 6423 6749
rect 7561 6749 7573 6752
rect 7607 6780 7619 6783
rect 7742 6780 7748 6792
rect 7607 6752 7748 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 7742 6740 7748 6752
rect 7800 6780 7806 6792
rect 9416 6789 9444 6820
rect 10689 6817 10701 6820
rect 10735 6848 10747 6851
rect 10778 6848 10784 6860
rect 10735 6820 10784 6848
rect 10735 6817 10747 6820
rect 10689 6811 10747 6817
rect 10778 6808 10784 6820
rect 10836 6808 10842 6860
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 11701 6851 11759 6857
rect 11701 6848 11713 6851
rect 11112 6820 11713 6848
rect 11112 6808 11118 6820
rect 11701 6817 11713 6820
rect 11747 6848 11759 6851
rect 12158 6848 12164 6860
rect 11747 6820 12164 6848
rect 11747 6817 11759 6820
rect 11701 6811 11759 6817
rect 12158 6808 12164 6820
rect 12216 6808 12222 6860
rect 12986 6808 12992 6860
rect 13044 6848 13050 6860
rect 13464 6848 13492 6879
rect 21082 6876 21088 6928
rect 21140 6916 21146 6928
rect 22094 6916 22100 6928
rect 21140 6888 22100 6916
rect 21140 6876 21146 6888
rect 22094 6876 22100 6888
rect 22152 6916 22158 6928
rect 23106 6916 23112 6928
rect 22152 6888 23112 6916
rect 22152 6876 22158 6888
rect 13044 6820 13492 6848
rect 16016 6851 16074 6857
rect 13044 6808 13050 6820
rect 16016 6817 16028 6851
rect 16062 6848 16074 6851
rect 16482 6848 16488 6860
rect 16062 6820 16488 6848
rect 16062 6817 16074 6820
rect 16016 6811 16074 6817
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 17402 6808 17408 6860
rect 17460 6848 17466 6860
rect 22296 6857 22324 6888
rect 23106 6876 23112 6888
rect 23164 6876 23170 6928
rect 25409 6919 25467 6925
rect 25409 6885 25421 6919
rect 25455 6885 25467 6919
rect 25409 6879 25467 6885
rect 18489 6851 18547 6857
rect 18489 6848 18501 6851
rect 17460 6820 18501 6848
rect 17460 6808 17466 6820
rect 18489 6817 18501 6820
rect 18535 6817 18547 6851
rect 18489 6811 18547 6817
rect 22281 6851 22339 6857
rect 22281 6817 22293 6851
rect 22327 6817 22339 6851
rect 22281 6811 22339 6817
rect 22370 6808 22376 6860
rect 22428 6848 22434 6860
rect 22537 6851 22595 6857
rect 22537 6848 22549 6851
rect 22428 6820 22549 6848
rect 22428 6808 22434 6820
rect 22537 6817 22549 6820
rect 22583 6817 22595 6851
rect 24210 6848 24216 6860
rect 24171 6820 24216 6848
rect 22537 6811 22595 6817
rect 24210 6808 24216 6820
rect 24268 6808 24274 6860
rect 25222 6808 25228 6860
rect 25280 6848 25286 6860
rect 25424 6848 25452 6879
rect 27080 6860 27108 6947
rect 27246 6944 27252 6996
rect 27304 6984 27310 6996
rect 28077 6987 28135 6993
rect 28077 6984 28089 6987
rect 27304 6956 28089 6984
rect 27304 6944 27310 6956
rect 28077 6953 28089 6956
rect 28123 6953 28135 6987
rect 32306 6984 32312 6996
rect 32267 6956 32312 6984
rect 28077 6947 28135 6953
rect 32306 6944 32312 6956
rect 32364 6944 32370 6996
rect 33778 6984 33784 6996
rect 33739 6956 33784 6984
rect 33778 6944 33784 6956
rect 33836 6944 33842 6996
rect 29086 6916 29092 6928
rect 28920 6888 29092 6916
rect 25280 6820 25452 6848
rect 25280 6808 25286 6820
rect 26786 6808 26792 6860
rect 26844 6848 26850 6860
rect 26881 6851 26939 6857
rect 26881 6848 26893 6851
rect 26844 6820 26893 6848
rect 26844 6808 26850 6820
rect 26881 6817 26893 6820
rect 26927 6817 26939 6851
rect 26881 6811 26939 6817
rect 27062 6808 27068 6860
rect 27120 6808 27126 6860
rect 28813 6851 28871 6857
rect 28813 6817 28825 6851
rect 28859 6848 28871 6851
rect 28920 6848 28948 6888
rect 29086 6876 29092 6888
rect 29144 6876 29150 6928
rect 30650 6916 30656 6928
rect 30300 6888 30656 6916
rect 28859 6820 28948 6848
rect 28859 6817 28871 6820
rect 28813 6811 28871 6817
rect 29178 6808 29184 6860
rect 29236 6848 29242 6860
rect 29362 6857 29368 6860
rect 29345 6851 29368 6857
rect 29345 6848 29357 6851
rect 29236 6820 29357 6848
rect 29236 6808 29242 6820
rect 29345 6817 29357 6820
rect 29420 6848 29426 6860
rect 30300 6848 30328 6888
rect 30650 6876 30656 6888
rect 30708 6876 30714 6928
rect 33321 6919 33379 6925
rect 33321 6885 33333 6919
rect 33367 6885 33379 6919
rect 33321 6879 33379 6885
rect 33413 6919 33471 6925
rect 33413 6885 33425 6919
rect 33459 6916 33471 6919
rect 33594 6916 33600 6928
rect 33459 6888 33600 6916
rect 33459 6885 33471 6888
rect 33413 6879 33471 6885
rect 29420 6820 30328 6848
rect 29345 6811 29368 6817
rect 29362 6808 29368 6811
rect 29420 6808 29426 6820
rect 33134 6808 33140 6860
rect 33192 6848 33198 6860
rect 33336 6848 33364 6879
rect 33594 6876 33600 6888
rect 33652 6876 33658 6928
rect 34882 6916 34888 6928
rect 34843 6888 34888 6916
rect 34882 6876 34888 6888
rect 34940 6876 34946 6928
rect 36078 6876 36084 6928
rect 36136 6916 36142 6928
rect 36354 6916 36360 6928
rect 36136 6888 36360 6916
rect 36136 6876 36142 6888
rect 36354 6876 36360 6888
rect 36412 6916 36418 6928
rect 36449 6919 36507 6925
rect 36449 6916 36461 6919
rect 36412 6888 36461 6916
rect 36412 6876 36418 6888
rect 36449 6885 36461 6888
rect 36495 6885 36507 6919
rect 36449 6879 36507 6885
rect 33192 6820 33364 6848
rect 33192 6808 33198 6820
rect 34054 6808 34060 6860
rect 34112 6848 34118 6860
rect 34330 6848 34336 6860
rect 34112 6820 34336 6848
rect 34112 6808 34118 6820
rect 34330 6808 34336 6820
rect 34388 6848 34394 6860
rect 34977 6851 35035 6857
rect 34977 6848 34989 6851
rect 34388 6820 34989 6848
rect 34388 6808 34394 6820
rect 34977 6817 34989 6820
rect 35023 6848 35035 6851
rect 35526 6848 35532 6860
rect 35023 6820 35532 6848
rect 35023 6817 35035 6820
rect 34977 6811 35035 6817
rect 35526 6808 35532 6820
rect 35584 6848 35590 6860
rect 35713 6851 35771 6857
rect 35713 6848 35725 6851
rect 35584 6820 35725 6848
rect 35584 6808 35590 6820
rect 35713 6817 35725 6820
rect 35759 6848 35771 6851
rect 36541 6851 36599 6857
rect 36541 6848 36553 6851
rect 35759 6820 36553 6848
rect 35759 6817 35771 6820
rect 35713 6811 35771 6817
rect 36541 6817 36553 6820
rect 36587 6817 36599 6851
rect 36541 6811 36599 6817
rect 8297 6783 8355 6789
rect 8297 6780 8309 6783
rect 7800 6752 8309 6780
rect 7800 6740 7806 6752
rect 8297 6749 8309 6752
rect 8343 6780 8355 6783
rect 9401 6783 9459 6789
rect 9401 6780 9413 6783
rect 8343 6752 9413 6780
rect 8343 6749 8355 6752
rect 8297 6743 8355 6749
rect 9401 6749 9413 6752
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 9582 6740 9588 6792
rect 9640 6780 9646 6792
rect 9858 6780 9864 6792
rect 9640 6752 9864 6780
rect 9640 6740 9646 6752
rect 9858 6740 9864 6752
rect 9916 6780 9922 6792
rect 10321 6783 10379 6789
rect 10321 6780 10333 6783
rect 9916 6752 10333 6780
rect 9916 6740 9922 6752
rect 10321 6749 10333 6752
rect 10367 6749 10379 6783
rect 10321 6743 10379 6749
rect 11146 6740 11152 6792
rect 11204 6780 11210 6792
rect 11204 6752 11468 6780
rect 11204 6740 11210 6752
rect 4154 6672 4160 6724
rect 4212 6712 4218 6724
rect 4249 6715 4307 6721
rect 4249 6712 4261 6715
rect 4212 6684 4261 6712
rect 4212 6672 4218 6684
rect 4249 6681 4261 6684
rect 4295 6681 4307 6715
rect 4249 6675 4307 6681
rect 5718 6672 5724 6724
rect 5776 6712 5782 6724
rect 11440 6721 11468 6752
rect 11974 6740 11980 6792
rect 12032 6780 12038 6792
rect 13354 6780 13360 6792
rect 12032 6752 12077 6780
rect 13315 6752 13360 6780
rect 12032 6740 12038 6752
rect 13354 6740 13360 6752
rect 13412 6740 13418 6792
rect 13538 6780 13544 6792
rect 13499 6752 13544 6780
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 15102 6740 15108 6792
rect 15160 6780 15166 6792
rect 15654 6780 15660 6792
rect 15160 6752 15660 6780
rect 15160 6740 15166 6752
rect 15654 6740 15660 6752
rect 15712 6780 15718 6792
rect 15749 6783 15807 6789
rect 15749 6780 15761 6783
rect 15712 6752 15761 6780
rect 15712 6740 15718 6752
rect 15749 6749 15761 6752
rect 15795 6749 15807 6783
rect 18230 6780 18236 6792
rect 18191 6752 18236 6780
rect 15749 6743 15807 6749
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 25406 6780 25412 6792
rect 25367 6752 25412 6780
rect 25406 6740 25412 6752
rect 25464 6740 25470 6792
rect 25498 6740 25504 6792
rect 25556 6780 25562 6792
rect 27157 6783 27215 6789
rect 27157 6780 27169 6783
rect 25556 6752 27169 6780
rect 25556 6740 25562 6752
rect 27157 6749 27169 6752
rect 27203 6780 27215 6783
rect 27525 6783 27583 6789
rect 27525 6780 27537 6783
rect 27203 6752 27537 6780
rect 27203 6749 27215 6752
rect 27157 6743 27215 6749
rect 27525 6749 27537 6752
rect 27571 6780 27583 6783
rect 27798 6780 27804 6792
rect 27571 6752 27804 6780
rect 27571 6749 27583 6752
rect 27525 6743 27583 6749
rect 27798 6740 27804 6752
rect 27856 6740 27862 6792
rect 28994 6740 29000 6792
rect 29052 6780 29058 6792
rect 29089 6783 29147 6789
rect 29089 6780 29101 6783
rect 29052 6752 29101 6780
rect 29052 6740 29058 6752
rect 29089 6749 29101 6752
rect 29135 6749 29147 6783
rect 29089 6743 29147 6749
rect 33321 6783 33379 6789
rect 33321 6749 33333 6783
rect 33367 6780 33379 6783
rect 33686 6780 33692 6792
rect 33367 6752 33692 6780
rect 33367 6749 33379 6752
rect 33321 6743 33379 6749
rect 33686 6740 33692 6752
rect 33744 6780 33750 6792
rect 34146 6780 34152 6792
rect 33744 6752 34152 6780
rect 33744 6740 33750 6752
rect 34146 6740 34152 6752
rect 34204 6740 34210 6792
rect 34885 6783 34943 6789
rect 34885 6749 34897 6783
rect 34931 6780 34943 6783
rect 35066 6780 35072 6792
rect 34931 6752 35072 6780
rect 34931 6749 34943 6752
rect 34885 6743 34943 6749
rect 35066 6740 35072 6752
rect 35124 6740 35130 6792
rect 36354 6780 36360 6792
rect 36315 6752 36360 6780
rect 36354 6740 36360 6752
rect 36412 6740 36418 6792
rect 7009 6715 7067 6721
rect 7009 6712 7021 6715
rect 5776 6684 7021 6712
rect 5776 6672 5782 6684
rect 7009 6681 7021 6684
rect 7055 6681 7067 6715
rect 7009 6675 7067 6681
rect 11425 6715 11483 6721
rect 11425 6681 11437 6715
rect 11471 6681 11483 6715
rect 11425 6675 11483 6681
rect 11514 6672 11520 6724
rect 11572 6712 11578 6724
rect 12989 6715 13047 6721
rect 12989 6712 13001 6715
rect 11572 6684 13001 6712
rect 11572 6672 11578 6684
rect 12989 6681 13001 6684
rect 13035 6681 13047 6715
rect 24946 6712 24952 6724
rect 24907 6684 24952 6712
rect 12989 6675 13047 6681
rect 24946 6672 24952 6684
rect 25004 6712 25010 6724
rect 26237 6715 26295 6721
rect 26237 6712 26249 6715
rect 25004 6684 26249 6712
rect 25004 6672 25010 6684
rect 26237 6681 26249 6684
rect 26283 6681 26295 6715
rect 26237 6675 26295 6681
rect 30926 6672 30932 6724
rect 30984 6712 30990 6724
rect 32861 6715 32919 6721
rect 32861 6712 32873 6715
rect 30984 6684 32873 6712
rect 30984 6672 30990 6684
rect 32861 6681 32873 6684
rect 32907 6681 32919 6715
rect 32861 6675 32919 6681
rect 3513 6647 3571 6653
rect 3513 6613 3525 6647
rect 3559 6644 3571 6647
rect 3878 6644 3884 6656
rect 3559 6616 3884 6644
rect 3559 6613 3571 6616
rect 3513 6607 3571 6613
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 5442 6644 5448 6656
rect 5403 6616 5448 6644
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 9769 6647 9827 6653
rect 9769 6644 9781 6647
rect 9732 6616 9781 6644
rect 9732 6604 9738 6616
rect 9769 6613 9781 6616
rect 9815 6613 9827 6647
rect 9769 6607 9827 6613
rect 11149 6647 11207 6653
rect 11149 6613 11161 6647
rect 11195 6644 11207 6647
rect 11330 6644 11336 6656
rect 11195 6616 11336 6644
rect 11195 6613 11207 6616
rect 11149 6607 11207 6613
rect 11330 6604 11336 6616
rect 11388 6604 11394 6656
rect 12618 6644 12624 6656
rect 12579 6616 12624 6644
rect 12618 6604 12624 6616
rect 12676 6604 12682 6656
rect 15378 6604 15384 6656
rect 15436 6644 15442 6656
rect 15473 6647 15531 6653
rect 15473 6644 15485 6647
rect 15436 6616 15485 6644
rect 15436 6604 15442 6616
rect 15473 6613 15485 6616
rect 15519 6613 15531 6647
rect 15473 6607 15531 6613
rect 17586 6604 17592 6656
rect 17644 6644 17650 6656
rect 17773 6647 17831 6653
rect 17773 6644 17785 6647
rect 17644 6616 17785 6644
rect 17644 6604 17650 6616
rect 17773 6613 17785 6616
rect 17819 6644 17831 6647
rect 18049 6647 18107 6653
rect 18049 6644 18061 6647
rect 17819 6616 18061 6644
rect 17819 6613 17831 6616
rect 17773 6607 17831 6613
rect 18049 6613 18061 6616
rect 18095 6644 18107 6647
rect 18506 6644 18512 6656
rect 18095 6616 18512 6644
rect 18095 6613 18107 6616
rect 18049 6607 18107 6613
rect 18506 6604 18512 6616
rect 18564 6644 18570 6656
rect 19613 6647 19671 6653
rect 19613 6644 19625 6647
rect 18564 6616 19625 6644
rect 18564 6604 18570 6616
rect 19613 6613 19625 6616
rect 19659 6613 19671 6647
rect 26602 6644 26608 6656
rect 26563 6616 26608 6644
rect 19613 6607 19671 6613
rect 26602 6604 26608 6616
rect 26660 6604 26666 6656
rect 27890 6644 27896 6656
rect 27851 6616 27896 6644
rect 27890 6604 27896 6616
rect 27948 6604 27954 6656
rect 30466 6644 30472 6656
rect 30427 6616 30472 6644
rect 30466 6604 30472 6616
rect 30524 6604 30530 6656
rect 33870 6604 33876 6656
rect 33928 6644 33934 6656
rect 34425 6647 34483 6653
rect 34425 6644 34437 6647
rect 33928 6616 34437 6644
rect 33928 6604 33934 6616
rect 34425 6613 34437 6616
rect 34471 6613 34483 6647
rect 34425 6607 34483 6613
rect 35250 6604 35256 6656
rect 35308 6644 35314 6656
rect 35345 6647 35403 6653
rect 35345 6644 35357 6647
rect 35308 6616 35357 6644
rect 35308 6604 35314 6616
rect 35345 6613 35357 6616
rect 35391 6613 35403 6647
rect 35986 6644 35992 6656
rect 35947 6616 35992 6644
rect 35345 6607 35403 6613
rect 35986 6604 35992 6616
rect 36044 6604 36050 6656
rect 36538 6604 36544 6656
rect 36596 6644 36602 6656
rect 36909 6647 36967 6653
rect 36909 6644 36921 6647
rect 36596 6616 36921 6644
rect 36596 6604 36602 6616
rect 36909 6613 36921 6616
rect 36955 6613 36967 6647
rect 36909 6607 36967 6613
rect 1104 6554 38824 6576
rect 1104 6502 7648 6554
rect 7700 6502 7712 6554
rect 7764 6502 7776 6554
rect 7828 6502 7840 6554
rect 7892 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 34315 6554
rect 34367 6502 34379 6554
rect 34431 6502 34443 6554
rect 34495 6502 34507 6554
rect 34559 6502 38824 6554
rect 1104 6480 38824 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 1452 6412 1593 6440
rect 1452 6400 1458 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 1581 6403 1639 6409
rect 2041 6443 2099 6449
rect 2041 6409 2053 6443
rect 2087 6440 2099 6443
rect 2590 6440 2596 6452
rect 2087 6412 2596 6440
rect 2087 6409 2099 6412
rect 2041 6403 2099 6409
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2056 6236 2084 6403
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 3786 6400 3792 6452
rect 3844 6440 3850 6452
rect 4525 6443 4583 6449
rect 4525 6440 4537 6443
rect 3844 6412 4537 6440
rect 3844 6400 3850 6412
rect 4525 6409 4537 6412
rect 4571 6409 4583 6443
rect 5074 6440 5080 6452
rect 5035 6412 5080 6440
rect 4525 6403 4583 6409
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 6270 6440 6276 6452
rect 6231 6412 6276 6440
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 6638 6440 6644 6452
rect 6551 6412 6644 6440
rect 6638 6400 6644 6412
rect 6696 6440 6702 6452
rect 7006 6440 7012 6452
rect 6696 6412 7012 6440
rect 6696 6400 6702 6412
rect 7006 6400 7012 6412
rect 7064 6440 7070 6452
rect 8110 6440 8116 6452
rect 7064 6412 8116 6440
rect 7064 6400 7070 6412
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 9401 6443 9459 6449
rect 9401 6409 9413 6443
rect 9447 6440 9459 6443
rect 9766 6440 9772 6452
rect 9447 6412 9772 6440
rect 9447 6409 9459 6412
rect 9401 6403 9459 6409
rect 9766 6400 9772 6412
rect 9824 6400 9830 6452
rect 10134 6440 10140 6452
rect 10095 6412 10140 6440
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 11790 6440 11796 6452
rect 11751 6412 11796 6440
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 12158 6440 12164 6452
rect 12119 6412 12164 6440
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 13538 6400 13544 6452
rect 13596 6440 13602 6452
rect 14553 6443 14611 6449
rect 14553 6440 14565 6443
rect 13596 6412 14565 6440
rect 13596 6400 13602 6412
rect 14553 6409 14565 6412
rect 14599 6409 14611 6443
rect 17402 6440 17408 6452
rect 17363 6412 17408 6440
rect 14553 6403 14611 6409
rect 17402 6400 17408 6412
rect 17460 6400 17466 6452
rect 18230 6400 18236 6452
rect 18288 6440 18294 6452
rect 19061 6443 19119 6449
rect 19061 6440 19073 6443
rect 18288 6412 19073 6440
rect 18288 6400 18294 6412
rect 19061 6409 19073 6412
rect 19107 6409 19119 6443
rect 19061 6403 19119 6409
rect 20993 6443 21051 6449
rect 20993 6409 21005 6443
rect 21039 6440 21051 6443
rect 22094 6440 22100 6452
rect 21039 6412 22100 6440
rect 21039 6409 21051 6412
rect 20993 6403 21051 6409
rect 5261 6375 5319 6381
rect 5261 6341 5273 6375
rect 5307 6372 5319 6375
rect 5994 6372 6000 6384
rect 5307 6344 6000 6372
rect 5307 6341 5319 6344
rect 5261 6335 5319 6341
rect 5994 6332 6000 6344
rect 6052 6332 6058 6384
rect 10873 6375 10931 6381
rect 10873 6341 10885 6375
rect 10919 6372 10931 6375
rect 11054 6372 11060 6384
rect 10919 6344 11060 6372
rect 10919 6341 10931 6344
rect 10873 6335 10931 6341
rect 11054 6332 11060 6344
rect 11112 6332 11118 6384
rect 13998 6372 14004 6384
rect 13959 6344 14004 6372
rect 13998 6332 14004 6344
rect 14056 6332 14062 6384
rect 18138 6372 18144 6384
rect 18099 6344 18144 6372
rect 18138 6332 18144 6344
rect 18196 6332 18202 6384
rect 5442 6264 5448 6316
rect 5500 6304 5506 6316
rect 5721 6307 5779 6313
rect 5721 6304 5733 6307
rect 5500 6276 5733 6304
rect 5500 6264 5506 6276
rect 5721 6273 5733 6276
rect 5767 6304 5779 6307
rect 9769 6307 9827 6313
rect 5767 6276 6960 6304
rect 5767 6273 5779 6276
rect 5721 6267 5779 6273
rect 1443 6208 2084 6236
rect 2409 6239 2467 6245
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2409 6205 2421 6239
rect 2455 6236 2467 6239
rect 2593 6239 2651 6245
rect 2593 6236 2605 6239
rect 2455 6208 2605 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 2593 6205 2605 6208
rect 2639 6236 2651 6239
rect 3786 6236 3792 6248
rect 2639 6208 3792 6236
rect 2639 6205 2651 6208
rect 2593 6199 2651 6205
rect 3786 6196 3792 6208
rect 3844 6196 3850 6248
rect 5810 6236 5816 6248
rect 5771 6208 5816 6236
rect 5810 6196 5816 6208
rect 5868 6196 5874 6248
rect 6730 6196 6736 6248
rect 6788 6236 6794 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6788 6208 6837 6236
rect 6788 6196 6794 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 6932 6236 6960 6276
rect 9769 6273 9781 6307
rect 9815 6304 9827 6307
rect 9858 6304 9864 6316
rect 9815 6276 9864 6304
rect 9815 6273 9827 6276
rect 9769 6267 9827 6273
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 11333 6307 11391 6313
rect 11333 6304 11345 6307
rect 10100 6276 11345 6304
rect 10100 6264 10106 6276
rect 11333 6273 11345 6276
rect 11379 6304 11391 6307
rect 11514 6304 11520 6316
rect 11379 6276 11520 6304
rect 11379 6273 11391 6276
rect 11333 6267 11391 6273
rect 11514 6264 11520 6276
rect 11572 6264 11578 6316
rect 12618 6304 12624 6316
rect 12579 6276 12624 6304
rect 12618 6264 12624 6276
rect 12676 6264 12682 6316
rect 14016 6304 14044 6332
rect 21100 6313 21128 6412
rect 22094 6400 22100 6412
rect 22152 6400 22158 6452
rect 22370 6400 22376 6452
rect 22428 6440 22434 6452
rect 22465 6443 22523 6449
rect 22465 6440 22477 6443
rect 22428 6412 22477 6440
rect 22428 6400 22434 6412
rect 22465 6409 22477 6412
rect 22511 6409 22523 6443
rect 23106 6440 23112 6452
rect 23067 6412 23112 6440
rect 22465 6403 22523 6409
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 23934 6440 23940 6452
rect 23895 6412 23940 6440
rect 23934 6400 23940 6412
rect 23992 6400 23998 6452
rect 24118 6440 24124 6452
rect 24079 6412 24124 6440
rect 24118 6400 24124 6412
rect 24176 6400 24182 6452
rect 25133 6443 25191 6449
rect 25133 6409 25145 6443
rect 25179 6440 25191 6443
rect 25406 6440 25412 6452
rect 25179 6412 25412 6440
rect 25179 6409 25191 6412
rect 25133 6403 25191 6409
rect 25406 6400 25412 6412
rect 25464 6400 25470 6452
rect 27062 6400 27068 6452
rect 27120 6440 27126 6452
rect 27525 6443 27583 6449
rect 27525 6440 27537 6443
rect 27120 6412 27537 6440
rect 27120 6400 27126 6412
rect 27525 6409 27537 6412
rect 27571 6440 27583 6443
rect 28626 6440 28632 6452
rect 27571 6412 28632 6440
rect 27571 6409 27583 6412
rect 27525 6403 27583 6409
rect 28626 6400 28632 6412
rect 28684 6400 28690 6452
rect 28994 6440 29000 6452
rect 28955 6412 29000 6440
rect 28994 6400 29000 6412
rect 29052 6400 29058 6452
rect 33134 6400 33140 6452
rect 33192 6440 33198 6452
rect 33321 6443 33379 6449
rect 33321 6440 33333 6443
rect 33192 6412 33333 6440
rect 33192 6400 33198 6412
rect 33321 6409 33333 6412
rect 33367 6409 33379 6443
rect 34054 6440 34060 6452
rect 34015 6412 34060 6440
rect 33321 6403 33379 6409
rect 34054 6400 34060 6412
rect 34112 6400 34118 6452
rect 36538 6400 36544 6452
rect 36596 6440 36602 6452
rect 36633 6443 36691 6449
rect 36633 6440 36645 6443
rect 36596 6412 36645 6440
rect 36596 6400 36602 6412
rect 36633 6409 36645 6412
rect 36679 6409 36691 6443
rect 36633 6403 36691 6409
rect 27798 6332 27804 6384
rect 27856 6372 27862 6384
rect 27893 6375 27951 6381
rect 27893 6372 27905 6375
rect 27856 6344 27905 6372
rect 27856 6332 27862 6344
rect 27893 6341 27905 6344
rect 27939 6341 27951 6375
rect 27893 6335 27951 6341
rect 29365 6375 29423 6381
rect 29365 6341 29377 6375
rect 29411 6372 29423 6375
rect 30190 6372 30196 6384
rect 29411 6344 30196 6372
rect 29411 6341 29423 6344
rect 29365 6335 29423 6341
rect 30190 6332 30196 6344
rect 30248 6332 30254 6384
rect 33045 6375 33103 6381
rect 33045 6341 33057 6375
rect 33091 6372 33103 6375
rect 33594 6372 33600 6384
rect 33091 6344 33600 6372
rect 33091 6341 33103 6344
rect 33045 6335 33103 6341
rect 33594 6332 33600 6344
rect 33652 6332 33658 6384
rect 21085 6307 21143 6313
rect 14016 6276 15240 6304
rect 8757 6239 8815 6245
rect 8757 6236 8769 6239
rect 6932 6208 8769 6236
rect 6825 6199 6883 6205
rect 8757 6205 8769 6208
rect 8803 6205 8815 6239
rect 8757 6199 8815 6205
rect 10689 6239 10747 6245
rect 10689 6205 10701 6239
rect 10735 6236 10747 6239
rect 10778 6236 10784 6248
rect 10735 6208 10784 6236
rect 10735 6205 10747 6208
rect 10689 6199 10747 6205
rect 10778 6196 10784 6208
rect 10836 6236 10842 6248
rect 11422 6236 11428 6248
rect 10836 6208 11428 6236
rect 10836 6196 10842 6208
rect 11422 6196 11428 6208
rect 11480 6196 11486 6248
rect 12636 6236 12664 6264
rect 14921 6239 14979 6245
rect 14921 6236 14933 6239
rect 12636 6208 14933 6236
rect 14921 6205 14933 6208
rect 14967 6236 14979 6239
rect 15102 6236 15108 6248
rect 14967 6208 15108 6236
rect 14967 6205 14979 6208
rect 14921 6199 14979 6205
rect 15102 6196 15108 6208
rect 15160 6196 15166 6248
rect 15212 6236 15240 6276
rect 21085 6273 21097 6307
rect 21131 6273 21143 6307
rect 24486 6304 24492 6316
rect 24447 6276 24492 6304
rect 21085 6267 21143 6273
rect 24486 6264 24492 6276
rect 24544 6264 24550 6316
rect 24670 6304 24676 6316
rect 24631 6276 24676 6304
rect 24670 6264 24676 6276
rect 24728 6264 24734 6316
rect 25222 6264 25228 6316
rect 25280 6304 25286 6316
rect 25409 6307 25467 6313
rect 25409 6304 25421 6307
rect 25280 6276 25421 6304
rect 25280 6264 25286 6276
rect 25409 6273 25421 6276
rect 25455 6273 25467 6307
rect 29822 6304 29828 6316
rect 29783 6276 29828 6304
rect 25409 6267 25467 6273
rect 29822 6264 29828 6276
rect 29880 6264 29886 6316
rect 33226 6264 33232 6316
rect 33284 6304 33290 6316
rect 34333 6307 34391 6313
rect 34333 6304 34345 6307
rect 33284 6276 34345 6304
rect 33284 6264 33290 6276
rect 34333 6273 34345 6276
rect 34379 6304 34391 6307
rect 34882 6304 34888 6316
rect 34379 6276 34888 6304
rect 34379 6273 34391 6276
rect 34333 6267 34391 6273
rect 34882 6264 34888 6276
rect 34940 6264 34946 6316
rect 35066 6304 35072 6316
rect 35027 6276 35072 6304
rect 35066 6264 35072 6276
rect 35124 6264 35130 6316
rect 15378 6245 15384 6248
rect 15361 6239 15384 6245
rect 15361 6236 15373 6239
rect 15212 6208 15373 6236
rect 15361 6205 15373 6208
rect 15436 6236 15442 6248
rect 19429 6239 19487 6245
rect 19429 6236 19441 6239
rect 15436 6208 15509 6236
rect 18616 6208 19441 6236
rect 15361 6199 15384 6205
rect 15378 6196 15384 6199
rect 15436 6196 15442 6208
rect 18616 6180 18644 6208
rect 19429 6205 19441 6208
rect 19475 6205 19487 6239
rect 19429 6199 19487 6205
rect 23477 6239 23535 6245
rect 23477 6205 23489 6239
rect 23523 6236 23535 6239
rect 23523 6208 24624 6236
rect 23523 6205 23535 6208
rect 23477 6199 23535 6205
rect 24596 6180 24624 6208
rect 24854 6196 24860 6248
rect 24912 6236 24918 6248
rect 25593 6239 25651 6245
rect 25593 6236 25605 6239
rect 24912 6208 25605 6236
rect 24912 6196 24918 6208
rect 25593 6205 25605 6208
rect 25639 6236 25651 6239
rect 25682 6236 25688 6248
rect 25639 6208 25688 6236
rect 25639 6205 25651 6208
rect 25593 6199 25651 6205
rect 25682 6196 25688 6208
rect 25740 6196 25746 6248
rect 28721 6239 28779 6245
rect 28721 6205 28733 6239
rect 28767 6236 28779 6239
rect 29914 6236 29920 6248
rect 28767 6208 29920 6236
rect 28767 6205 28779 6208
rect 28721 6199 28779 6205
rect 29914 6196 29920 6208
rect 29972 6196 29978 6248
rect 30929 6239 30987 6245
rect 30929 6205 30941 6239
rect 30975 6236 30987 6239
rect 31021 6239 31079 6245
rect 31021 6236 31033 6239
rect 30975 6208 31033 6236
rect 30975 6205 30987 6208
rect 30929 6199 30987 6205
rect 31021 6205 31033 6208
rect 31067 6236 31079 6239
rect 32306 6236 32312 6248
rect 31067 6208 32312 6236
rect 31067 6205 31079 6208
rect 31021 6199 31079 6205
rect 32306 6196 32312 6208
rect 32364 6196 32370 6248
rect 34054 6196 34060 6248
rect 34112 6236 34118 6248
rect 34606 6236 34612 6248
rect 34112 6208 34612 6236
rect 34112 6196 34118 6208
rect 34606 6196 34612 6208
rect 34664 6236 34670 6248
rect 35250 6236 35256 6248
rect 34664 6208 35256 6236
rect 34664 6196 34670 6208
rect 35250 6196 35256 6208
rect 35308 6196 35314 6248
rect 35526 6245 35532 6248
rect 35520 6236 35532 6245
rect 35487 6208 35532 6236
rect 35520 6199 35532 6208
rect 35584 6236 35590 6248
rect 37185 6239 37243 6245
rect 37185 6236 37197 6239
rect 35584 6208 37197 6236
rect 35526 6196 35532 6199
rect 35584 6196 35590 6208
rect 37185 6205 37197 6208
rect 37231 6205 37243 6239
rect 37185 6199 37243 6205
rect 1762 6128 1768 6180
rect 1820 6168 1826 6180
rect 2860 6171 2918 6177
rect 1820 6140 2084 6168
rect 1820 6128 1826 6140
rect 2056 6100 2084 6140
rect 2860 6137 2872 6171
rect 2906 6168 2918 6171
rect 3050 6168 3056 6180
rect 2906 6140 3056 6168
rect 2906 6137 2918 6140
rect 2860 6131 2918 6137
rect 3050 6128 3056 6140
rect 3108 6128 3114 6180
rect 5718 6168 5724 6180
rect 5679 6140 5724 6168
rect 5718 6128 5724 6140
rect 5776 6128 5782 6180
rect 7006 6128 7012 6180
rect 7064 6177 7070 6180
rect 7064 6171 7128 6177
rect 7064 6137 7082 6171
rect 7116 6137 7128 6171
rect 11330 6168 11336 6180
rect 11291 6140 11336 6168
rect 7064 6131 7128 6137
rect 7064 6128 7070 6131
rect 11330 6128 11336 6140
rect 11388 6128 11394 6180
rect 12526 6128 12532 6180
rect 12584 6168 12590 6180
rect 12888 6171 12946 6177
rect 12888 6168 12900 6171
rect 12584 6140 12900 6168
rect 12584 6128 12590 6140
rect 12888 6137 12900 6140
rect 12934 6168 12946 6171
rect 13538 6168 13544 6180
rect 12934 6140 13544 6168
rect 12934 6137 12946 6140
rect 12888 6131 12946 6137
rect 13538 6128 13544 6140
rect 13596 6128 13602 6180
rect 18414 6168 18420 6180
rect 18327 6140 18420 6168
rect 18414 6128 18420 6140
rect 18472 6128 18478 6180
rect 18598 6168 18604 6180
rect 18559 6140 18604 6168
rect 18598 6128 18604 6140
rect 18656 6128 18662 6180
rect 18690 6128 18696 6180
rect 18748 6168 18754 6180
rect 20625 6171 20683 6177
rect 18748 6140 18793 6168
rect 18748 6128 18754 6140
rect 20625 6137 20637 6171
rect 20671 6168 20683 6171
rect 21330 6171 21388 6177
rect 21330 6168 21342 6171
rect 20671 6140 21342 6168
rect 20671 6137 20683 6140
rect 20625 6131 20683 6137
rect 21330 6137 21342 6140
rect 21376 6168 21388 6171
rect 21726 6168 21732 6180
rect 21376 6140 21732 6168
rect 21376 6137 21388 6140
rect 21330 6131 21388 6137
rect 21726 6128 21732 6140
rect 21784 6128 21790 6180
rect 24578 6168 24584 6180
rect 24539 6140 24584 6168
rect 24578 6128 24584 6140
rect 24636 6128 24642 6180
rect 25860 6171 25918 6177
rect 25860 6137 25872 6171
rect 25906 6168 25918 6171
rect 25958 6168 25964 6180
rect 25906 6140 25964 6168
rect 25906 6137 25918 6140
rect 25860 6131 25918 6137
rect 25958 6128 25964 6140
rect 26016 6128 26022 6180
rect 28169 6171 28227 6177
rect 28169 6137 28181 6171
rect 28215 6168 28227 6171
rect 28902 6168 28908 6180
rect 28215 6140 28908 6168
rect 28215 6137 28227 6140
rect 28169 6131 28227 6137
rect 28902 6128 28908 6140
rect 28960 6128 28966 6180
rect 30742 6128 30748 6180
rect 30800 6168 30806 6180
rect 31266 6171 31324 6177
rect 31266 6168 31278 6171
rect 30800 6140 31278 6168
rect 30800 6128 30806 6140
rect 31266 6137 31278 6140
rect 31312 6137 31324 6171
rect 31266 6131 31324 6137
rect 3970 6100 3976 6112
rect 2056 6072 3976 6100
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 8018 6060 8024 6112
rect 8076 6100 8082 6112
rect 8205 6103 8263 6109
rect 8205 6100 8217 6103
rect 8076 6072 8217 6100
rect 8076 6060 8082 6072
rect 8205 6069 8217 6072
rect 8251 6069 8263 6103
rect 16482 6100 16488 6112
rect 16443 6072 16488 6100
rect 8205 6063 8263 6069
rect 16482 6060 16488 6072
rect 16540 6100 16546 6112
rect 17037 6103 17095 6109
rect 17037 6100 17049 6103
rect 16540 6072 17049 6100
rect 16540 6060 16546 6072
rect 17037 6069 17049 6072
rect 17083 6069 17095 6103
rect 17037 6063 17095 6069
rect 17678 6060 17684 6112
rect 17736 6100 17742 6112
rect 17773 6103 17831 6109
rect 17773 6100 17785 6103
rect 17736 6072 17785 6100
rect 17736 6060 17742 6072
rect 17773 6069 17785 6072
rect 17819 6100 17831 6103
rect 18432 6100 18460 6128
rect 26970 6100 26976 6112
rect 17819 6072 18460 6100
rect 26931 6072 26976 6100
rect 17819 6069 17831 6072
rect 17773 6063 17831 6069
rect 26970 6060 26976 6072
rect 27028 6060 27034 6112
rect 29730 6060 29736 6112
rect 29788 6100 29794 6112
rect 29825 6103 29883 6109
rect 29825 6100 29837 6103
rect 29788 6072 29837 6100
rect 29788 6060 29794 6072
rect 29825 6069 29837 6072
rect 29871 6100 29883 6103
rect 30285 6103 30343 6109
rect 30285 6100 30297 6103
rect 29871 6072 30297 6100
rect 29871 6069 29883 6072
rect 29825 6063 29883 6069
rect 30285 6069 30297 6072
rect 30331 6069 30343 6103
rect 30285 6063 30343 6069
rect 32122 6060 32128 6112
rect 32180 6100 32186 6112
rect 32401 6103 32459 6109
rect 32401 6100 32413 6103
rect 32180 6072 32413 6100
rect 32180 6060 32186 6072
rect 32401 6069 32413 6072
rect 32447 6069 32459 6103
rect 32401 6063 32459 6069
rect 1104 6010 38824 6032
rect 1104 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 27648 6010
rect 27700 5958 27712 6010
rect 27764 5958 27776 6010
rect 27828 5958 27840 6010
rect 27892 5958 38824 6010
rect 1104 5936 38824 5958
rect 4249 5899 4307 5905
rect 4249 5865 4261 5899
rect 4295 5896 4307 5899
rect 4430 5896 4436 5908
rect 4295 5868 4436 5896
rect 4295 5865 4307 5868
rect 4249 5859 4307 5865
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 5445 5899 5503 5905
rect 5445 5865 5457 5899
rect 5491 5896 5503 5899
rect 5902 5896 5908 5908
rect 5491 5868 5908 5896
rect 5491 5865 5503 5868
rect 5445 5859 5503 5865
rect 5902 5856 5908 5868
rect 5960 5856 5966 5908
rect 6086 5896 6092 5908
rect 6047 5868 6092 5896
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 7009 5899 7067 5905
rect 7009 5865 7021 5899
rect 7055 5896 7067 5899
rect 7098 5896 7104 5908
rect 7055 5868 7104 5896
rect 7055 5865 7067 5868
rect 7009 5859 7067 5865
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 10042 5896 10048 5908
rect 10003 5868 10048 5896
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 11330 5856 11336 5908
rect 11388 5896 11394 5908
rect 11959 5899 12017 5905
rect 11959 5896 11971 5899
rect 11388 5868 11971 5896
rect 11388 5856 11394 5868
rect 11959 5865 11971 5868
rect 12005 5865 12017 5899
rect 11959 5859 12017 5865
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 12986 5896 12992 5908
rect 12492 5868 12537 5896
rect 12947 5868 12992 5896
rect 12492 5856 12498 5868
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 13354 5896 13360 5908
rect 13315 5868 13360 5896
rect 13354 5856 13360 5868
rect 13412 5856 13418 5908
rect 15654 5856 15660 5908
rect 15712 5896 15718 5908
rect 15749 5899 15807 5905
rect 15749 5896 15761 5899
rect 15712 5868 15761 5896
rect 15712 5856 15718 5868
rect 15749 5865 15761 5868
rect 15795 5865 15807 5899
rect 16666 5896 16672 5908
rect 16579 5868 16672 5896
rect 15749 5859 15807 5865
rect 16666 5856 16672 5868
rect 16724 5896 16730 5908
rect 17310 5896 17316 5908
rect 16724 5868 17316 5896
rect 16724 5856 16730 5868
rect 17310 5856 17316 5868
rect 17368 5856 17374 5908
rect 21634 5896 21640 5908
rect 21595 5868 21640 5896
rect 21634 5856 21640 5868
rect 21692 5856 21698 5908
rect 22370 5896 22376 5908
rect 22331 5868 22376 5896
rect 22370 5856 22376 5868
rect 22428 5896 22434 5908
rect 24857 5899 24915 5905
rect 24857 5896 24869 5899
rect 22428 5868 24869 5896
rect 22428 5856 22434 5868
rect 24857 5865 24869 5868
rect 24903 5896 24915 5899
rect 25498 5896 25504 5908
rect 24903 5868 25504 5896
rect 24903 5865 24915 5868
rect 24857 5859 24915 5865
rect 25498 5856 25504 5868
rect 25556 5856 25562 5908
rect 26786 5896 26792 5908
rect 26747 5868 26792 5896
rect 26786 5856 26792 5868
rect 26844 5856 26850 5908
rect 27430 5896 27436 5908
rect 27391 5868 27436 5896
rect 27430 5856 27436 5868
rect 27488 5856 27494 5908
rect 28527 5899 28585 5905
rect 28527 5865 28539 5899
rect 28573 5896 28585 5899
rect 29822 5896 29828 5908
rect 28573 5868 29828 5896
rect 28573 5865 28585 5868
rect 28527 5859 28585 5865
rect 29822 5856 29828 5868
rect 29880 5856 29886 5908
rect 30374 5856 30380 5908
rect 30432 5896 30438 5908
rect 30561 5899 30619 5905
rect 30561 5896 30573 5899
rect 30432 5868 30573 5896
rect 30432 5856 30438 5868
rect 30561 5865 30573 5868
rect 30607 5865 30619 5899
rect 33134 5896 33140 5908
rect 33047 5868 33140 5896
rect 30561 5859 30619 5865
rect 33134 5856 33140 5868
rect 33192 5896 33198 5908
rect 33870 5896 33876 5908
rect 33192 5868 33876 5896
rect 33192 5856 33198 5868
rect 33870 5856 33876 5868
rect 33928 5856 33934 5908
rect 35526 5896 35532 5908
rect 35487 5868 35532 5896
rect 35526 5856 35532 5868
rect 35584 5856 35590 5908
rect 36078 5896 36084 5908
rect 36039 5868 36084 5896
rect 36078 5856 36084 5868
rect 36136 5856 36142 5908
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5828 2835 5831
rect 2866 5828 2872 5840
rect 2823 5800 2872 5828
rect 2823 5797 2835 5800
rect 2777 5791 2835 5797
rect 2866 5788 2872 5800
rect 2924 5828 2930 5840
rect 3605 5831 3663 5837
rect 3605 5828 3617 5831
rect 2924 5800 3617 5828
rect 2924 5788 2930 5800
rect 3605 5797 3617 5800
rect 3651 5797 3663 5831
rect 3605 5791 3663 5797
rect 3970 5788 3976 5840
rect 4028 5828 4034 5840
rect 4617 5831 4675 5837
rect 4617 5828 4629 5831
rect 4028 5800 4629 5828
rect 4028 5788 4034 5800
rect 4617 5797 4629 5800
rect 4663 5828 4675 5831
rect 4982 5828 4988 5840
rect 4663 5800 4988 5828
rect 4663 5797 4675 5800
rect 4617 5791 4675 5797
rect 4982 5788 4988 5800
rect 5040 5788 5046 5840
rect 7368 5831 7426 5837
rect 7368 5797 7380 5831
rect 7414 5828 7426 5831
rect 8018 5828 8024 5840
rect 7414 5800 8024 5828
rect 7414 5797 7426 5800
rect 7368 5791 7426 5797
rect 8018 5788 8024 5800
rect 8076 5788 8082 5840
rect 10134 5788 10140 5840
rect 10192 5828 10198 5840
rect 10689 5831 10747 5837
rect 10689 5828 10701 5831
rect 10192 5800 10701 5828
rect 10192 5788 10198 5800
rect 10689 5797 10701 5800
rect 10735 5797 10747 5831
rect 10689 5791 10747 5797
rect 10778 5788 10784 5840
rect 10836 5828 10842 5840
rect 12250 5828 12256 5840
rect 10836 5800 10881 5828
rect 12211 5800 12256 5828
rect 10836 5788 10842 5800
rect 12250 5788 12256 5800
rect 12308 5788 12314 5840
rect 12526 5788 12532 5840
rect 12584 5828 12590 5840
rect 13998 5828 14004 5840
rect 12584 5800 12629 5828
rect 13959 5800 14004 5828
rect 12584 5788 12590 5800
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 14182 5828 14188 5840
rect 14143 5800 14188 5828
rect 14182 5788 14188 5800
rect 14240 5788 14246 5840
rect 14277 5831 14335 5837
rect 14277 5797 14289 5831
rect 14323 5828 14335 5831
rect 15102 5828 15108 5840
rect 14323 5800 15108 5828
rect 14323 5797 14335 5800
rect 14277 5791 14335 5797
rect 2406 5720 2412 5772
rect 2464 5760 2470 5772
rect 2593 5763 2651 5769
rect 2593 5760 2605 5763
rect 2464 5732 2605 5760
rect 2464 5720 2470 5732
rect 2593 5729 2605 5732
rect 2639 5760 2651 5763
rect 4062 5760 4068 5772
rect 2639 5732 3648 5760
rect 4023 5732 4068 5760
rect 2639 5729 2651 5732
rect 2593 5723 2651 5729
rect 2130 5652 2136 5704
rect 2188 5692 2194 5704
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 2188 5664 2881 5692
rect 2188 5652 2194 5664
rect 2869 5661 2881 5664
rect 2915 5692 2927 5695
rect 3050 5692 3056 5704
rect 2915 5664 3056 5692
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3620 5692 3648 5732
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 5626 5720 5632 5772
rect 5684 5760 5690 5772
rect 6181 5763 6239 5769
rect 6181 5760 6193 5763
rect 5684 5732 6193 5760
rect 5684 5720 5690 5732
rect 6181 5729 6193 5732
rect 6227 5760 6239 5763
rect 6549 5763 6607 5769
rect 6549 5760 6561 5763
rect 6227 5732 6561 5760
rect 6227 5729 6239 5732
rect 6181 5723 6239 5729
rect 6549 5729 6561 5732
rect 6595 5760 6607 5763
rect 7006 5760 7012 5772
rect 6595 5732 7012 5760
rect 6595 5729 6607 5732
rect 6549 5723 6607 5729
rect 7006 5720 7012 5732
rect 7064 5720 7070 5772
rect 10502 5760 10508 5772
rect 10463 5732 10508 5760
rect 10502 5720 10508 5732
rect 10560 5720 10566 5772
rect 11425 5763 11483 5769
rect 11425 5729 11437 5763
rect 11471 5760 11483 5763
rect 11974 5760 11980 5772
rect 11471 5732 11980 5760
rect 11471 5729 11483 5732
rect 11425 5723 11483 5729
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 13814 5720 13820 5772
rect 13872 5760 13878 5772
rect 14292 5760 14320 5791
rect 15102 5788 15108 5800
rect 15160 5788 15166 5840
rect 16758 5788 16764 5840
rect 16816 5828 16822 5840
rect 18046 5828 18052 5840
rect 16816 5800 16861 5828
rect 18007 5800 18052 5828
rect 16816 5788 16822 5800
rect 18046 5788 18052 5800
rect 18104 5788 18110 5840
rect 18230 5828 18236 5840
rect 18191 5800 18236 5828
rect 18230 5788 18236 5800
rect 18288 5788 18294 5840
rect 21726 5788 21732 5840
rect 21784 5828 21790 5840
rect 22462 5828 22468 5840
rect 21784 5800 22468 5828
rect 21784 5788 21790 5800
rect 22462 5788 22468 5800
rect 22520 5788 22526 5840
rect 23106 5828 23112 5840
rect 22664 5800 23112 5828
rect 13872 5732 14320 5760
rect 20717 5763 20775 5769
rect 13872 5720 13878 5732
rect 20717 5729 20729 5763
rect 20763 5760 20775 5763
rect 21450 5760 21456 5772
rect 20763 5732 21456 5760
rect 20763 5729 20775 5732
rect 20717 5723 20775 5729
rect 21450 5720 21456 5732
rect 21508 5720 21514 5772
rect 21818 5760 21824 5772
rect 21560 5732 21824 5760
rect 4522 5692 4528 5704
rect 3620 5664 4528 5692
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 5994 5692 6000 5704
rect 5955 5664 6000 5692
rect 5994 5652 6000 5664
rect 6052 5652 6058 5704
rect 6730 5652 6736 5704
rect 6788 5692 6794 5704
rect 7101 5695 7159 5701
rect 7101 5692 7113 5695
rect 6788 5664 7113 5692
rect 6788 5652 6794 5664
rect 7101 5661 7113 5664
rect 7147 5661 7159 5695
rect 7101 5655 7159 5661
rect 16390 5652 16396 5704
rect 16448 5692 16454 5704
rect 16669 5695 16727 5701
rect 16669 5692 16681 5695
rect 16448 5664 16681 5692
rect 16448 5652 16454 5664
rect 16669 5661 16681 5664
rect 16715 5692 16727 5695
rect 16850 5692 16856 5704
rect 16715 5664 16856 5692
rect 16715 5661 16727 5664
rect 16669 5655 16727 5661
rect 16850 5652 16856 5664
rect 16908 5652 16914 5704
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5661 18383 5695
rect 19794 5692 19800 5704
rect 19755 5664 19800 5692
rect 18325 5655 18383 5661
rect 5629 5627 5687 5633
rect 5629 5593 5641 5627
rect 5675 5624 5687 5627
rect 6822 5624 6828 5636
rect 5675 5596 6828 5624
rect 5675 5593 5687 5596
rect 5629 5587 5687 5593
rect 6822 5584 6828 5596
rect 6880 5584 6886 5636
rect 13722 5624 13728 5636
rect 13683 5596 13728 5624
rect 13722 5584 13728 5596
rect 13780 5584 13786 5636
rect 1673 5559 1731 5565
rect 1673 5525 1685 5559
rect 1719 5556 1731 5559
rect 1762 5556 1768 5568
rect 1719 5528 1768 5556
rect 1719 5525 1731 5528
rect 1673 5519 1731 5525
rect 1762 5516 1768 5528
rect 1820 5516 1826 5568
rect 2130 5556 2136 5568
rect 2091 5528 2136 5556
rect 2130 5516 2136 5528
rect 2188 5516 2194 5568
rect 2317 5559 2375 5565
rect 2317 5525 2329 5559
rect 2363 5556 2375 5559
rect 2682 5556 2688 5568
rect 2363 5528 2688 5556
rect 2363 5525 2375 5528
rect 2317 5519 2375 5525
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 3142 5516 3148 5568
rect 3200 5556 3206 5568
rect 3237 5559 3295 5565
rect 3237 5556 3249 5559
rect 3200 5528 3249 5556
rect 3200 5516 3206 5528
rect 3237 5525 3249 5528
rect 3283 5525 3295 5559
rect 3237 5519 3295 5525
rect 4890 5516 4896 5568
rect 4948 5556 4954 5568
rect 4985 5559 5043 5565
rect 4985 5556 4997 5559
rect 4948 5528 4997 5556
rect 4948 5516 4954 5528
rect 4985 5525 4997 5528
rect 5031 5525 5043 5559
rect 4985 5519 5043 5525
rect 8481 5559 8539 5565
rect 8481 5525 8493 5559
rect 8527 5556 8539 5559
rect 9490 5556 9496 5568
rect 8527 5528 9496 5556
rect 8527 5525 8539 5528
rect 8481 5519 8539 5525
rect 9490 5516 9496 5528
rect 9548 5516 9554 5568
rect 10226 5556 10232 5568
rect 10187 5528 10232 5556
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 16206 5556 16212 5568
rect 16167 5528 16212 5556
rect 16206 5516 16212 5528
rect 16264 5516 16270 5568
rect 16574 5516 16580 5568
rect 16632 5556 16638 5568
rect 17773 5559 17831 5565
rect 17773 5556 17785 5559
rect 16632 5528 17785 5556
rect 16632 5516 16638 5528
rect 17773 5525 17785 5528
rect 17819 5525 17831 5559
rect 18340 5556 18368 5655
rect 19794 5652 19800 5664
rect 19852 5652 19858 5704
rect 20806 5652 20812 5704
rect 20864 5692 20870 5704
rect 21560 5701 21588 5732
rect 21818 5720 21824 5732
rect 21876 5720 21882 5772
rect 22002 5720 22008 5772
rect 22060 5760 22066 5772
rect 22664 5769 22692 5800
rect 23106 5788 23112 5800
rect 23164 5788 23170 5840
rect 28997 5831 29055 5837
rect 28997 5797 29009 5831
rect 29043 5828 29055 5831
rect 29178 5828 29184 5840
rect 29043 5800 29184 5828
rect 29043 5797 29055 5800
rect 28997 5791 29055 5797
rect 29178 5788 29184 5800
rect 29236 5788 29242 5840
rect 29362 5788 29368 5840
rect 29420 5828 29426 5840
rect 29457 5831 29515 5837
rect 29457 5828 29469 5831
rect 29420 5800 29469 5828
rect 29420 5788 29426 5800
rect 29457 5797 29469 5800
rect 29503 5797 29515 5831
rect 29457 5791 29515 5797
rect 32493 5831 32551 5837
rect 32493 5797 32505 5831
rect 32539 5828 32551 5831
rect 32953 5831 33011 5837
rect 32953 5828 32965 5831
rect 32539 5800 32965 5828
rect 32539 5797 32551 5800
rect 32493 5791 32551 5797
rect 32953 5797 32965 5800
rect 32999 5828 33011 5831
rect 33042 5828 33048 5840
rect 32999 5800 33048 5828
rect 32999 5797 33011 5800
rect 32953 5791 33011 5797
rect 33042 5788 33048 5800
rect 33100 5788 33106 5840
rect 33226 5828 33232 5840
rect 33187 5800 33232 5828
rect 33226 5788 33232 5800
rect 33284 5788 33290 5840
rect 33686 5828 33692 5840
rect 33647 5800 33692 5828
rect 33686 5788 33692 5800
rect 33744 5788 33750 5840
rect 34146 5788 34152 5840
rect 34204 5828 34210 5840
rect 34394 5831 34452 5837
rect 34394 5828 34406 5831
rect 34204 5800 34406 5828
rect 34204 5788 34210 5800
rect 34394 5797 34406 5800
rect 34440 5797 34452 5831
rect 34394 5791 34452 5797
rect 22922 5769 22928 5772
rect 22649 5763 22707 5769
rect 22649 5760 22661 5763
rect 22060 5732 22661 5760
rect 22060 5720 22066 5732
rect 22649 5729 22661 5732
rect 22695 5729 22707 5763
rect 22916 5760 22928 5769
rect 22883 5732 22928 5760
rect 22649 5723 22707 5729
rect 22916 5723 22928 5732
rect 22922 5720 22928 5723
rect 22980 5720 22986 5772
rect 26970 5720 26976 5772
rect 27028 5760 27034 5772
rect 27525 5763 27583 5769
rect 27525 5760 27537 5763
rect 27028 5732 27537 5760
rect 27028 5720 27034 5732
rect 27525 5729 27537 5732
rect 27571 5760 27583 5763
rect 27706 5760 27712 5772
rect 27571 5732 27712 5760
rect 27571 5729 27583 5732
rect 27525 5723 27583 5729
rect 27706 5720 27712 5732
rect 27764 5760 27770 5772
rect 27893 5763 27951 5769
rect 27893 5760 27905 5763
rect 27764 5732 27905 5760
rect 27764 5720 27770 5732
rect 27893 5729 27905 5732
rect 27939 5729 27951 5763
rect 27893 5723 27951 5729
rect 28442 5720 28448 5772
rect 28500 5760 28506 5772
rect 28813 5763 28871 5769
rect 28813 5760 28825 5763
rect 28500 5732 28825 5760
rect 28500 5720 28506 5732
rect 28813 5729 28825 5732
rect 28859 5729 28871 5763
rect 30653 5763 30711 5769
rect 30653 5760 30665 5763
rect 28813 5723 28871 5729
rect 29104 5732 30665 5760
rect 21545 5695 21603 5701
rect 21545 5692 21557 5695
rect 20864 5664 21557 5692
rect 20864 5652 20870 5664
rect 21545 5661 21557 5664
rect 21591 5661 21603 5695
rect 21545 5655 21603 5661
rect 24854 5652 24860 5704
rect 24912 5692 24918 5704
rect 25225 5695 25283 5701
rect 25225 5692 25237 5695
rect 24912 5664 25237 5692
rect 24912 5652 24918 5664
rect 25225 5661 25237 5664
rect 25271 5661 25283 5695
rect 27430 5692 27436 5704
rect 27343 5664 27436 5692
rect 25225 5655 25283 5661
rect 27430 5652 27436 5664
rect 27488 5692 27494 5704
rect 28166 5692 28172 5704
rect 27488 5664 28172 5692
rect 27488 5652 27494 5664
rect 28166 5652 28172 5664
rect 28224 5652 28230 5704
rect 28994 5652 29000 5704
rect 29052 5692 29058 5704
rect 29104 5701 29132 5732
rect 30653 5729 30665 5732
rect 30699 5760 30711 5763
rect 30742 5760 30748 5772
rect 30699 5732 30748 5760
rect 30699 5729 30711 5732
rect 30653 5723 30711 5729
rect 30742 5720 30748 5732
rect 30800 5760 30806 5772
rect 31021 5763 31079 5769
rect 31021 5760 31033 5763
rect 30800 5732 31033 5760
rect 30800 5720 30806 5732
rect 31021 5729 31033 5732
rect 31067 5729 31079 5763
rect 31021 5723 31079 5729
rect 29089 5695 29147 5701
rect 29089 5692 29101 5695
rect 29052 5664 29101 5692
rect 29052 5652 29058 5664
rect 29089 5661 29101 5664
rect 29135 5661 29147 5695
rect 30466 5692 30472 5704
rect 30427 5664 30472 5692
rect 29089 5655 29147 5661
rect 30466 5652 30472 5664
rect 30524 5652 30530 5704
rect 34054 5652 34060 5704
rect 34112 5692 34118 5704
rect 34149 5695 34207 5701
rect 34149 5692 34161 5695
rect 34112 5664 34161 5692
rect 34112 5652 34118 5664
rect 34149 5661 34161 5664
rect 34195 5661 34207 5695
rect 34149 5655 34207 5661
rect 20714 5584 20720 5636
rect 20772 5624 20778 5636
rect 21177 5627 21235 5633
rect 21177 5624 21189 5627
rect 20772 5596 21189 5624
rect 20772 5584 20778 5596
rect 21177 5593 21189 5596
rect 21223 5593 21235 5627
rect 26050 5624 26056 5636
rect 25963 5596 26056 5624
rect 21177 5587 21235 5593
rect 26050 5584 26056 5596
rect 26108 5624 26114 5636
rect 26973 5627 27031 5633
rect 26973 5624 26985 5627
rect 26108 5596 26985 5624
rect 26108 5584 26114 5596
rect 26973 5593 26985 5596
rect 27019 5593 27031 5627
rect 26973 5587 27031 5593
rect 31846 5584 31852 5636
rect 31904 5624 31910 5636
rect 32677 5627 32735 5633
rect 32677 5624 32689 5627
rect 31904 5596 32689 5624
rect 31904 5584 31910 5596
rect 32677 5593 32689 5596
rect 32723 5593 32735 5627
rect 32677 5587 32735 5593
rect 35894 5584 35900 5636
rect 35952 5624 35958 5636
rect 36354 5624 36360 5636
rect 35952 5596 36360 5624
rect 35952 5584 35958 5596
rect 36354 5584 36360 5596
rect 36412 5624 36418 5636
rect 36449 5627 36507 5633
rect 36449 5624 36461 5627
rect 36412 5596 36461 5624
rect 36412 5584 36418 5596
rect 36449 5593 36461 5596
rect 36495 5593 36507 5627
rect 36449 5587 36507 5593
rect 18690 5556 18696 5568
rect 18340 5528 18696 5556
rect 17773 5519 17831 5525
rect 18690 5516 18696 5528
rect 18748 5516 18754 5568
rect 24029 5559 24087 5565
rect 24029 5525 24041 5559
rect 24075 5556 24087 5559
rect 24302 5556 24308 5568
rect 24075 5528 24308 5556
rect 24075 5525 24087 5528
rect 24029 5519 24087 5525
rect 24302 5516 24308 5528
rect 24360 5516 24366 5568
rect 25682 5556 25688 5568
rect 25595 5528 25688 5556
rect 25682 5516 25688 5528
rect 25740 5556 25746 5568
rect 26142 5556 26148 5568
rect 25740 5528 26148 5556
rect 25740 5516 25746 5528
rect 26142 5516 26148 5528
rect 26200 5516 26206 5568
rect 30098 5556 30104 5568
rect 30059 5528 30104 5556
rect 30098 5516 30104 5528
rect 30156 5516 30162 5568
rect 1104 5466 38824 5488
rect 1104 5414 7648 5466
rect 7700 5414 7712 5466
rect 7764 5414 7776 5466
rect 7828 5414 7840 5466
rect 7892 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 34315 5466
rect 34367 5414 34379 5466
rect 34431 5414 34443 5466
rect 34495 5414 34507 5466
rect 34559 5414 38824 5466
rect 1104 5392 38824 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 1670 5352 1676 5364
rect 1627 5324 1676 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 1670 5312 1676 5324
rect 1728 5312 1734 5364
rect 2222 5312 2228 5364
rect 2280 5352 2286 5364
rect 2317 5355 2375 5361
rect 2317 5352 2329 5355
rect 2280 5324 2329 5352
rect 2280 5312 2286 5324
rect 2317 5321 2329 5324
rect 2363 5352 2375 5355
rect 2406 5352 2412 5364
rect 2363 5324 2412 5352
rect 2363 5321 2375 5324
rect 2317 5315 2375 5321
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 2866 5352 2872 5364
rect 2827 5324 2872 5352
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 4338 5312 4344 5364
rect 4396 5352 4402 5364
rect 4433 5355 4491 5361
rect 4433 5352 4445 5355
rect 4396 5324 4445 5352
rect 4396 5312 4402 5324
rect 4433 5321 4445 5324
rect 4479 5321 4491 5355
rect 5626 5352 5632 5364
rect 5587 5324 5632 5352
rect 4433 5315 4491 5321
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 6546 5352 6552 5364
rect 6507 5324 6552 5352
rect 6546 5312 6552 5324
rect 6604 5352 6610 5364
rect 10870 5352 10876 5364
rect 6604 5324 7788 5352
rect 10831 5324 10876 5352
rect 6604 5312 6610 5324
rect 6181 5287 6239 5293
rect 6181 5253 6193 5287
rect 6227 5284 6239 5287
rect 6730 5284 6736 5296
rect 6227 5256 6736 5284
rect 6227 5253 6239 5256
rect 6181 5247 6239 5253
rect 6730 5244 6736 5256
rect 6788 5244 6794 5296
rect 7374 5284 7380 5296
rect 7335 5256 7380 5284
rect 7374 5244 7380 5256
rect 7432 5244 7438 5296
rect 4982 5216 4988 5228
rect 4943 5188 4988 5216
rect 4982 5176 4988 5188
rect 5040 5176 5046 5228
rect 7760 5225 7788 5324
rect 10870 5312 10876 5324
rect 10928 5312 10934 5364
rect 11977 5355 12035 5361
rect 11977 5321 11989 5355
rect 12023 5352 12035 5355
rect 12250 5352 12256 5364
rect 12023 5324 12256 5352
rect 12023 5321 12035 5324
rect 11977 5315 12035 5321
rect 12250 5312 12256 5324
rect 12308 5312 12314 5364
rect 12526 5312 12532 5364
rect 12584 5352 12590 5364
rect 12897 5355 12955 5361
rect 12897 5352 12909 5355
rect 12584 5324 12909 5352
rect 12584 5312 12590 5324
rect 12897 5321 12909 5324
rect 12943 5321 12955 5355
rect 13722 5352 13728 5364
rect 13683 5324 13728 5352
rect 12897 5315 12955 5321
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 14093 5355 14151 5361
rect 14093 5321 14105 5355
rect 14139 5352 14151 5355
rect 14182 5352 14188 5364
rect 14139 5324 14188 5352
rect 14139 5321 14151 5324
rect 14093 5315 14151 5321
rect 14182 5312 14188 5324
rect 14240 5352 14246 5364
rect 15749 5355 15807 5361
rect 15749 5352 15761 5355
rect 14240 5324 15761 5352
rect 14240 5312 14246 5324
rect 15749 5321 15761 5324
rect 15795 5321 15807 5355
rect 15749 5315 15807 5321
rect 16758 5312 16764 5364
rect 16816 5352 16822 5364
rect 17037 5355 17095 5361
rect 17037 5352 17049 5355
rect 16816 5324 17049 5352
rect 16816 5312 16822 5324
rect 17037 5321 17049 5324
rect 17083 5321 17095 5355
rect 17402 5352 17408 5364
rect 17363 5324 17408 5352
rect 17037 5315 17095 5321
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 17770 5352 17776 5364
rect 17731 5324 17776 5352
rect 17770 5312 17776 5324
rect 17828 5312 17834 5364
rect 19518 5352 19524 5364
rect 19479 5324 19524 5352
rect 19518 5312 19524 5324
rect 19576 5312 19582 5364
rect 20806 5352 20812 5364
rect 20767 5324 20812 5352
rect 20806 5312 20812 5324
rect 20864 5312 20870 5364
rect 21085 5355 21143 5361
rect 21085 5321 21097 5355
rect 21131 5352 21143 5355
rect 21542 5352 21548 5364
rect 21131 5324 21548 5352
rect 21131 5321 21143 5324
rect 21085 5315 21143 5321
rect 21542 5312 21548 5324
rect 21600 5312 21606 5364
rect 22373 5355 22431 5361
rect 22373 5321 22385 5355
rect 22419 5352 22431 5355
rect 22462 5352 22468 5364
rect 22419 5324 22468 5352
rect 22419 5321 22431 5324
rect 22373 5315 22431 5321
rect 22462 5312 22468 5324
rect 22520 5312 22526 5364
rect 22741 5355 22799 5361
rect 22741 5321 22753 5355
rect 22787 5352 22799 5355
rect 23106 5352 23112 5364
rect 22787 5324 23112 5352
rect 22787 5321 22799 5324
rect 22741 5315 22799 5321
rect 23106 5312 23112 5324
rect 23164 5312 23170 5364
rect 23198 5312 23204 5364
rect 23256 5352 23262 5364
rect 23256 5324 24440 5352
rect 23256 5312 23262 5324
rect 8941 5287 8999 5293
rect 8941 5253 8953 5287
rect 8987 5284 8999 5287
rect 9398 5284 9404 5296
rect 8987 5256 9404 5284
rect 8987 5253 8999 5256
rect 8941 5247 8999 5253
rect 9398 5244 9404 5256
rect 9456 5244 9462 5296
rect 10229 5287 10287 5293
rect 10229 5253 10241 5287
rect 10275 5284 10287 5287
rect 10778 5284 10784 5296
rect 10275 5256 10784 5284
rect 10275 5253 10287 5256
rect 10229 5247 10287 5253
rect 10778 5244 10784 5256
rect 10836 5244 10842 5296
rect 13998 5244 14004 5296
rect 14056 5284 14062 5296
rect 14369 5287 14427 5293
rect 14369 5284 14381 5287
rect 14056 5256 14381 5284
rect 14056 5244 14062 5256
rect 14369 5253 14381 5256
rect 14415 5253 14427 5287
rect 14369 5247 14427 5253
rect 15565 5287 15623 5293
rect 15565 5253 15577 5287
rect 15611 5284 15623 5287
rect 16390 5284 16396 5296
rect 15611 5256 16396 5284
rect 15611 5253 15623 5256
rect 15565 5247 15623 5253
rect 16390 5244 16396 5256
rect 16448 5244 16454 5296
rect 7745 5219 7803 5225
rect 7745 5185 7757 5219
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 10689 5219 10747 5225
rect 10689 5185 10701 5219
rect 10735 5216 10747 5219
rect 11422 5216 11428 5228
rect 10735 5188 11428 5216
rect 10735 5185 10747 5188
rect 10689 5179 10747 5185
rect 11422 5176 11428 5188
rect 11480 5176 11486 5228
rect 12437 5219 12495 5225
rect 12437 5185 12449 5219
rect 12483 5216 12495 5219
rect 13354 5216 13360 5228
rect 12483 5188 13360 5216
rect 12483 5185 12495 5188
rect 12437 5179 12495 5185
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 14829 5219 14887 5225
rect 14829 5185 14841 5219
rect 14875 5216 14887 5219
rect 15838 5216 15844 5228
rect 14875 5188 15844 5216
rect 14875 5185 14887 5188
rect 14829 5179 14887 5185
rect 15838 5176 15844 5188
rect 15896 5216 15902 5228
rect 16117 5219 16175 5225
rect 16117 5216 16129 5219
rect 15896 5188 16129 5216
rect 15896 5176 15902 5188
rect 16117 5185 16129 5188
rect 16163 5185 16175 5219
rect 16117 5179 16175 5185
rect 16761 5219 16819 5225
rect 16761 5185 16773 5219
rect 16807 5216 16819 5219
rect 17310 5216 17316 5228
rect 16807 5188 17316 5216
rect 16807 5185 16819 5188
rect 16761 5179 16819 5185
rect 17310 5176 17316 5188
rect 17368 5176 17374 5228
rect 17788 5216 17816 5312
rect 18138 5284 18144 5296
rect 18099 5256 18144 5284
rect 18138 5244 18144 5256
rect 18196 5244 18202 5296
rect 19797 5287 19855 5293
rect 19797 5253 19809 5287
rect 19843 5284 19855 5287
rect 20346 5284 20352 5296
rect 19843 5256 20352 5284
rect 19843 5253 19855 5256
rect 19797 5247 19855 5253
rect 20346 5244 20352 5256
rect 20404 5284 20410 5296
rect 21174 5284 21180 5296
rect 20404 5256 21180 5284
rect 20404 5244 20410 5256
rect 21174 5244 21180 5256
rect 21232 5244 21238 5296
rect 21358 5284 21364 5296
rect 21319 5256 21364 5284
rect 21358 5244 21364 5256
rect 21416 5244 21422 5296
rect 21818 5244 21824 5296
rect 21876 5284 21882 5296
rect 23753 5287 23811 5293
rect 23753 5284 23765 5287
rect 21876 5256 23765 5284
rect 21876 5244 21882 5256
rect 23753 5253 23765 5256
rect 23799 5253 23811 5287
rect 24412 5284 24440 5324
rect 24486 5312 24492 5364
rect 24544 5352 24550 5364
rect 24673 5355 24731 5361
rect 24673 5352 24685 5355
rect 24544 5324 24685 5352
rect 24544 5312 24550 5324
rect 24673 5321 24685 5324
rect 24719 5321 24731 5355
rect 25590 5352 25596 5364
rect 25551 5324 25596 5352
rect 24673 5315 24731 5321
rect 25590 5312 25596 5324
rect 25648 5312 25654 5364
rect 26602 5352 26608 5364
rect 26515 5324 26608 5352
rect 26602 5312 26608 5324
rect 26660 5352 26666 5364
rect 27338 5352 27344 5364
rect 26660 5324 27344 5352
rect 26660 5312 26666 5324
rect 27338 5312 27344 5324
rect 27396 5312 27402 5364
rect 28166 5352 28172 5364
rect 28127 5324 28172 5352
rect 28166 5312 28172 5324
rect 28224 5312 28230 5364
rect 30374 5312 30380 5364
rect 30432 5352 30438 5364
rect 30926 5352 30932 5364
rect 30432 5324 30932 5352
rect 30432 5312 30438 5324
rect 30926 5312 30932 5324
rect 30984 5312 30990 5364
rect 31849 5355 31907 5361
rect 31849 5321 31861 5355
rect 31895 5352 31907 5355
rect 33042 5352 33048 5364
rect 31895 5324 33048 5352
rect 31895 5321 31907 5324
rect 31849 5315 31907 5321
rect 33042 5312 33048 5324
rect 33100 5312 33106 5364
rect 35618 5352 35624 5364
rect 35579 5324 35624 5352
rect 35618 5312 35624 5324
rect 35676 5312 35682 5364
rect 26789 5287 26847 5293
rect 26789 5284 26801 5287
rect 24412 5256 26801 5284
rect 23753 5247 23811 5253
rect 26789 5253 26801 5256
rect 26835 5284 26847 5287
rect 26881 5287 26939 5293
rect 26881 5284 26893 5287
rect 26835 5256 26893 5284
rect 26835 5253 26847 5256
rect 26789 5247 26847 5253
rect 26881 5253 26893 5256
rect 26927 5253 26939 5287
rect 26881 5247 26939 5253
rect 27157 5287 27215 5293
rect 27157 5253 27169 5287
rect 27203 5253 27215 5287
rect 27157 5247 27215 5253
rect 29641 5287 29699 5293
rect 29641 5253 29653 5287
rect 29687 5284 29699 5287
rect 30282 5284 30288 5296
rect 29687 5256 30288 5284
rect 29687 5253 29699 5256
rect 29641 5247 29699 5253
rect 18506 5216 18512 5228
rect 17788 5188 18512 5216
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 24210 5216 24216 5228
rect 24123 5188 24216 5216
rect 24210 5176 24216 5188
rect 24268 5216 24274 5228
rect 24762 5216 24768 5228
rect 24268 5188 24768 5216
rect 24268 5176 24274 5188
rect 24762 5176 24768 5188
rect 24820 5176 24826 5228
rect 26050 5216 26056 5228
rect 26011 5188 26056 5216
rect 26050 5176 26056 5188
rect 26108 5176 26114 5228
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 1670 5148 1676 5160
rect 1443 5120 1676 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 1670 5108 1676 5120
rect 1728 5148 1734 5160
rect 3142 5148 3148 5160
rect 1728 5120 3148 5148
rect 1728 5108 1734 5120
rect 3142 5108 3148 5120
rect 3200 5108 3206 5160
rect 4154 5148 4160 5160
rect 4067 5120 4160 5148
rect 4154 5108 4160 5120
rect 4212 5148 4218 5160
rect 5074 5148 5080 5160
rect 4212 5120 5080 5148
rect 4212 5108 4218 5120
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 9493 5151 9551 5157
rect 9493 5148 9505 5151
rect 8312 5120 9505 5148
rect 3418 5080 3424 5092
rect 3379 5052 3424 5080
rect 3418 5040 3424 5052
rect 3476 5040 3482 5092
rect 3878 5040 3884 5092
rect 3936 5080 3942 5092
rect 4709 5083 4767 5089
rect 4709 5080 4721 5083
rect 3936 5052 4721 5080
rect 3936 5040 3942 5052
rect 4709 5049 4721 5052
rect 4755 5049 4767 5083
rect 7926 5080 7932 5092
rect 7887 5052 7932 5080
rect 4709 5043 4767 5049
rect 7926 5040 7932 5052
rect 7984 5080 7990 5092
rect 8312 5089 8340 5120
rect 9493 5117 9505 5120
rect 9539 5117 9551 5151
rect 9493 5111 9551 5117
rect 11054 5108 11060 5160
rect 11112 5148 11118 5160
rect 11149 5151 11207 5157
rect 11149 5148 11161 5151
rect 11112 5120 11161 5148
rect 11112 5108 11118 5120
rect 11149 5117 11161 5120
rect 11195 5117 11207 5151
rect 11149 5111 11207 5117
rect 15197 5151 15255 5157
rect 15197 5117 15209 5151
rect 15243 5148 15255 5151
rect 19245 5151 19303 5157
rect 15243 5120 16252 5148
rect 15243 5117 15255 5120
rect 15197 5111 15255 5117
rect 16224 5092 16252 5120
rect 19245 5117 19257 5151
rect 19291 5148 19303 5151
rect 19794 5148 19800 5160
rect 19291 5120 19800 5148
rect 19291 5117 19303 5120
rect 19245 5111 19303 5117
rect 19794 5108 19800 5120
rect 19852 5148 19858 5160
rect 20073 5151 20131 5157
rect 20073 5148 20085 5151
rect 19852 5120 20085 5148
rect 19852 5108 19858 5120
rect 20073 5117 20085 5120
rect 20119 5117 20131 5151
rect 20073 5111 20131 5117
rect 20254 5108 20260 5160
rect 20312 5148 20318 5160
rect 20349 5151 20407 5157
rect 20349 5148 20361 5151
rect 20312 5120 20361 5148
rect 20312 5108 20318 5120
rect 20349 5117 20361 5120
rect 20395 5117 20407 5151
rect 20349 5111 20407 5117
rect 21450 5108 21456 5160
rect 21508 5148 21514 5160
rect 21637 5151 21695 5157
rect 21637 5148 21649 5151
rect 21508 5120 21649 5148
rect 21508 5108 21514 5120
rect 21637 5117 21649 5120
rect 21683 5117 21695 5151
rect 21637 5111 21695 5117
rect 23477 5151 23535 5157
rect 23477 5117 23489 5151
rect 23523 5148 23535 5151
rect 27172 5148 27200 5247
rect 30282 5244 30288 5256
rect 30340 5244 30346 5296
rect 27706 5216 27712 5228
rect 27667 5188 27712 5216
rect 27706 5176 27712 5188
rect 27764 5176 27770 5228
rect 29914 5176 29920 5228
rect 29972 5216 29978 5228
rect 30193 5219 30251 5225
rect 30193 5216 30205 5219
rect 29972 5188 30205 5216
rect 29972 5176 29978 5188
rect 30193 5185 30205 5188
rect 30239 5216 30251 5219
rect 32122 5216 32128 5228
rect 30239 5188 32128 5216
rect 30239 5185 30251 5188
rect 30193 5179 30251 5185
rect 32122 5176 32128 5188
rect 32180 5216 32186 5228
rect 32180 5188 32444 5216
rect 32180 5176 32186 5188
rect 28626 5148 28632 5160
rect 23523 5120 24348 5148
rect 23523 5117 23535 5120
rect 23477 5111 23535 5117
rect 24320 5092 24348 5120
rect 26068 5120 27200 5148
rect 27264 5120 28632 5148
rect 8297 5083 8355 5089
rect 8297 5080 8309 5083
rect 7984 5052 8309 5080
rect 7984 5040 7990 5052
rect 8297 5049 8309 5052
rect 8343 5049 8355 5083
rect 8297 5043 8355 5049
rect 8938 5040 8944 5092
rect 8996 5080 9002 5092
rect 9217 5083 9275 5089
rect 9217 5080 9229 5083
rect 8996 5052 9229 5080
rect 8996 5040 9002 5052
rect 9217 5049 9229 5052
rect 9263 5049 9275 5083
rect 9217 5043 9275 5049
rect 9401 5083 9459 5089
rect 9401 5049 9413 5083
rect 9447 5080 9459 5083
rect 9582 5080 9588 5092
rect 9447 5052 9588 5080
rect 9447 5049 9459 5052
rect 9401 5043 9459 5049
rect 2685 5015 2743 5021
rect 2685 4981 2697 5015
rect 2731 5012 2743 5015
rect 3142 5012 3148 5024
rect 2731 4984 3148 5012
rect 2731 4981 2743 4984
rect 2685 4975 2743 4981
rect 3142 4972 3148 4984
rect 3200 5012 3206 5024
rect 3329 5015 3387 5021
rect 3329 5012 3341 5015
rect 3200 4984 3341 5012
rect 3200 4972 3206 4984
rect 3329 4981 3341 4984
rect 3375 5012 3387 5015
rect 3510 5012 3516 5024
rect 3375 4984 3516 5012
rect 3375 4981 3387 4984
rect 3329 4975 3387 4981
rect 3510 4972 3516 4984
rect 3568 4972 3574 5024
rect 4890 5012 4896 5024
rect 4851 4984 4896 5012
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 6822 4972 6828 5024
rect 6880 5012 6886 5024
rect 7101 5015 7159 5021
rect 7101 5012 7113 5015
rect 6880 4984 7113 5012
rect 6880 4972 6886 4984
rect 7101 4981 7113 4984
rect 7147 5012 7159 5015
rect 7282 5012 7288 5024
rect 7147 4984 7288 5012
rect 7147 4981 7159 4984
rect 7101 4975 7159 4981
rect 7282 4972 7288 4984
rect 7340 5012 7346 5024
rect 7837 5015 7895 5021
rect 7837 5012 7849 5015
rect 7340 4984 7849 5012
rect 7340 4972 7346 4984
rect 7837 4981 7849 4984
rect 7883 4981 7895 5015
rect 8754 5012 8760 5024
rect 8667 4984 8760 5012
rect 7837 4975 7895 4981
rect 8754 4972 8760 4984
rect 8812 5012 8818 5024
rect 9416 5012 9444 5043
rect 9582 5040 9588 5052
rect 9640 5040 9646 5092
rect 16206 5080 16212 5092
rect 16167 5052 16212 5080
rect 16206 5040 16212 5052
rect 16264 5040 16270 5092
rect 16301 5083 16359 5089
rect 16301 5049 16313 5083
rect 16347 5049 16359 5083
rect 18598 5080 18604 5092
rect 18559 5052 18604 5080
rect 16301 5043 16359 5049
rect 8812 4984 9444 5012
rect 8812 4972 8818 4984
rect 10870 4972 10876 5024
rect 10928 5012 10934 5024
rect 11333 5015 11391 5021
rect 11333 5012 11345 5015
rect 10928 4984 11345 5012
rect 10928 4972 10934 4984
rect 11333 4981 11345 4984
rect 11379 4981 11391 5015
rect 11333 4975 11391 4981
rect 16114 4972 16120 5024
rect 16172 5012 16178 5024
rect 16316 5012 16344 5043
rect 18598 5040 18604 5052
rect 18656 5040 18662 5092
rect 18690 5040 18696 5092
rect 18748 5080 18754 5092
rect 21910 5080 21916 5092
rect 18748 5052 18793 5080
rect 21871 5052 21916 5080
rect 18748 5040 18754 5052
rect 21910 5040 21916 5052
rect 21968 5040 21974 5092
rect 24302 5080 24308 5092
rect 24263 5052 24308 5080
rect 24302 5040 24308 5052
rect 24360 5040 24366 5092
rect 25866 5040 25872 5092
rect 25924 5080 25930 5092
rect 26068 5089 26096 5120
rect 26053 5083 26111 5089
rect 26053 5080 26065 5083
rect 25924 5052 26065 5080
rect 25924 5040 25930 5052
rect 26053 5049 26065 5052
rect 26099 5049 26111 5083
rect 26053 5043 26111 5049
rect 26145 5083 26203 5089
rect 26145 5049 26157 5083
rect 26191 5080 26203 5083
rect 27264 5080 27292 5120
rect 28626 5108 28632 5120
rect 28684 5148 28690 5160
rect 28813 5151 28871 5157
rect 28813 5148 28825 5151
rect 28684 5120 28825 5148
rect 28684 5108 28690 5120
rect 28813 5117 28825 5120
rect 28859 5148 28871 5151
rect 28994 5148 29000 5160
rect 28859 5120 29000 5148
rect 28859 5117 28871 5120
rect 28813 5111 28871 5117
rect 28994 5108 29000 5120
rect 29052 5108 29058 5160
rect 31297 5151 31355 5157
rect 31297 5148 31309 5151
rect 30116 5120 31309 5148
rect 30116 5092 30144 5120
rect 31297 5117 31309 5120
rect 31343 5117 31355 5151
rect 31297 5111 31355 5117
rect 32217 5151 32275 5157
rect 32217 5117 32229 5151
rect 32263 5148 32275 5151
rect 32309 5151 32367 5157
rect 32309 5148 32321 5151
rect 32263 5120 32321 5148
rect 32263 5117 32275 5120
rect 32217 5111 32275 5117
rect 32309 5117 32321 5120
rect 32355 5117 32367 5151
rect 32416 5148 32444 5188
rect 32565 5151 32623 5157
rect 32565 5148 32577 5151
rect 32416 5120 32577 5148
rect 32309 5111 32367 5117
rect 32565 5117 32577 5120
rect 32611 5117 32623 5151
rect 34054 5148 34060 5160
rect 32565 5111 32623 5117
rect 32692 5120 34060 5148
rect 26191 5052 27292 5080
rect 26191 5049 26203 5052
rect 26145 5043 26203 5049
rect 16172 4984 16344 5012
rect 16172 4972 16178 4984
rect 19518 4972 19524 5024
rect 19576 5012 19582 5024
rect 20257 5015 20315 5021
rect 20257 5012 20269 5015
rect 19576 4984 20269 5012
rect 19576 4972 19582 4984
rect 20257 4981 20269 4984
rect 20303 5012 20315 5015
rect 20438 5012 20444 5024
rect 20303 4984 20444 5012
rect 20303 4981 20315 4984
rect 20257 4975 20315 4981
rect 20438 4972 20444 4984
rect 20496 4972 20502 5024
rect 21818 5012 21824 5024
rect 21779 4984 21824 5012
rect 21818 4972 21824 4984
rect 21876 4972 21882 5024
rect 23106 5012 23112 5024
rect 23067 4984 23112 5012
rect 23106 4972 23112 4984
rect 23164 4972 23170 5024
rect 24118 4972 24124 5024
rect 24176 5012 24182 5024
rect 24213 5015 24271 5021
rect 24213 5012 24225 5015
rect 24176 4984 24225 5012
rect 24176 4972 24182 4984
rect 24213 4981 24225 4984
rect 24259 4981 24271 5015
rect 24213 4975 24271 4981
rect 25409 5015 25467 5021
rect 25409 4981 25421 5015
rect 25455 5012 25467 5015
rect 26160 5012 26188 5043
rect 27338 5040 27344 5092
rect 27396 5080 27402 5092
rect 27433 5083 27491 5089
rect 27433 5080 27445 5083
rect 27396 5052 27445 5080
rect 27396 5040 27402 5052
rect 27433 5049 27445 5052
rect 27479 5049 27491 5083
rect 28442 5080 28448 5092
rect 28403 5052 28448 5080
rect 27433 5043 27491 5049
rect 28442 5040 28448 5052
rect 28500 5040 28506 5092
rect 29914 5080 29920 5092
rect 29875 5052 29920 5080
rect 29914 5040 29920 5052
rect 29972 5040 29978 5092
rect 30098 5080 30104 5092
rect 30059 5052 30104 5080
rect 30098 5040 30104 5052
rect 30156 5040 30162 5092
rect 32324 5080 32352 5111
rect 32692 5080 32720 5120
rect 34054 5108 34060 5120
rect 34112 5108 34118 5160
rect 35434 5148 35440 5160
rect 35395 5120 35440 5148
rect 35434 5108 35440 5120
rect 35492 5148 35498 5160
rect 35989 5151 36047 5157
rect 35989 5148 36001 5151
rect 35492 5120 36001 5148
rect 35492 5108 35498 5120
rect 35989 5117 36001 5120
rect 36035 5117 36047 5151
rect 35989 5111 36047 5117
rect 34146 5080 34152 5092
rect 32324 5052 32720 5080
rect 33704 5052 34152 5080
rect 33704 5024 33732 5052
rect 34146 5040 34152 5052
rect 34204 5080 34210 5092
rect 34609 5083 34667 5089
rect 34609 5080 34621 5083
rect 34204 5052 34621 5080
rect 34204 5040 34210 5052
rect 34609 5049 34621 5052
rect 34655 5049 34667 5083
rect 34609 5043 34667 5049
rect 25455 4984 26188 5012
rect 26789 5015 26847 5021
rect 25455 4981 25467 4984
rect 25409 4975 25467 4981
rect 26789 4981 26801 5015
rect 26835 5012 26847 5015
rect 27617 5015 27675 5021
rect 27617 5012 27629 5015
rect 26835 4984 27629 5012
rect 26835 4981 26847 4984
rect 26789 4975 26847 4981
rect 27617 4981 27629 4984
rect 27663 5012 27675 5015
rect 28534 5012 28540 5024
rect 27663 4984 28540 5012
rect 27663 4981 27675 4984
rect 27617 4975 27675 4981
rect 28534 4972 28540 4984
rect 28592 4972 28598 5024
rect 30466 4972 30472 5024
rect 30524 5012 30530 5024
rect 30561 5015 30619 5021
rect 30561 5012 30573 5015
rect 30524 4984 30573 5012
rect 30524 4972 30530 4984
rect 30561 4981 30573 4984
rect 30607 4981 30619 5015
rect 33686 5012 33692 5024
rect 33647 4984 33692 5012
rect 30561 4975 30619 4981
rect 33686 4972 33692 4984
rect 33744 4972 33750 5024
rect 34054 4972 34060 5024
rect 34112 5012 34118 5024
rect 34333 5015 34391 5021
rect 34333 5012 34345 5015
rect 34112 4984 34345 5012
rect 34112 4972 34118 4984
rect 34333 4981 34345 4984
rect 34379 5012 34391 5015
rect 34974 5012 34980 5024
rect 34379 4984 34980 5012
rect 34379 4981 34391 4984
rect 34333 4975 34391 4981
rect 34974 4972 34980 4984
rect 35032 4972 35038 5024
rect 1104 4922 38824 4944
rect 1104 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 27648 4922
rect 27700 4870 27712 4922
rect 27764 4870 27776 4922
rect 27828 4870 27840 4922
rect 27892 4870 38824 4922
rect 1104 4848 38824 4870
rect 1670 4808 1676 4820
rect 1631 4780 1676 4808
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 2130 4808 2136 4820
rect 2091 4780 2136 4808
rect 2130 4768 2136 4780
rect 2188 4768 2194 4820
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3878 4808 3884 4820
rect 2832 4780 3884 4808
rect 2832 4768 2838 4780
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 5718 4768 5724 4820
rect 5776 4808 5782 4820
rect 5997 4811 6055 4817
rect 5997 4808 6009 4811
rect 5776 4780 6009 4808
rect 5776 4768 5782 4780
rect 5997 4777 6009 4780
rect 6043 4777 6055 4811
rect 5997 4771 6055 4777
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 7745 4811 7803 4817
rect 7745 4808 7757 4811
rect 7248 4780 7757 4808
rect 7248 4768 7254 4780
rect 7745 4777 7757 4780
rect 7791 4808 7803 4811
rect 8202 4808 8208 4820
rect 7791 4780 8208 4808
rect 7791 4777 7803 4780
rect 7745 4771 7803 4777
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 10226 4768 10232 4820
rect 10284 4808 10290 4820
rect 10870 4808 10876 4820
rect 10284 4780 10876 4808
rect 10284 4768 10290 4780
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 11054 4768 11060 4820
rect 11112 4808 11118 4820
rect 11241 4811 11299 4817
rect 11241 4808 11253 4811
rect 11112 4780 11253 4808
rect 11112 4768 11118 4780
rect 11241 4777 11253 4780
rect 11287 4777 11299 4811
rect 11241 4771 11299 4777
rect 11977 4811 12035 4817
rect 11977 4777 11989 4811
rect 12023 4808 12035 4811
rect 12342 4808 12348 4820
rect 12023 4780 12348 4808
rect 12023 4777 12035 4780
rect 11977 4771 12035 4777
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 15749 4811 15807 4817
rect 15749 4777 15761 4811
rect 15795 4808 15807 4811
rect 16114 4808 16120 4820
rect 15795 4780 16120 4808
rect 15795 4777 15807 4780
rect 15749 4771 15807 4777
rect 16114 4768 16120 4780
rect 16172 4768 16178 4820
rect 16390 4808 16396 4820
rect 16351 4780 16396 4808
rect 16390 4768 16396 4780
rect 16448 4768 16454 4820
rect 17773 4811 17831 4817
rect 17773 4777 17785 4811
rect 17819 4808 17831 4811
rect 17862 4808 17868 4820
rect 17819 4780 17868 4808
rect 17819 4777 17831 4780
rect 17773 4771 17831 4777
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 18141 4811 18199 4817
rect 18141 4777 18153 4811
rect 18187 4808 18199 4811
rect 18598 4808 18604 4820
rect 18187 4780 18604 4808
rect 18187 4777 18199 4780
rect 18141 4771 18199 4777
rect 18598 4768 18604 4780
rect 18656 4768 18662 4820
rect 19797 4811 19855 4817
rect 19797 4777 19809 4811
rect 19843 4808 19855 4811
rect 20070 4808 20076 4820
rect 19843 4780 20076 4808
rect 19843 4777 19855 4780
rect 19797 4771 19855 4777
rect 20070 4768 20076 4780
rect 20128 4768 20134 4820
rect 20717 4811 20775 4817
rect 20717 4777 20729 4811
rect 20763 4808 20775 4811
rect 21818 4808 21824 4820
rect 20763 4780 21824 4808
rect 20763 4777 20775 4780
rect 20717 4771 20775 4777
rect 21818 4768 21824 4780
rect 21876 4768 21882 4820
rect 23198 4768 23204 4820
rect 23256 4808 23262 4820
rect 23753 4811 23811 4817
rect 23753 4808 23765 4811
rect 23256 4780 23765 4808
rect 23256 4768 23262 4780
rect 23753 4777 23765 4780
rect 23799 4777 23811 4811
rect 25685 4811 25743 4817
rect 25685 4808 25697 4811
rect 23753 4771 23811 4777
rect 25148 4780 25697 4808
rect 2869 4743 2927 4749
rect 2869 4709 2881 4743
rect 2915 4740 2927 4743
rect 2958 4740 2964 4752
rect 2915 4712 2964 4740
rect 2915 4709 2927 4712
rect 2869 4703 2927 4709
rect 2958 4700 2964 4712
rect 3016 4700 3022 4752
rect 7098 4700 7104 4752
rect 7156 4740 7162 4752
rect 7466 4740 7472 4752
rect 7156 4712 7472 4740
rect 7156 4700 7162 4712
rect 7466 4700 7472 4712
rect 7524 4740 7530 4752
rect 7561 4743 7619 4749
rect 7561 4740 7573 4743
rect 7524 4712 7573 4740
rect 7524 4700 7530 4712
rect 7561 4709 7573 4712
rect 7607 4709 7619 4743
rect 16132 4740 16160 4768
rect 18417 4743 18475 4749
rect 18417 4740 18429 4743
rect 16132 4712 18429 4740
rect 7561 4703 7619 4709
rect 18417 4709 18429 4712
rect 18463 4740 18475 4743
rect 18690 4740 18696 4752
rect 18463 4712 18696 4740
rect 18463 4709 18475 4712
rect 18417 4703 18475 4709
rect 18690 4700 18696 4712
rect 18748 4700 18754 4752
rect 21453 4743 21511 4749
rect 21453 4740 21465 4743
rect 20732 4712 21465 4740
rect 3418 4672 3424 4684
rect 3331 4644 3424 4672
rect 3418 4632 3424 4644
rect 3476 4672 3482 4684
rect 4332 4675 4390 4681
rect 4332 4672 4344 4675
rect 3476 4644 4344 4672
rect 3476 4632 3482 4644
rect 4332 4641 4344 4644
rect 4378 4672 4390 4675
rect 4706 4672 4712 4684
rect 4378 4644 4712 4672
rect 4378 4641 4390 4644
rect 4332 4635 4390 4641
rect 4706 4632 4712 4644
rect 4764 4632 4770 4684
rect 12345 4675 12403 4681
rect 12345 4641 12357 4675
rect 12391 4672 12403 4675
rect 12526 4672 12532 4684
rect 12391 4644 12532 4672
rect 12391 4641 12403 4644
rect 12345 4635 12403 4641
rect 12526 4632 12532 4644
rect 12584 4632 12590 4684
rect 15194 4632 15200 4684
rect 15252 4672 15258 4684
rect 15838 4672 15844 4684
rect 15252 4644 15844 4672
rect 15252 4632 15258 4644
rect 15838 4632 15844 4644
rect 15896 4672 15902 4684
rect 16485 4675 16543 4681
rect 16485 4672 16497 4675
rect 15896 4644 16497 4672
rect 15896 4632 15902 4644
rect 16485 4641 16497 4644
rect 16531 4641 16543 4675
rect 16485 4635 16543 4641
rect 2866 4604 2872 4616
rect 2827 4576 2872 4604
rect 2866 4564 2872 4576
rect 2924 4564 2930 4616
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4604 3019 4607
rect 3007 4576 3464 4604
rect 3007 4573 3019 4576
rect 2961 4567 3019 4573
rect 2406 4536 2412 4548
rect 2367 4508 2412 4536
rect 2406 4496 2412 4508
rect 2464 4496 2470 4548
rect 2130 4428 2136 4480
rect 2188 4468 2194 4480
rect 2976 4468 3004 4567
rect 3050 4468 3056 4480
rect 2188 4440 3056 4468
rect 2188 4428 2194 4440
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 3436 4468 3464 4576
rect 3878 4564 3884 4616
rect 3936 4604 3942 4616
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 3936 4576 4077 4604
rect 3936 4564 3942 4576
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4604 7895 4607
rect 7926 4604 7932 4616
rect 7883 4576 7932 4604
rect 7883 4573 7895 4576
rect 7837 4567 7895 4573
rect 7852 4536 7880 4567
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 10134 4604 10140 4616
rect 10095 4576 10140 4604
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 16390 4604 16396 4616
rect 16351 4576 16396 4604
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 19794 4604 19800 4616
rect 19755 4576 19800 4604
rect 19794 4564 19800 4576
rect 19852 4564 19858 4616
rect 19889 4607 19947 4613
rect 19889 4573 19901 4607
rect 19935 4604 19947 4607
rect 20254 4604 20260 4616
rect 19935 4576 20260 4604
rect 19935 4573 19947 4576
rect 19889 4567 19947 4573
rect 20254 4564 20260 4576
rect 20312 4564 20318 4616
rect 20732 4548 20760 4712
rect 21453 4709 21465 4712
rect 21499 4709 21511 4743
rect 21453 4703 21511 4709
rect 22922 4700 22928 4752
rect 22980 4740 22986 4752
rect 23569 4743 23627 4749
rect 23569 4740 23581 4743
rect 22980 4712 23581 4740
rect 22980 4700 22986 4712
rect 23569 4709 23581 4712
rect 23615 4740 23627 4743
rect 25148 4740 25176 4780
rect 25685 4777 25697 4780
rect 25731 4777 25743 4811
rect 25866 4808 25872 4820
rect 25827 4780 25872 4808
rect 25685 4771 25743 4777
rect 25866 4768 25872 4780
rect 25924 4768 25930 4820
rect 28626 4808 28632 4820
rect 28587 4780 28632 4808
rect 28626 4768 28632 4780
rect 28684 4768 28690 4820
rect 29641 4811 29699 4817
rect 29641 4777 29653 4811
rect 29687 4808 29699 4811
rect 29822 4808 29828 4820
rect 29687 4780 29828 4808
rect 29687 4777 29699 4780
rect 29641 4771 29699 4777
rect 29822 4768 29828 4780
rect 29880 4768 29886 4820
rect 30190 4768 30196 4820
rect 30248 4808 30254 4820
rect 30285 4811 30343 4817
rect 30285 4808 30297 4811
rect 30248 4780 30297 4808
rect 30248 4768 30254 4780
rect 30285 4777 30297 4780
rect 30331 4808 30343 4811
rect 30558 4808 30564 4820
rect 30331 4780 30564 4808
rect 30331 4777 30343 4780
rect 30285 4771 30343 4777
rect 30558 4768 30564 4780
rect 30616 4768 30622 4820
rect 30742 4808 30748 4820
rect 30703 4780 30748 4808
rect 30742 4768 30748 4780
rect 30800 4768 30806 4820
rect 32122 4768 32128 4820
rect 32180 4808 32186 4820
rect 32309 4811 32367 4817
rect 32309 4808 32321 4811
rect 32180 4780 32321 4808
rect 32180 4768 32186 4780
rect 32309 4777 32321 4780
rect 32355 4777 32367 4811
rect 32309 4771 32367 4777
rect 32769 4811 32827 4817
rect 32769 4777 32781 4811
rect 32815 4808 32827 4811
rect 33134 4808 33140 4820
rect 32815 4780 33140 4808
rect 32815 4777 32827 4780
rect 32769 4771 32827 4777
rect 25314 4740 25320 4752
rect 23615 4712 25176 4740
rect 25275 4712 25320 4740
rect 23615 4709 23627 4712
rect 23569 4703 23627 4709
rect 25314 4700 25320 4712
rect 25372 4700 25378 4752
rect 25409 4743 25467 4749
rect 25409 4709 25421 4743
rect 25455 4740 25467 4743
rect 25774 4740 25780 4752
rect 25455 4712 25780 4740
rect 25455 4709 25467 4712
rect 25409 4703 25467 4709
rect 21174 4632 21180 4684
rect 21232 4672 21238 4684
rect 21269 4675 21327 4681
rect 21269 4672 21281 4675
rect 21232 4644 21281 4672
rect 21232 4632 21238 4644
rect 21269 4641 21281 4644
rect 21315 4641 21327 4675
rect 23106 4672 23112 4684
rect 23019 4644 23112 4672
rect 21269 4635 21327 4641
rect 23106 4632 23112 4644
rect 23164 4672 23170 4684
rect 25130 4672 25136 4684
rect 23164 4644 23888 4672
rect 25091 4644 25136 4672
rect 23164 4632 23170 4644
rect 23860 4613 23888 4644
rect 25130 4632 25136 4644
rect 25188 4632 25194 4684
rect 21545 4607 21603 4613
rect 21545 4573 21557 4607
rect 21591 4604 21603 4607
rect 23845 4607 23903 4613
rect 21591 4576 21956 4604
rect 21591 4573 21603 4576
rect 21545 4567 21603 4573
rect 7024 4508 7880 4536
rect 5445 4471 5503 4477
rect 5445 4468 5457 4471
rect 3436 4440 5457 4468
rect 5445 4437 5457 4440
rect 5491 4437 5503 4471
rect 6638 4468 6644 4480
rect 6599 4440 6644 4468
rect 5445 4431 5503 4437
rect 6638 4428 6644 4440
rect 6696 4468 6702 4480
rect 7024 4477 7052 4508
rect 15746 4496 15752 4548
rect 15804 4536 15810 4548
rect 15933 4539 15991 4545
rect 15933 4536 15945 4539
rect 15804 4508 15945 4536
rect 15804 4496 15810 4508
rect 15933 4505 15945 4508
rect 15979 4505 15991 4539
rect 15933 4499 15991 4505
rect 19337 4539 19395 4545
rect 19337 4505 19349 4539
rect 19383 4536 19395 4539
rect 20714 4536 20720 4548
rect 19383 4508 20720 4536
rect 19383 4505 19395 4508
rect 19337 4499 19395 4505
rect 20714 4496 20720 4508
rect 20772 4496 20778 4548
rect 21928 4480 21956 4576
rect 23845 4573 23857 4607
rect 23891 4604 23903 4607
rect 25424 4604 25452 4703
rect 25774 4700 25780 4712
rect 25832 4700 25838 4752
rect 27522 4749 27528 4752
rect 26789 4743 26847 4749
rect 26789 4709 26801 4743
rect 26835 4740 26847 4743
rect 27516 4740 27528 4749
rect 26835 4712 27528 4740
rect 26835 4709 26847 4712
rect 26789 4703 26847 4709
rect 27516 4703 27528 4712
rect 27522 4700 27528 4703
rect 27580 4700 27586 4752
rect 30374 4700 30380 4752
rect 30432 4740 30438 4752
rect 30432 4712 30477 4740
rect 30432 4700 30438 4712
rect 25685 4675 25743 4681
rect 25685 4641 25697 4675
rect 25731 4672 25743 4675
rect 27065 4675 27123 4681
rect 27065 4672 27077 4675
rect 25731 4644 27077 4672
rect 25731 4641 25743 4644
rect 25685 4635 25743 4641
rect 27065 4641 27077 4644
rect 27111 4672 27123 4675
rect 27338 4672 27344 4684
rect 27111 4644 27344 4672
rect 27111 4641 27123 4644
rect 27065 4635 27123 4641
rect 27338 4632 27344 4644
rect 27396 4632 27402 4684
rect 33060 4672 33088 4780
rect 33134 4768 33140 4780
rect 33192 4768 33198 4820
rect 33410 4808 33416 4820
rect 33371 4780 33416 4808
rect 33410 4768 33416 4780
rect 33468 4768 33474 4820
rect 33226 4740 33232 4752
rect 33187 4712 33232 4740
rect 33226 4700 33232 4712
rect 33284 4700 33290 4752
rect 33505 4675 33563 4681
rect 33505 4672 33517 4675
rect 33060 4644 33517 4672
rect 33505 4641 33517 4644
rect 33551 4641 33563 4675
rect 33505 4635 33563 4641
rect 23891 4576 25452 4604
rect 23891 4573 23903 4576
rect 23845 4567 23903 4573
rect 26234 4564 26240 4616
rect 26292 4604 26298 4616
rect 26786 4604 26792 4616
rect 26292 4576 26792 4604
rect 26292 4564 26298 4576
rect 26786 4564 26792 4576
rect 26844 4604 26850 4616
rect 27249 4607 27307 4613
rect 27249 4604 27261 4607
rect 26844 4576 27261 4604
rect 26844 4564 26850 4576
rect 27249 4573 27261 4576
rect 27295 4573 27307 4607
rect 30282 4604 30288 4616
rect 30243 4576 30288 4604
rect 27249 4567 27307 4573
rect 30282 4564 30288 4576
rect 30340 4564 30346 4616
rect 23293 4539 23351 4545
rect 23293 4505 23305 4539
rect 23339 4536 23351 4539
rect 24118 4536 24124 4548
rect 23339 4508 24124 4536
rect 23339 4505 23351 4508
rect 23293 4499 23351 4505
rect 24118 4496 24124 4508
rect 24176 4536 24182 4548
rect 24581 4539 24639 4545
rect 24581 4536 24593 4539
rect 24176 4508 24593 4536
rect 24176 4496 24182 4508
rect 24581 4505 24593 4508
rect 24627 4505 24639 4539
rect 24581 4499 24639 4505
rect 29638 4496 29644 4548
rect 29696 4536 29702 4548
rect 29825 4539 29883 4545
rect 29825 4536 29837 4539
rect 29696 4508 29837 4536
rect 29696 4496 29702 4508
rect 29825 4505 29837 4508
rect 29871 4505 29883 4539
rect 32950 4536 32956 4548
rect 32911 4508 32956 4536
rect 29825 4499 29883 4505
rect 32950 4496 32956 4508
rect 33008 4496 33014 4548
rect 7009 4471 7067 4477
rect 7009 4468 7021 4471
rect 6696 4440 7021 4468
rect 6696 4428 6702 4440
rect 7009 4437 7021 4440
rect 7055 4437 7067 4471
rect 7282 4468 7288 4480
rect 7243 4440 7288 4468
rect 7009 4431 7067 4437
rect 7282 4428 7288 4440
rect 7340 4428 7346 4480
rect 8938 4468 8944 4480
rect 8899 4440 8944 4468
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 10502 4468 10508 4480
rect 10463 4440 10508 4468
rect 10502 4428 10508 4440
rect 10560 4428 10566 4480
rect 20254 4468 20260 4480
rect 20215 4440 20260 4468
rect 20254 4428 20260 4440
rect 20312 4428 20318 4480
rect 20806 4428 20812 4480
rect 20864 4468 20870 4480
rect 20993 4471 21051 4477
rect 20993 4468 21005 4471
rect 20864 4440 21005 4468
rect 20864 4428 20870 4440
rect 20993 4437 21005 4440
rect 21039 4437 21051 4471
rect 21910 4468 21916 4480
rect 21871 4440 21916 4468
rect 20993 4431 21051 4437
rect 21910 4428 21916 4440
rect 21968 4428 21974 4480
rect 24302 4468 24308 4480
rect 24263 4440 24308 4468
rect 24302 4428 24308 4440
rect 24360 4428 24366 4480
rect 24854 4468 24860 4480
rect 24815 4440 24860 4468
rect 24854 4428 24860 4440
rect 24912 4428 24918 4480
rect 29178 4468 29184 4480
rect 29139 4440 29184 4468
rect 29178 4428 29184 4440
rect 29236 4428 29242 4480
rect 31110 4468 31116 4480
rect 31071 4440 31116 4468
rect 31110 4428 31116 4440
rect 31168 4428 31174 4480
rect 1104 4378 38824 4400
rect 1104 4326 7648 4378
rect 7700 4326 7712 4378
rect 7764 4326 7776 4378
rect 7828 4326 7840 4378
rect 7892 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 34315 4378
rect 34367 4326 34379 4378
rect 34431 4326 34443 4378
rect 34495 4326 34507 4378
rect 34559 4326 38824 4378
rect 1104 4304 38824 4326
rect 2866 4224 2872 4276
rect 2924 4264 2930 4276
rect 3602 4264 3608 4276
rect 2924 4236 3608 4264
rect 2924 4224 2930 4236
rect 3602 4224 3608 4236
rect 3660 4264 3666 4276
rect 4065 4267 4123 4273
rect 4065 4264 4077 4267
rect 3660 4236 4077 4264
rect 3660 4224 3666 4236
rect 4065 4233 4077 4236
rect 4111 4233 4123 4267
rect 6638 4264 6644 4276
rect 6599 4236 6644 4264
rect 4065 4227 4123 4233
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 7190 4264 7196 4276
rect 7151 4236 7196 4264
rect 7190 4224 7196 4236
rect 7248 4224 7254 4276
rect 7377 4267 7435 4273
rect 7377 4233 7389 4267
rect 7423 4264 7435 4267
rect 7466 4264 7472 4276
rect 7423 4236 7472 4264
rect 7423 4233 7435 4236
rect 7377 4227 7435 4233
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 15838 4264 15844 4276
rect 15799 4236 15844 4264
rect 15838 4224 15844 4236
rect 15896 4224 15902 4276
rect 16298 4264 16304 4276
rect 16259 4236 16304 4264
rect 16298 4224 16304 4236
rect 16356 4224 16362 4276
rect 19705 4267 19763 4273
rect 19705 4233 19717 4267
rect 19751 4264 19763 4267
rect 20070 4264 20076 4276
rect 19751 4236 20076 4264
rect 19751 4233 19763 4236
rect 19705 4227 19763 4233
rect 20070 4224 20076 4236
rect 20128 4224 20134 4276
rect 21450 4224 21456 4276
rect 21508 4264 21514 4276
rect 23753 4267 23811 4273
rect 23753 4264 23765 4267
rect 21508 4236 23765 4264
rect 21508 4224 21514 4236
rect 23753 4233 23765 4236
rect 23799 4233 23811 4267
rect 23753 4227 23811 4233
rect 25593 4267 25651 4273
rect 25593 4233 25605 4267
rect 25639 4264 25651 4267
rect 25774 4264 25780 4276
rect 25639 4236 25780 4264
rect 25639 4233 25651 4236
rect 25593 4227 25651 4233
rect 25774 4224 25780 4236
rect 25832 4224 25838 4276
rect 26786 4264 26792 4276
rect 26747 4236 26792 4264
rect 26786 4224 26792 4236
rect 26844 4224 26850 4276
rect 27341 4267 27399 4273
rect 27341 4233 27353 4267
rect 27387 4264 27399 4267
rect 29178 4264 29184 4276
rect 27387 4236 29184 4264
rect 27387 4233 27399 4236
rect 27341 4227 27399 4233
rect 29178 4224 29184 4236
rect 29236 4224 29242 4276
rect 29914 4264 29920 4276
rect 29827 4236 29920 4264
rect 29914 4224 29920 4236
rect 29972 4264 29978 4276
rect 31110 4264 31116 4276
rect 29972 4236 31116 4264
rect 29972 4224 29978 4236
rect 31110 4224 31116 4236
rect 31168 4224 31174 4276
rect 33134 4224 33140 4276
rect 33192 4264 33198 4276
rect 33321 4267 33379 4273
rect 33321 4264 33333 4267
rect 33192 4236 33333 4264
rect 33192 4224 33198 4236
rect 33321 4233 33333 4236
rect 33367 4233 33379 4267
rect 33321 4227 33379 4233
rect 33410 4224 33416 4276
rect 33468 4264 33474 4276
rect 33597 4267 33655 4273
rect 33597 4264 33609 4267
rect 33468 4236 33609 4264
rect 33468 4224 33474 4236
rect 33597 4233 33609 4236
rect 33643 4233 33655 4267
rect 33597 4227 33655 4233
rect 2501 4199 2559 4205
rect 2501 4165 2513 4199
rect 2547 4165 2559 4199
rect 2501 4159 2559 4165
rect 8941 4199 8999 4205
rect 8941 4165 8953 4199
rect 8987 4165 8999 4199
rect 10502 4196 10508 4208
rect 8941 4159 8999 4165
rect 9600 4168 10508 4196
rect 2406 4088 2412 4140
rect 2464 4128 2470 4140
rect 2516 4128 2544 4159
rect 2866 4128 2872 4140
rect 2464 4100 2544 4128
rect 2827 4100 2872 4128
rect 2464 4088 2470 4100
rect 2866 4088 2872 4100
rect 2924 4088 2930 4140
rect 3050 4128 3056 4140
rect 3011 4100 3056 4128
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4128 3571 4131
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 3559 4100 4537 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 4525 4097 4537 4100
rect 4571 4128 4583 4131
rect 4614 4128 4620 4140
rect 4571 4100 4620 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 5994 4128 6000 4140
rect 5955 4100 6000 4128
rect 5994 4088 6000 4100
rect 6052 4088 6058 4140
rect 7929 4131 7987 4137
rect 7929 4097 7941 4131
rect 7975 4128 7987 4131
rect 8956 4128 8984 4159
rect 9600 4128 9628 4168
rect 10502 4156 10508 4168
rect 10560 4156 10566 4208
rect 19334 4156 19340 4208
rect 19392 4196 19398 4208
rect 19794 4196 19800 4208
rect 19392 4168 19800 4196
rect 19392 4156 19398 4168
rect 19794 4156 19800 4168
rect 19852 4156 19858 4208
rect 22830 4196 22836 4208
rect 22791 4168 22836 4196
rect 22830 4156 22836 4168
rect 22888 4156 22894 4208
rect 23198 4196 23204 4208
rect 23159 4168 23204 4196
rect 23198 4156 23204 4168
rect 23256 4156 23262 4208
rect 24857 4199 24915 4205
rect 24857 4165 24869 4199
rect 24903 4196 24915 4199
rect 25314 4196 25320 4208
rect 24903 4168 25320 4196
rect 24903 4165 24915 4168
rect 24857 4159 24915 4165
rect 25314 4156 25320 4168
rect 25372 4156 25378 4208
rect 26694 4156 26700 4208
rect 26752 4196 26758 4208
rect 26973 4199 27031 4205
rect 26973 4196 26985 4199
rect 26752 4168 26985 4196
rect 26752 4156 26758 4168
rect 26973 4165 26985 4168
rect 27019 4196 27031 4199
rect 27065 4199 27123 4205
rect 27065 4196 27077 4199
rect 27019 4168 27077 4196
rect 27019 4165 27031 4168
rect 26973 4159 27031 4165
rect 27065 4165 27077 4168
rect 27111 4165 27123 4199
rect 30466 4196 30472 4208
rect 27065 4159 27123 4165
rect 30392 4168 30472 4196
rect 16574 4128 16580 4140
rect 7975 4100 8892 4128
rect 8956 4100 9628 4128
rect 16535 4100 16580 4128
rect 7975 4097 7987 4100
rect 7929 4091 7987 4097
rect 1949 4063 2007 4069
rect 1949 4029 1961 4063
rect 1995 4060 2007 4063
rect 2774 4060 2780 4072
rect 1995 4032 2780 4060
rect 1995 4029 2007 4032
rect 1949 4023 2007 4029
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4060 5687 4063
rect 6086 4060 6092 4072
rect 5675 4032 6092 4060
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 7282 4020 7288 4072
rect 7340 4060 7346 4072
rect 7653 4063 7711 4069
rect 7653 4060 7665 4063
rect 7340 4032 7665 4060
rect 7340 4020 7346 4032
rect 7653 4029 7665 4032
rect 7699 4029 7711 4063
rect 8297 4063 8355 4069
rect 8297 4060 8309 4063
rect 7653 4023 7711 4029
rect 7852 4032 8309 4060
rect 2038 3952 2044 4004
rect 2096 3992 2102 4004
rect 2317 3995 2375 4001
rect 2317 3992 2329 3995
rect 2096 3964 2329 3992
rect 2096 3952 2102 3964
rect 2317 3961 2329 3964
rect 2363 3992 2375 3995
rect 2866 3992 2872 4004
rect 2363 3964 2872 3992
rect 2363 3961 2375 3964
rect 2317 3955 2375 3961
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 3786 3952 3792 4004
rect 3844 3992 3850 4004
rect 3881 3995 3939 4001
rect 3881 3992 3893 3995
rect 3844 3964 3893 3992
rect 3844 3952 3850 3964
rect 3881 3961 3893 3964
rect 3927 3992 3939 3995
rect 4522 3992 4528 4004
rect 3927 3964 4528 3992
rect 3927 3961 3939 3964
rect 3881 3955 3939 3961
rect 4522 3952 4528 3964
rect 4580 3952 4586 4004
rect 4617 3995 4675 4001
rect 4617 3961 4629 3995
rect 4663 3961 4675 3995
rect 4617 3955 4675 3961
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 2961 3927 3019 3933
rect 2961 3924 2973 3927
rect 2832 3896 2973 3924
rect 2832 3884 2838 3896
rect 2961 3893 2973 3896
rect 3007 3924 3019 3927
rect 3694 3924 3700 3936
rect 3007 3896 3700 3924
rect 3007 3893 3019 3896
rect 2961 3887 3019 3893
rect 3694 3884 3700 3896
rect 3752 3884 3758 3936
rect 4632 3924 4660 3955
rect 7374 3952 7380 4004
rect 7432 3992 7438 4004
rect 7852 4001 7880 4032
rect 8297 4029 8309 4032
rect 8343 4029 8355 4063
rect 8864 4060 8892 4100
rect 16574 4088 16580 4100
rect 16632 4088 16638 4140
rect 20073 4131 20131 4137
rect 20073 4097 20085 4131
rect 20119 4128 20131 4131
rect 20254 4128 20260 4140
rect 20119 4100 20260 4128
rect 20119 4097 20131 4100
rect 20073 4091 20131 4097
rect 20254 4088 20260 4100
rect 20312 4128 20318 4140
rect 25130 4128 25136 4140
rect 20312 4100 20944 4128
rect 25091 4100 25136 4128
rect 20312 4088 20318 4100
rect 9490 4060 9496 4072
rect 8864 4032 9496 4060
rect 8297 4023 8355 4029
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 20809 4063 20867 4069
rect 20809 4029 20821 4063
rect 20855 4029 20867 4063
rect 20916 4060 20944 4100
rect 25130 4088 25136 4100
rect 25188 4088 25194 4140
rect 26421 4131 26479 4137
rect 26421 4097 26433 4131
rect 26467 4128 26479 4131
rect 27522 4128 27528 4140
rect 26467 4100 27528 4128
rect 26467 4097 26479 4100
rect 26421 4091 26479 4097
rect 27522 4088 27528 4100
rect 27580 4128 27586 4140
rect 27893 4131 27951 4137
rect 27893 4128 27905 4131
rect 27580 4100 27905 4128
rect 27580 4088 27586 4100
rect 27893 4097 27905 4100
rect 27939 4097 27951 4131
rect 27893 4091 27951 4097
rect 29089 4131 29147 4137
rect 29089 4097 29101 4131
rect 29135 4128 29147 4131
rect 30392 4128 30420 4168
rect 30466 4156 30472 4168
rect 30524 4156 30530 4208
rect 33226 4196 33232 4208
rect 33060 4168 33232 4196
rect 29135 4100 30420 4128
rect 29135 4097 29147 4100
rect 29089 4091 29147 4097
rect 30558 4088 30564 4140
rect 30616 4128 30622 4140
rect 30837 4131 30895 4137
rect 30837 4128 30849 4131
rect 30616 4100 30849 4128
rect 30616 4088 30622 4100
rect 30837 4097 30849 4100
rect 30883 4097 30895 4131
rect 30837 4091 30895 4097
rect 32953 4131 33011 4137
rect 32953 4097 32965 4131
rect 32999 4128 33011 4131
rect 33060 4128 33088 4168
rect 33226 4156 33232 4168
rect 33284 4156 33290 4208
rect 32999 4100 33088 4128
rect 32999 4097 33011 4100
rect 32953 4091 33011 4097
rect 21082 4069 21088 4072
rect 21076 4060 21088 4069
rect 20916 4032 21088 4060
rect 20809 4023 20867 4029
rect 21076 4023 21088 4032
rect 7837 3995 7895 4001
rect 7837 3992 7849 3995
rect 7432 3964 7849 3992
rect 7432 3952 7438 3964
rect 7837 3961 7849 3964
rect 7883 3961 7895 3995
rect 9214 3992 9220 4004
rect 9127 3964 9220 3992
rect 7837 3955 7895 3961
rect 9214 3952 9220 3964
rect 9272 3952 9278 4004
rect 9398 3992 9404 4004
rect 9359 3964 9404 3992
rect 9398 3952 9404 3964
rect 9456 3952 9462 4004
rect 20717 3995 20775 4001
rect 20717 3961 20729 3995
rect 20763 3992 20775 3995
rect 20824 3992 20852 4023
rect 21082 4020 21088 4023
rect 21140 4020 21146 4072
rect 24026 4060 24032 4072
rect 23987 4032 24032 4060
rect 24026 4020 24032 4032
rect 24084 4020 24090 4072
rect 24854 4060 24860 4072
rect 24228 4032 24860 4060
rect 22002 3992 22008 4004
rect 20763 3964 22008 3992
rect 20763 3961 20775 3964
rect 20717 3955 20775 3961
rect 22002 3952 22008 3964
rect 22060 3952 22066 4004
rect 24228 4001 24256 4032
rect 24854 4020 24860 4032
rect 24912 4020 24918 4072
rect 30469 4063 30527 4069
rect 30469 4029 30481 4063
rect 30515 4060 30527 4063
rect 30742 4060 30748 4072
rect 30515 4032 30748 4060
rect 30515 4029 30527 4032
rect 30469 4023 30527 4029
rect 30742 4020 30748 4032
rect 30800 4020 30806 4072
rect 24213 3995 24271 4001
rect 24213 3961 24225 3995
rect 24259 3961 24271 3995
rect 24213 3955 24271 3961
rect 24302 3952 24308 4004
rect 24360 3992 24366 4004
rect 24360 3964 24405 3992
rect 24360 3952 24366 3964
rect 25038 3952 25044 4004
rect 25096 3992 25102 4004
rect 27338 3992 27344 4004
rect 25096 3964 27344 3992
rect 25096 3952 25102 3964
rect 27338 3952 27344 3964
rect 27396 3992 27402 4004
rect 27617 3995 27675 4001
rect 27617 3992 27629 3995
rect 27396 3964 27629 3992
rect 27396 3952 27402 3964
rect 27617 3961 27629 3964
rect 27663 3961 27675 3995
rect 30190 3992 30196 4004
rect 30151 3964 30196 3992
rect 27617 3955 27675 3961
rect 30190 3952 30196 3964
rect 30248 3952 30254 4004
rect 4706 3924 4712 3936
rect 4632 3896 4712 3924
rect 4706 3884 4712 3896
rect 4764 3924 4770 3936
rect 4985 3927 5043 3933
rect 4985 3924 4997 3927
rect 4764 3896 4997 3924
rect 4764 3884 4770 3896
rect 4985 3893 4997 3896
rect 5031 3893 5043 3927
rect 8662 3924 8668 3936
rect 8623 3896 8668 3924
rect 4985 3887 5043 3893
rect 8662 3884 8668 3896
rect 8720 3924 8726 3936
rect 9232 3924 9260 3952
rect 8720 3896 9260 3924
rect 8720 3884 8726 3896
rect 21910 3884 21916 3936
rect 21968 3924 21974 3936
rect 22189 3927 22247 3933
rect 22189 3924 22201 3927
rect 21968 3896 22201 3924
rect 21968 3884 21974 3896
rect 22189 3893 22201 3896
rect 22235 3893 22247 3927
rect 22189 3887 22247 3893
rect 26973 3927 27031 3933
rect 26973 3893 26985 3927
rect 27019 3924 27031 3927
rect 27801 3927 27859 3933
rect 27801 3924 27813 3927
rect 27019 3896 27813 3924
rect 27019 3893 27031 3896
rect 26973 3887 27031 3893
rect 27801 3893 27813 3896
rect 27847 3893 27859 3927
rect 29638 3924 29644 3936
rect 29599 3896 29644 3924
rect 27801 3887 27859 3893
rect 29638 3884 29644 3896
rect 29696 3924 29702 3936
rect 30377 3927 30435 3933
rect 30377 3924 30389 3927
rect 29696 3896 30389 3924
rect 29696 3884 29702 3896
rect 30377 3893 30389 3896
rect 30423 3924 30435 3927
rect 30558 3924 30564 3936
rect 30423 3896 30564 3924
rect 30423 3893 30435 3896
rect 30377 3887 30435 3893
rect 30558 3884 30564 3896
rect 30616 3884 30622 3936
rect 1104 3834 38824 3856
rect 1104 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 27648 3834
rect 27700 3782 27712 3834
rect 27764 3782 27776 3834
rect 27828 3782 27840 3834
rect 27892 3782 38824 3834
rect 1104 3760 38824 3782
rect 2498 3680 2504 3732
rect 2556 3720 2562 3732
rect 3050 3720 3056 3732
rect 2556 3692 3056 3720
rect 2556 3680 2562 3692
rect 3050 3680 3056 3692
rect 3108 3720 3114 3732
rect 3237 3723 3295 3729
rect 3237 3720 3249 3723
rect 3108 3692 3249 3720
rect 3108 3680 3114 3692
rect 3237 3689 3249 3692
rect 3283 3689 3295 3723
rect 3602 3720 3608 3732
rect 3563 3692 3608 3720
rect 3237 3683 3295 3689
rect 3602 3680 3608 3692
rect 3660 3680 3666 3732
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 7193 3723 7251 3729
rect 7193 3720 7205 3723
rect 7156 3692 7205 3720
rect 7156 3680 7162 3692
rect 7193 3689 7205 3692
rect 7239 3689 7251 3723
rect 7193 3683 7251 3689
rect 7282 3680 7288 3732
rect 7340 3720 7346 3732
rect 7929 3723 7987 3729
rect 7929 3720 7941 3723
rect 7340 3692 7941 3720
rect 7340 3680 7346 3692
rect 7929 3689 7941 3692
rect 7975 3689 7987 3723
rect 7929 3683 7987 3689
rect 9309 3723 9367 3729
rect 9309 3689 9321 3723
rect 9355 3720 9367 3723
rect 9398 3720 9404 3732
rect 9355 3692 9404 3720
rect 9355 3689 9367 3692
rect 9309 3683 9367 3689
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 20346 3720 20352 3732
rect 20307 3692 20352 3720
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 20714 3720 20720 3732
rect 20675 3692 20720 3720
rect 20714 3680 20720 3692
rect 20772 3680 20778 3732
rect 21082 3720 21088 3732
rect 21043 3692 21088 3720
rect 21082 3680 21088 3692
rect 21140 3680 21146 3732
rect 23753 3723 23811 3729
rect 23753 3689 23765 3723
rect 23799 3720 23811 3723
rect 24026 3720 24032 3732
rect 23799 3692 24032 3720
rect 23799 3689 23811 3692
rect 23753 3683 23811 3689
rect 24026 3680 24032 3692
rect 24084 3680 24090 3732
rect 24578 3680 24584 3732
rect 24636 3720 24642 3732
rect 24673 3723 24731 3729
rect 24673 3720 24685 3723
rect 24636 3692 24685 3720
rect 24636 3680 24642 3692
rect 24673 3689 24685 3692
rect 24719 3689 24731 3723
rect 24673 3683 24731 3689
rect 24854 3680 24860 3732
rect 24912 3720 24918 3732
rect 25133 3723 25191 3729
rect 25133 3720 25145 3723
rect 24912 3692 25145 3720
rect 24912 3680 24918 3692
rect 25133 3689 25145 3692
rect 25179 3689 25191 3723
rect 25133 3683 25191 3689
rect 27522 3680 27528 3732
rect 27580 3720 27586 3732
rect 27617 3723 27675 3729
rect 27617 3720 27629 3723
rect 27580 3692 27629 3720
rect 27580 3680 27586 3692
rect 27617 3689 27629 3692
rect 27663 3689 27675 3723
rect 27617 3683 27675 3689
rect 28994 3680 29000 3732
rect 29052 3720 29058 3732
rect 29825 3723 29883 3729
rect 29825 3720 29837 3723
rect 29052 3692 29837 3720
rect 29052 3680 29058 3692
rect 29825 3689 29837 3692
rect 29871 3720 29883 3723
rect 30190 3720 30196 3732
rect 29871 3692 30196 3720
rect 29871 3689 29883 3692
rect 29825 3683 29883 3689
rect 30190 3680 30196 3692
rect 30248 3680 30254 3732
rect 30374 3680 30380 3732
rect 30432 3720 30438 3732
rect 30561 3723 30619 3729
rect 30561 3720 30573 3723
rect 30432 3692 30573 3720
rect 30432 3680 30438 3692
rect 30561 3689 30573 3692
rect 30607 3689 30619 3723
rect 30561 3683 30619 3689
rect 1946 3612 1952 3664
rect 2004 3652 2010 3664
rect 2406 3652 2412 3664
rect 2004 3624 2412 3652
rect 2004 3612 2010 3624
rect 2406 3612 2412 3624
rect 2464 3612 2470 3664
rect 7653 3655 7711 3661
rect 7653 3621 7665 3655
rect 7699 3652 7711 3655
rect 8941 3655 8999 3661
rect 8941 3652 8953 3655
rect 7699 3624 8953 3652
rect 7699 3621 7711 3624
rect 7653 3615 7711 3621
rect 8941 3621 8953 3624
rect 8987 3652 8999 3655
rect 9490 3652 9496 3664
rect 8987 3624 9496 3652
rect 8987 3621 8999 3624
rect 8941 3615 8999 3621
rect 9490 3612 9496 3624
rect 9548 3612 9554 3664
rect 24762 3612 24768 3664
rect 24820 3652 24826 3664
rect 25774 3652 25780 3664
rect 24820 3624 25780 3652
rect 24820 3612 24826 3624
rect 25774 3612 25780 3624
rect 25832 3612 25838 3664
rect 30285 3655 30343 3661
rect 30285 3621 30297 3655
rect 30331 3652 30343 3655
rect 30742 3652 30748 3664
rect 30331 3624 30748 3652
rect 30331 3621 30343 3624
rect 30285 3615 30343 3621
rect 30742 3612 30748 3624
rect 30800 3612 30806 3664
rect 1765 3587 1823 3593
rect 1765 3553 1777 3587
rect 1811 3584 1823 3587
rect 2958 3584 2964 3596
rect 1811 3556 2964 3584
rect 1811 3553 1823 3556
rect 1765 3547 1823 3553
rect 2958 3544 2964 3556
rect 3016 3544 3022 3596
rect 21910 3593 21916 3596
rect 21545 3587 21603 3593
rect 21545 3553 21557 3587
rect 21591 3584 21603 3587
rect 21904 3584 21916 3593
rect 21591 3556 21916 3584
rect 21591 3553 21603 3556
rect 21545 3547 21603 3553
rect 21904 3547 21916 3556
rect 21910 3544 21916 3547
rect 21968 3544 21974 3596
rect 2314 3516 2320 3528
rect 2275 3488 2320 3516
rect 2314 3476 2320 3488
rect 2372 3476 2378 3528
rect 2406 3476 2412 3528
rect 2464 3516 2470 3528
rect 2501 3519 2559 3525
rect 2501 3516 2513 3519
rect 2464 3488 2513 3516
rect 2464 3476 2470 3488
rect 2501 3485 2513 3488
rect 2547 3485 2559 3519
rect 2501 3479 2559 3485
rect 21637 3519 21695 3525
rect 21637 3485 21649 3519
rect 21683 3485 21695 3519
rect 24670 3516 24676 3528
rect 24631 3488 24676 3516
rect 21637 3479 21695 3485
rect 1854 3408 1860 3460
rect 1912 3448 1918 3460
rect 1949 3451 2007 3457
rect 1949 3448 1961 3451
rect 1912 3420 1961 3448
rect 1912 3408 1918 3420
rect 1949 3417 1961 3420
rect 1995 3417 2007 3451
rect 1949 3411 2007 3417
rect 2866 3408 2872 3460
rect 2924 3448 2930 3460
rect 9582 3448 9588 3460
rect 2924 3420 9588 3448
rect 2924 3408 2930 3420
rect 9582 3408 9588 3420
rect 9640 3408 9646 3460
rect 21652 3392 21680 3479
rect 24670 3476 24676 3488
rect 24728 3476 24734 3528
rect 24210 3448 24216 3460
rect 24171 3420 24216 3448
rect 24210 3408 24216 3420
rect 24268 3408 24274 3460
rect 2961 3383 3019 3389
rect 2961 3349 2973 3383
rect 3007 3380 3019 3383
rect 3510 3380 3516 3392
rect 3007 3352 3516 3380
rect 3007 3349 3019 3352
rect 2961 3343 3019 3349
rect 3510 3340 3516 3352
rect 3568 3340 3574 3392
rect 3878 3340 3884 3392
rect 3936 3380 3942 3392
rect 4154 3380 4160 3392
rect 3936 3352 4160 3380
rect 3936 3340 3942 3352
rect 4154 3340 4160 3352
rect 4212 3380 4218 3392
rect 4249 3383 4307 3389
rect 4249 3380 4261 3383
rect 4212 3352 4261 3380
rect 4212 3340 4218 3352
rect 4249 3349 4261 3352
rect 4295 3349 4307 3383
rect 4706 3380 4712 3392
rect 4667 3352 4712 3380
rect 4249 3343 4307 3349
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 21634 3380 21640 3392
rect 21547 3352 21640 3380
rect 21634 3340 21640 3352
rect 21692 3380 21698 3392
rect 22002 3380 22008 3392
rect 21692 3352 22008 3380
rect 21692 3340 21698 3352
rect 22002 3340 22008 3352
rect 22060 3340 22066 3392
rect 23014 3380 23020 3392
rect 22975 3352 23020 3380
rect 23014 3340 23020 3352
rect 23072 3340 23078 3392
rect 27338 3380 27344 3392
rect 27299 3352 27344 3380
rect 27338 3340 27344 3352
rect 27396 3340 27402 3392
rect 1104 3290 38824 3312
rect 1104 3238 7648 3290
rect 7700 3238 7712 3290
rect 7764 3238 7776 3290
rect 7828 3238 7840 3290
rect 7892 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 34315 3290
rect 34367 3238 34379 3290
rect 34431 3238 34443 3290
rect 34495 3238 34507 3290
rect 34559 3238 38824 3290
rect 1104 3216 38824 3238
rect 2409 3179 2467 3185
rect 2409 3145 2421 3179
rect 2455 3176 2467 3179
rect 2498 3176 2504 3188
rect 2455 3148 2504 3176
rect 2455 3145 2467 3148
rect 2409 3139 2467 3145
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 2958 3176 2964 3188
rect 2919 3148 2964 3176
rect 2958 3136 2964 3148
rect 3016 3136 3022 3188
rect 6546 3176 6552 3188
rect 3436 3148 6552 3176
rect 1762 3000 1768 3052
rect 1820 3040 1826 3052
rect 1949 3043 2007 3049
rect 1949 3040 1961 3043
rect 1820 3012 1961 3040
rect 1820 3000 1826 3012
rect 1949 3009 1961 3012
rect 1995 3040 2007 3043
rect 2406 3040 2412 3052
rect 1995 3012 2412 3040
rect 1995 3009 2007 3012
rect 1949 3003 2007 3009
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 2958 3000 2964 3052
rect 3016 3040 3022 3052
rect 3436 3049 3464 3148
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 21634 3176 21640 3188
rect 21595 3148 21640 3176
rect 21634 3136 21640 3148
rect 21692 3136 21698 3188
rect 21910 3136 21916 3188
rect 21968 3176 21974 3188
rect 22005 3179 22063 3185
rect 22005 3176 22017 3179
rect 21968 3148 22017 3176
rect 21968 3136 21974 3148
rect 22005 3145 22017 3148
rect 22051 3145 22063 3179
rect 22005 3139 22063 3145
rect 24581 3179 24639 3185
rect 24581 3145 24593 3179
rect 24627 3176 24639 3179
rect 24670 3176 24676 3188
rect 24627 3148 24676 3176
rect 24627 3145 24639 3148
rect 24581 3139 24639 3145
rect 24670 3136 24676 3148
rect 24728 3136 24734 3188
rect 24762 3136 24768 3188
rect 24820 3176 24826 3188
rect 24857 3179 24915 3185
rect 24857 3176 24869 3179
rect 24820 3148 24869 3176
rect 24820 3136 24826 3148
rect 24857 3145 24869 3148
rect 24903 3145 24915 3179
rect 24857 3139 24915 3145
rect 20530 3108 20536 3120
rect 20491 3080 20536 3108
rect 20530 3068 20536 3080
rect 20588 3068 20594 3120
rect 3421 3043 3479 3049
rect 3421 3040 3433 3043
rect 3016 3012 3433 3040
rect 3016 3000 3022 3012
rect 3421 3009 3433 3012
rect 3467 3009 3479 3043
rect 5258 3040 5264 3052
rect 3421 3003 3479 3009
rect 4448 3012 5264 3040
rect 4448 2981 4476 3012
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 20349 3043 20407 3049
rect 20349 3009 20361 3043
rect 20395 3040 20407 3043
rect 21085 3043 21143 3049
rect 21085 3040 21097 3043
rect 20395 3012 21097 3040
rect 20395 3009 20407 3012
rect 20349 3003 20407 3009
rect 21085 3009 21097 3012
rect 21131 3040 21143 3043
rect 23014 3040 23020 3052
rect 21131 3012 23020 3040
rect 21131 3009 21143 3012
rect 21085 3003 21143 3009
rect 23014 3000 23020 3012
rect 23072 3000 23078 3052
rect 24213 3043 24271 3049
rect 24213 3009 24225 3043
rect 24259 3040 24271 3043
rect 24578 3040 24584 3052
rect 24259 3012 24584 3040
rect 24259 3009 24271 3012
rect 24213 3003 24271 3009
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 4433 2975 4491 2981
rect 4433 2941 4445 2975
rect 4479 2941 4491 2975
rect 4433 2935 4491 2941
rect 19981 2975 20039 2981
rect 19981 2941 19993 2975
rect 20027 2972 20039 2975
rect 20806 2972 20812 2984
rect 20027 2944 20812 2972
rect 20027 2941 20039 2944
rect 19981 2935 20039 2941
rect 20806 2932 20812 2944
rect 20864 2932 20870 2984
rect 3510 2864 3516 2916
rect 3568 2904 3574 2916
rect 4614 2904 4620 2916
rect 3568 2876 4620 2904
rect 3568 2864 3574 2876
rect 4614 2864 4620 2876
rect 4672 2864 4678 2916
rect 4709 2907 4767 2913
rect 4709 2873 4721 2907
rect 4755 2904 4767 2907
rect 4982 2904 4988 2916
rect 4755 2876 4988 2904
rect 4755 2873 4767 2876
rect 4709 2867 4767 2873
rect 4982 2864 4988 2876
rect 5040 2864 5046 2916
rect 20622 2864 20628 2916
rect 20680 2904 20686 2916
rect 20993 2907 21051 2913
rect 20993 2904 21005 2907
rect 20680 2876 21005 2904
rect 20680 2864 20686 2876
rect 20993 2873 21005 2876
rect 21039 2904 21051 2907
rect 21358 2904 21364 2916
rect 21039 2876 21364 2904
rect 21039 2873 21051 2876
rect 20993 2867 21051 2873
rect 21358 2864 21364 2876
rect 21416 2864 21422 2916
rect 2682 2836 2688 2848
rect 2643 2808 2688 2836
rect 2682 2796 2688 2808
rect 2740 2836 2746 2848
rect 3421 2839 3479 2845
rect 3421 2836 3433 2839
rect 2740 2808 3433 2836
rect 2740 2796 2746 2808
rect 3421 2805 3433 2808
rect 3467 2836 3479 2839
rect 6822 2836 6828 2848
rect 3467 2808 6828 2836
rect 3467 2805 3479 2808
rect 3421 2799 3479 2805
rect 6822 2796 6828 2808
rect 6880 2796 6886 2848
rect 1104 2746 38824 2768
rect 1104 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 27648 2746
rect 27700 2694 27712 2746
rect 27764 2694 27776 2746
rect 27828 2694 27840 2746
rect 27892 2694 38824 2746
rect 1104 2672 38824 2694
rect 1946 2632 1952 2644
rect 1907 2604 1952 2632
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 2314 2632 2320 2644
rect 2275 2604 2320 2632
rect 2314 2592 2320 2604
rect 2372 2592 2378 2644
rect 2958 2632 2964 2644
rect 2919 2604 2964 2632
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 5445 2635 5503 2641
rect 5445 2632 5457 2635
rect 4764 2604 5457 2632
rect 4764 2592 4770 2604
rect 5445 2601 5457 2604
rect 5491 2601 5503 2635
rect 5445 2595 5503 2601
rect 20533 2635 20591 2641
rect 20533 2601 20545 2635
rect 20579 2632 20591 2635
rect 20622 2632 20628 2644
rect 20579 2604 20628 2632
rect 20579 2601 20591 2604
rect 20533 2595 20591 2601
rect 20622 2592 20628 2604
rect 20680 2592 20686 2644
rect 4338 2505 4344 2508
rect 3881 2499 3939 2505
rect 3881 2465 3893 2499
rect 3927 2496 3939 2499
rect 4332 2496 4344 2505
rect 3927 2468 4344 2496
rect 3927 2465 3939 2468
rect 3881 2459 3939 2465
rect 4332 2459 4344 2468
rect 4338 2456 4344 2459
rect 4396 2456 4402 2508
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2428 3571 2431
rect 4062 2428 4068 2440
rect 3559 2400 4068 2428
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 4062 2388 4068 2400
rect 4120 2388 4126 2440
rect 1104 2202 38824 2224
rect 1104 2150 7648 2202
rect 7700 2150 7712 2202
rect 7764 2150 7776 2202
rect 7828 2150 7840 2202
rect 7892 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 34315 2202
rect 34367 2150 34379 2202
rect 34431 2150 34443 2202
rect 34495 2150 34507 2202
rect 34559 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 3424 14016 3476 14068
rect 7196 14016 7248 14068
rect 4068 13948 4120 14000
rect 6460 13948 6512 14000
rect 3332 13880 3384 13932
rect 7012 13880 7064 13932
rect 32864 13880 32916 13932
rect 34796 13880 34848 13932
rect 3056 13812 3108 13864
rect 7104 13812 7156 13864
rect 25412 13812 25464 13864
rect 31760 13812 31812 13864
rect 34612 13812 34664 13864
rect 35164 13744 35216 13796
rect 23572 13676 23624 13728
rect 30932 13676 30984 13728
rect 31208 13676 31260 13728
rect 31668 13676 31720 13728
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 27648 13574 27700 13626
rect 27712 13574 27764 13626
rect 27776 13574 27828 13626
rect 27840 13574 27892 13626
rect 2780 13472 2832 13524
rect 4344 13472 4396 13524
rect 2136 13404 2188 13456
rect 4620 13404 4672 13456
rect 24032 13472 24084 13524
rect 26148 13472 26200 13524
rect 25504 13404 25556 13456
rect 28540 13472 28592 13524
rect 31760 13472 31812 13524
rect 34520 13472 34572 13524
rect 36728 13515 36780 13524
rect 36728 13481 36737 13515
rect 36737 13481 36771 13515
rect 36771 13481 36780 13515
rect 36728 13472 36780 13481
rect 26608 13404 26660 13456
rect 28908 13404 28960 13456
rect 35072 13404 35124 13456
rect 5172 13379 5224 13388
rect 5172 13345 5181 13379
rect 5181 13345 5215 13379
rect 5215 13345 5224 13379
rect 5172 13336 5224 13345
rect 8024 13336 8076 13388
rect 17868 13336 17920 13388
rect 22468 13336 22520 13388
rect 22652 13379 22704 13388
rect 22652 13345 22661 13379
rect 22661 13345 22695 13379
rect 22695 13345 22704 13379
rect 22652 13336 22704 13345
rect 28724 13336 28776 13388
rect 30104 13379 30156 13388
rect 30104 13345 30113 13379
rect 30113 13345 30147 13379
rect 30147 13345 30156 13379
rect 30104 13336 30156 13345
rect 2044 13268 2096 13320
rect 2320 13268 2372 13320
rect 22836 13268 22888 13320
rect 25412 13268 25464 13320
rect 25688 13311 25740 13320
rect 25688 13277 25697 13311
rect 25697 13277 25731 13311
rect 25731 13277 25740 13311
rect 25688 13268 25740 13277
rect 7104 13243 7156 13252
rect 7104 13209 7113 13243
rect 7113 13209 7147 13243
rect 7147 13209 7156 13243
rect 7104 13200 7156 13209
rect 24584 13200 24636 13252
rect 27436 13268 27488 13320
rect 27988 13268 28040 13320
rect 30380 13311 30432 13320
rect 30380 13277 30389 13311
rect 30389 13277 30423 13311
rect 30423 13277 30432 13311
rect 30380 13268 30432 13277
rect 31208 13311 31260 13320
rect 31208 13277 31217 13311
rect 31217 13277 31251 13311
rect 31251 13277 31260 13311
rect 31208 13268 31260 13277
rect 25964 13200 26016 13252
rect 26056 13200 26108 13252
rect 32128 13336 32180 13388
rect 33416 13336 33468 13388
rect 34152 13336 34204 13388
rect 35532 13336 35584 13388
rect 36544 13379 36596 13388
rect 36544 13345 36553 13379
rect 36553 13345 36587 13379
rect 36587 13345 36596 13379
rect 36544 13336 36596 13345
rect 34704 13200 34756 13252
rect 1676 13132 1728 13184
rect 13728 13132 13780 13184
rect 16948 13132 17000 13184
rect 24308 13175 24360 13184
rect 24308 13141 24317 13175
rect 24317 13141 24351 13175
rect 24351 13141 24360 13175
rect 24308 13132 24360 13141
rect 24860 13132 24912 13184
rect 25044 13175 25096 13184
rect 25044 13141 25053 13175
rect 25053 13141 25087 13175
rect 25087 13141 25096 13175
rect 25044 13132 25096 13141
rect 25228 13175 25280 13184
rect 25228 13141 25237 13175
rect 25237 13141 25271 13175
rect 25271 13141 25280 13175
rect 25228 13132 25280 13141
rect 25596 13132 25648 13184
rect 26608 13175 26660 13184
rect 26608 13141 26617 13175
rect 26617 13141 26651 13175
rect 26651 13141 26660 13175
rect 26976 13175 27028 13184
rect 26608 13132 26660 13141
rect 26976 13141 26985 13175
rect 26985 13141 27019 13175
rect 27019 13141 27028 13175
rect 26976 13132 27028 13141
rect 27068 13132 27120 13184
rect 28908 13132 28960 13184
rect 29000 13132 29052 13184
rect 29828 13175 29880 13184
rect 29828 13141 29837 13175
rect 29837 13141 29871 13175
rect 29871 13141 29880 13175
rect 29828 13132 29880 13141
rect 35624 13175 35676 13184
rect 35624 13141 35633 13175
rect 35633 13141 35667 13175
rect 35667 13141 35676 13175
rect 35624 13132 35676 13141
rect 7648 13030 7700 13082
rect 7712 13030 7764 13082
rect 7776 13030 7828 13082
rect 7840 13030 7892 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 34315 13030 34367 13082
rect 34379 13030 34431 13082
rect 34443 13030 34495 13082
rect 34507 13030 34559 13082
rect 4620 12971 4672 12980
rect 4620 12937 4629 12971
rect 4629 12937 4663 12971
rect 4663 12937 4672 12971
rect 4620 12928 4672 12937
rect 5172 12971 5224 12980
rect 5172 12937 5181 12971
rect 5181 12937 5215 12971
rect 5215 12937 5224 12971
rect 5172 12928 5224 12937
rect 7012 12971 7064 12980
rect 7012 12937 7021 12971
rect 7021 12937 7055 12971
rect 7055 12937 7064 12971
rect 7012 12928 7064 12937
rect 2412 12860 2464 12912
rect 1216 12792 1268 12844
rect 4068 12792 4120 12844
rect 5632 12792 5684 12844
rect 6184 12792 6236 12844
rect 1492 12724 1544 12776
rect 5356 12724 5408 12776
rect 22836 12928 22888 12980
rect 25504 12971 25556 12980
rect 25504 12937 25513 12971
rect 25513 12937 25547 12971
rect 25547 12937 25556 12971
rect 25504 12928 25556 12937
rect 8024 12860 8076 12912
rect 14832 12903 14884 12912
rect 14832 12869 14841 12903
rect 14841 12869 14875 12903
rect 14875 12869 14884 12903
rect 14832 12860 14884 12869
rect 14924 12860 14976 12912
rect 17040 12860 17092 12912
rect 21548 12903 21600 12912
rect 21548 12869 21557 12903
rect 21557 12869 21591 12903
rect 21591 12869 21600 12903
rect 21548 12860 21600 12869
rect 24032 12903 24084 12912
rect 24032 12869 24041 12903
rect 24041 12869 24075 12903
rect 24075 12869 24084 12903
rect 24032 12860 24084 12869
rect 24584 12903 24636 12912
rect 24584 12869 24593 12903
rect 24593 12869 24627 12903
rect 24627 12869 24636 12903
rect 24584 12860 24636 12869
rect 26240 12860 26292 12912
rect 11152 12792 11204 12844
rect 16212 12792 16264 12844
rect 18420 12792 18472 12844
rect 23572 12792 23624 12844
rect 23664 12792 23716 12844
rect 24952 12792 25004 12844
rect 29368 12928 29420 12980
rect 29460 12928 29512 12980
rect 34612 12928 34664 12980
rect 35808 12928 35860 12980
rect 36544 12928 36596 12980
rect 27804 12860 27856 12912
rect 28448 12792 28500 12844
rect 28908 12860 28960 12912
rect 29736 12860 29788 12912
rect 31392 12860 31444 12912
rect 34796 12860 34848 12912
rect 30196 12835 30248 12844
rect 30196 12801 30205 12835
rect 30205 12801 30239 12835
rect 30239 12801 30248 12835
rect 30196 12792 30248 12801
rect 30380 12792 30432 12844
rect 30656 12835 30708 12844
rect 30656 12801 30665 12835
rect 30665 12801 30699 12835
rect 30699 12801 30708 12835
rect 30656 12792 30708 12801
rect 30932 12835 30984 12844
rect 30932 12801 30941 12835
rect 30941 12801 30975 12835
rect 30975 12801 30984 12835
rect 30932 12792 30984 12801
rect 31668 12792 31720 12844
rect 33600 12792 33652 12844
rect 35532 12792 35584 12844
rect 1400 12588 1452 12640
rect 2872 12699 2924 12708
rect 2872 12665 2881 12699
rect 2881 12665 2915 12699
rect 2915 12665 2924 12699
rect 2872 12656 2924 12665
rect 3516 12588 3568 12640
rect 10876 12631 10928 12640
rect 10876 12597 10885 12631
rect 10885 12597 10919 12631
rect 10919 12597 10928 12631
rect 10876 12588 10928 12597
rect 12532 12588 12584 12640
rect 13728 12724 13780 12776
rect 15016 12588 15068 12640
rect 15384 12699 15436 12708
rect 15384 12665 15393 12699
rect 15393 12665 15427 12699
rect 15427 12665 15436 12699
rect 16948 12724 17000 12776
rect 15384 12656 15436 12665
rect 20444 12656 20496 12708
rect 22376 12724 22428 12776
rect 22652 12724 22704 12776
rect 22192 12656 22244 12708
rect 15752 12588 15804 12640
rect 20536 12631 20588 12640
rect 20536 12597 20545 12631
rect 20545 12597 20579 12631
rect 20579 12597 20588 12631
rect 20536 12588 20588 12597
rect 20812 12588 20864 12640
rect 22468 12588 22520 12640
rect 23020 12588 23072 12640
rect 24308 12724 24360 12776
rect 26700 12724 26752 12776
rect 25044 12656 25096 12708
rect 25780 12588 25832 12640
rect 25872 12631 25924 12640
rect 25872 12597 25881 12631
rect 25881 12597 25915 12631
rect 25915 12597 25924 12631
rect 26424 12656 26476 12708
rect 28356 12656 28408 12708
rect 29092 12656 29144 12708
rect 29920 12699 29972 12708
rect 29920 12665 29929 12699
rect 29929 12665 29963 12699
rect 29963 12665 29972 12699
rect 29920 12656 29972 12665
rect 31208 12724 31260 12776
rect 32128 12767 32180 12776
rect 31760 12699 31812 12708
rect 31760 12665 31769 12699
rect 31769 12665 31803 12699
rect 31803 12665 31812 12699
rect 32128 12733 32137 12767
rect 32137 12733 32171 12767
rect 32171 12733 32180 12767
rect 32128 12724 32180 12733
rect 35440 12767 35492 12776
rect 35440 12733 35449 12767
rect 35449 12733 35483 12767
rect 35483 12733 35492 12767
rect 35440 12724 35492 12733
rect 31760 12656 31812 12665
rect 25872 12588 25924 12597
rect 26976 12588 27028 12640
rect 28264 12588 28316 12640
rect 29644 12588 29696 12640
rect 33416 12631 33468 12640
rect 33416 12597 33425 12631
rect 33425 12597 33459 12631
rect 33459 12597 33468 12631
rect 33416 12588 33468 12597
rect 34244 12631 34296 12640
rect 34244 12597 34253 12631
rect 34253 12597 34287 12631
rect 34287 12597 34296 12631
rect 34244 12588 34296 12597
rect 34796 12588 34848 12640
rect 35440 12588 35492 12640
rect 36728 12631 36780 12640
rect 36728 12597 36737 12631
rect 36737 12597 36771 12631
rect 36771 12597 36780 12631
rect 36728 12588 36780 12597
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 27648 12486 27700 12538
rect 27712 12486 27764 12538
rect 27776 12486 27828 12538
rect 27840 12486 27892 12538
rect 4160 12384 4212 12436
rect 6460 12427 6512 12436
rect 6460 12393 6469 12427
rect 6469 12393 6503 12427
rect 6503 12393 6512 12427
rect 6460 12384 6512 12393
rect 7196 12384 7248 12436
rect 20536 12384 20588 12436
rect 22192 12384 22244 12436
rect 26332 12384 26384 12436
rect 27528 12384 27580 12436
rect 28264 12427 28316 12436
rect 28264 12393 28273 12427
rect 28273 12393 28307 12427
rect 28307 12393 28316 12427
rect 28264 12384 28316 12393
rect 29920 12384 29972 12436
rect 31392 12384 31444 12436
rect 31668 12384 31720 12436
rect 32864 12427 32916 12436
rect 32864 12393 32873 12427
rect 32873 12393 32907 12427
rect 32907 12393 32916 12427
rect 32864 12384 32916 12393
rect 2504 12316 2556 12368
rect 12072 12316 12124 12368
rect 13636 12316 13688 12368
rect 17040 12316 17092 12368
rect 18696 12316 18748 12368
rect 20628 12316 20680 12368
rect 21732 12359 21784 12368
rect 21732 12325 21741 12359
rect 21741 12325 21775 12359
rect 21775 12325 21784 12359
rect 21732 12316 21784 12325
rect 23296 12359 23348 12368
rect 23296 12325 23305 12359
rect 23305 12325 23339 12359
rect 23339 12325 23348 12359
rect 23296 12316 23348 12325
rect 24952 12316 25004 12368
rect 25780 12316 25832 12368
rect 26240 12316 26292 12368
rect 28356 12359 28408 12368
rect 28356 12325 28365 12359
rect 28365 12325 28399 12359
rect 28399 12325 28408 12359
rect 28356 12316 28408 12325
rect 29828 12359 29880 12368
rect 29828 12325 29837 12359
rect 29837 12325 29871 12359
rect 29871 12325 29880 12359
rect 29828 12316 29880 12325
rect 34060 12359 34112 12368
rect 34060 12325 34069 12359
rect 34069 12325 34103 12359
rect 34103 12325 34112 12359
rect 34060 12316 34112 12325
rect 3424 12248 3476 12300
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5172 12248 5224 12257
rect 6184 12248 6236 12300
rect 7380 12291 7432 12300
rect 7380 12257 7389 12291
rect 7389 12257 7423 12291
rect 7423 12257 7432 12291
rect 7380 12248 7432 12257
rect 12348 12291 12400 12300
rect 12348 12257 12357 12291
rect 12357 12257 12391 12291
rect 12391 12257 12400 12291
rect 12348 12248 12400 12257
rect 13912 12248 13964 12300
rect 14832 12248 14884 12300
rect 17960 12291 18012 12300
rect 17960 12257 17969 12291
rect 17969 12257 18003 12291
rect 18003 12257 18012 12291
rect 17960 12248 18012 12257
rect 19524 12291 19576 12300
rect 19524 12257 19533 12291
rect 19533 12257 19567 12291
rect 19567 12257 19576 12291
rect 19524 12248 19576 12257
rect 21548 12291 21600 12300
rect 21548 12257 21557 12291
rect 21557 12257 21591 12291
rect 21591 12257 21600 12291
rect 21548 12248 21600 12257
rect 22928 12248 22980 12300
rect 25504 12291 25556 12300
rect 2320 12112 2372 12164
rect 2872 12180 2924 12232
rect 3516 12180 3568 12232
rect 3884 12180 3936 12232
rect 12716 12180 12768 12232
rect 4252 12155 4304 12164
rect 4252 12121 4261 12155
rect 4261 12121 4295 12155
rect 4295 12121 4304 12155
rect 4252 12112 4304 12121
rect 16120 12112 16172 12164
rect 2228 12087 2280 12096
rect 2228 12053 2237 12087
rect 2237 12053 2271 12087
rect 2271 12053 2280 12087
rect 2228 12044 2280 12053
rect 3608 12087 3660 12096
rect 3608 12053 3617 12087
rect 3617 12053 3651 12087
rect 3651 12053 3660 12087
rect 3608 12044 3660 12053
rect 6828 12087 6880 12096
rect 6828 12053 6837 12087
rect 6837 12053 6871 12087
rect 6871 12053 6880 12087
rect 6828 12044 6880 12053
rect 9496 12044 9548 12096
rect 12992 12087 13044 12096
rect 12992 12053 13001 12087
rect 13001 12053 13035 12087
rect 13035 12053 13044 12087
rect 12992 12044 13044 12053
rect 15108 12044 15160 12096
rect 16028 12044 16080 12096
rect 17132 12180 17184 12232
rect 21824 12223 21876 12232
rect 21824 12189 21833 12223
rect 21833 12189 21867 12223
rect 21867 12189 21876 12223
rect 21824 12180 21876 12189
rect 23848 12180 23900 12232
rect 24584 12112 24636 12164
rect 25504 12257 25513 12291
rect 25513 12257 25547 12291
rect 25547 12257 25556 12291
rect 25504 12248 25556 12257
rect 26976 12223 27028 12232
rect 26976 12189 26985 12223
rect 26985 12189 27019 12223
rect 27019 12189 27028 12223
rect 26976 12180 27028 12189
rect 27436 12180 27488 12232
rect 28816 12180 28868 12232
rect 29000 12180 29052 12232
rect 30196 12248 30248 12300
rect 30656 12291 30708 12300
rect 30656 12257 30665 12291
rect 30665 12257 30699 12291
rect 30699 12257 30708 12291
rect 30656 12248 30708 12257
rect 32680 12291 32732 12300
rect 29828 12223 29880 12232
rect 29828 12189 29837 12223
rect 29837 12189 29871 12223
rect 29871 12189 29880 12223
rect 29828 12180 29880 12189
rect 29920 12223 29972 12232
rect 29920 12189 29929 12223
rect 29929 12189 29963 12223
rect 29963 12189 29972 12223
rect 29920 12180 29972 12189
rect 30564 12180 30616 12232
rect 32680 12257 32689 12291
rect 32689 12257 32723 12291
rect 32723 12257 32732 12291
rect 32680 12248 32732 12257
rect 33784 12291 33836 12300
rect 33784 12257 33793 12291
rect 33793 12257 33827 12291
rect 33827 12257 33836 12291
rect 33784 12248 33836 12257
rect 34980 12248 35032 12300
rect 36452 12248 36504 12300
rect 25596 12112 25648 12164
rect 28448 12112 28500 12164
rect 28632 12112 28684 12164
rect 29368 12155 29420 12164
rect 29368 12121 29377 12155
rect 29377 12121 29411 12155
rect 29411 12121 29420 12155
rect 29368 12112 29420 12121
rect 21272 12087 21324 12096
rect 21272 12053 21281 12087
rect 21281 12053 21315 12087
rect 21315 12053 21324 12087
rect 21272 12044 21324 12053
rect 21732 12044 21784 12096
rect 24400 12087 24452 12096
rect 24400 12053 24409 12087
rect 24409 12053 24443 12087
rect 24443 12053 24452 12087
rect 24400 12044 24452 12053
rect 25688 12044 25740 12096
rect 26424 12044 26476 12096
rect 27804 12087 27856 12096
rect 27804 12053 27813 12087
rect 27813 12053 27847 12087
rect 27847 12053 27856 12087
rect 27804 12044 27856 12053
rect 33324 12087 33376 12096
rect 33324 12053 33333 12087
rect 33333 12053 33367 12087
rect 33367 12053 33376 12087
rect 33324 12044 33376 12053
rect 33692 12087 33744 12096
rect 33692 12053 33701 12087
rect 33701 12053 33735 12087
rect 33735 12053 33744 12087
rect 33692 12044 33744 12053
rect 35624 12087 35676 12096
rect 35624 12053 35633 12087
rect 35633 12053 35667 12087
rect 35667 12053 35676 12087
rect 35624 12044 35676 12053
rect 37188 12044 37240 12096
rect 7648 11942 7700 11994
rect 7712 11942 7764 11994
rect 7776 11942 7828 11994
rect 7840 11942 7892 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 34315 11942 34367 11994
rect 34379 11942 34431 11994
rect 34443 11942 34495 11994
rect 34507 11942 34559 11994
rect 5172 11840 5224 11892
rect 5632 11840 5684 11892
rect 12072 11883 12124 11892
rect 12072 11849 12081 11883
rect 12081 11849 12115 11883
rect 12115 11849 12124 11883
rect 12072 11840 12124 11849
rect 13912 11883 13964 11892
rect 13912 11849 13921 11883
rect 13921 11849 13955 11883
rect 13955 11849 13964 11883
rect 13912 11840 13964 11849
rect 1584 11815 1636 11824
rect 1584 11781 1593 11815
rect 1593 11781 1627 11815
rect 1627 11781 1636 11815
rect 1584 11772 1636 11781
rect 3792 11772 3844 11824
rect 4620 11772 4672 11824
rect 9220 11815 9272 11824
rect 9220 11781 9229 11815
rect 9229 11781 9263 11815
rect 9263 11781 9272 11815
rect 9220 11772 9272 11781
rect 12440 11772 12492 11824
rect 3516 11704 3568 11756
rect 4528 11747 4580 11756
rect 4528 11713 4537 11747
rect 4537 11713 4571 11747
rect 4571 11713 4580 11747
rect 4528 11704 4580 11713
rect 6276 11747 6328 11756
rect 1584 11636 1636 11688
rect 6276 11713 6285 11747
rect 6285 11713 6319 11747
rect 6319 11713 6328 11747
rect 6276 11704 6328 11713
rect 8668 11704 8720 11756
rect 9496 11704 9548 11756
rect 12900 11747 12952 11756
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 2596 11568 2648 11620
rect 3148 11611 3200 11620
rect 3148 11577 3157 11611
rect 3157 11577 3191 11611
rect 3191 11577 3200 11611
rect 3148 11568 3200 11577
rect 6828 11679 6880 11688
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 6828 11636 6880 11645
rect 9128 11636 9180 11688
rect 19524 11840 19576 11892
rect 21824 11883 21876 11892
rect 21824 11849 21833 11883
rect 21833 11849 21867 11883
rect 21867 11849 21876 11883
rect 21824 11840 21876 11849
rect 23296 11883 23348 11892
rect 23296 11849 23305 11883
rect 23305 11849 23339 11883
rect 23339 11849 23348 11883
rect 23296 11840 23348 11849
rect 16488 11815 16540 11824
rect 16488 11781 16497 11815
rect 16497 11781 16531 11815
rect 16531 11781 16540 11815
rect 16488 11772 16540 11781
rect 15384 11747 15436 11756
rect 15384 11713 15393 11747
rect 15393 11713 15427 11747
rect 15427 11713 15436 11747
rect 15384 11704 15436 11713
rect 15936 11704 15988 11756
rect 21732 11772 21784 11824
rect 26516 11840 26568 11892
rect 29460 11883 29512 11892
rect 29460 11849 29469 11883
rect 29469 11849 29503 11883
rect 29503 11849 29512 11883
rect 29460 11840 29512 11849
rect 31760 11883 31812 11892
rect 31760 11849 31769 11883
rect 31769 11849 31803 11883
rect 31803 11849 31812 11883
rect 31760 11840 31812 11849
rect 33784 11840 33836 11892
rect 28356 11772 28408 11824
rect 29920 11772 29972 11824
rect 21272 11747 21324 11756
rect 21272 11713 21281 11747
rect 21281 11713 21315 11747
rect 21315 11713 21324 11747
rect 21272 11704 21324 11713
rect 22376 11747 22428 11756
rect 22376 11713 22385 11747
rect 22385 11713 22419 11747
rect 22419 11713 22428 11747
rect 22376 11704 22428 11713
rect 24584 11747 24636 11756
rect 24584 11713 24593 11747
rect 24593 11713 24627 11747
rect 24627 11713 24636 11747
rect 24584 11704 24636 11713
rect 28908 11704 28960 11756
rect 33692 11747 33744 11756
rect 33692 11713 33701 11747
rect 33701 11713 33735 11747
rect 33735 11713 33744 11747
rect 33692 11704 33744 11713
rect 4712 11611 4764 11620
rect 4712 11577 4721 11611
rect 4721 11577 4755 11611
rect 4755 11577 4764 11611
rect 4712 11568 4764 11577
rect 3332 11500 3384 11552
rect 3424 11500 3476 11552
rect 6276 11500 6328 11552
rect 7380 11500 7432 11552
rect 8024 11500 8076 11552
rect 8944 11543 8996 11552
rect 8944 11509 8953 11543
rect 8953 11509 8987 11543
rect 8987 11509 8996 11543
rect 9588 11568 9640 11620
rect 16304 11636 16356 11688
rect 17868 11679 17920 11688
rect 9864 11568 9916 11620
rect 12716 11568 12768 11620
rect 12992 11611 13044 11620
rect 12992 11577 13001 11611
rect 13001 11577 13035 11611
rect 13035 11577 13044 11611
rect 12992 11568 13044 11577
rect 15108 11568 15160 11620
rect 17868 11645 17877 11679
rect 17877 11645 17911 11679
rect 17911 11645 17920 11679
rect 22928 11679 22980 11688
rect 17868 11636 17920 11645
rect 22928 11645 22937 11679
rect 22937 11645 22971 11679
rect 22971 11645 22980 11679
rect 22928 11636 22980 11645
rect 24032 11636 24084 11688
rect 13452 11543 13504 11552
rect 8944 11500 8996 11509
rect 13452 11509 13461 11543
rect 13461 11509 13495 11543
rect 13495 11509 13504 11543
rect 13452 11500 13504 11509
rect 15200 11500 15252 11552
rect 17132 11568 17184 11620
rect 17500 11611 17552 11620
rect 17500 11577 17509 11611
rect 17509 11577 17543 11611
rect 17543 11577 17552 11611
rect 17500 11568 17552 11577
rect 18604 11611 18656 11620
rect 18604 11577 18613 11611
rect 18613 11577 18647 11611
rect 18647 11577 18656 11611
rect 18604 11568 18656 11577
rect 18696 11611 18748 11620
rect 18696 11577 18705 11611
rect 18705 11577 18739 11611
rect 18739 11577 18748 11611
rect 18696 11568 18748 11577
rect 21456 11611 21508 11620
rect 21456 11577 21465 11611
rect 21465 11577 21499 11611
rect 21499 11577 21508 11611
rect 21456 11568 21508 11577
rect 21824 11568 21876 11620
rect 22376 11568 22428 11620
rect 24400 11568 24452 11620
rect 29184 11636 29236 11688
rect 30380 11679 30432 11688
rect 30380 11645 30389 11679
rect 30389 11645 30423 11679
rect 30423 11645 30432 11679
rect 30380 11636 30432 11645
rect 30656 11679 30708 11688
rect 30656 11645 30690 11679
rect 30690 11645 30708 11679
rect 30656 11636 30708 11645
rect 35256 11636 35308 11688
rect 36268 11636 36320 11688
rect 25780 11611 25832 11620
rect 25780 11577 25814 11611
rect 25814 11577 25832 11611
rect 25780 11568 25832 11577
rect 28264 11568 28316 11620
rect 28908 11568 28960 11620
rect 21732 11500 21784 11552
rect 22192 11543 22244 11552
rect 22192 11509 22201 11543
rect 22201 11509 22235 11543
rect 22235 11509 22244 11543
rect 22192 11500 22244 11509
rect 24952 11543 25004 11552
rect 24952 11509 24961 11543
rect 24961 11509 24995 11543
rect 24995 11509 25004 11543
rect 24952 11500 25004 11509
rect 25320 11543 25372 11552
rect 25320 11509 25329 11543
rect 25329 11509 25363 11543
rect 25363 11509 25372 11543
rect 25320 11500 25372 11509
rect 28816 11500 28868 11552
rect 30564 11500 30616 11552
rect 32404 11543 32456 11552
rect 32404 11509 32413 11543
rect 32413 11509 32447 11543
rect 32447 11509 32456 11543
rect 32404 11500 32456 11509
rect 32680 11543 32732 11552
rect 32680 11509 32689 11543
rect 32689 11509 32723 11543
rect 32723 11509 32732 11543
rect 32680 11500 32732 11509
rect 33324 11568 33376 11620
rect 33784 11611 33836 11620
rect 33784 11577 33793 11611
rect 33793 11577 33827 11611
rect 33827 11577 33836 11611
rect 33784 11568 33836 11577
rect 34704 11543 34756 11552
rect 34704 11509 34713 11543
rect 34713 11509 34747 11543
rect 34747 11509 34756 11543
rect 34704 11500 34756 11509
rect 34980 11500 35032 11552
rect 35808 11500 35860 11552
rect 36452 11543 36504 11552
rect 36452 11509 36461 11543
rect 36461 11509 36495 11543
rect 36495 11509 36504 11543
rect 36452 11500 36504 11509
rect 36728 11543 36780 11552
rect 36728 11509 36737 11543
rect 36737 11509 36771 11543
rect 36771 11509 36780 11543
rect 36728 11500 36780 11509
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 27648 11398 27700 11450
rect 27712 11398 27764 11450
rect 27776 11398 27828 11450
rect 27840 11398 27892 11450
rect 2228 11296 2280 11348
rect 3792 11339 3844 11348
rect 1584 11092 1636 11144
rect 2320 11092 2372 11144
rect 2136 11067 2188 11076
rect 2136 11033 2145 11067
rect 2145 11033 2179 11067
rect 2179 11033 2188 11067
rect 2136 11024 2188 11033
rect 2504 11160 2556 11212
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 9128 11339 9180 11348
rect 9128 11305 9137 11339
rect 9137 11305 9171 11339
rect 9171 11305 9180 11339
rect 9128 11296 9180 11305
rect 12348 11296 12400 11348
rect 15936 11339 15988 11348
rect 15936 11305 15945 11339
rect 15945 11305 15979 11339
rect 15979 11305 15988 11339
rect 15936 11296 15988 11305
rect 17040 11339 17092 11348
rect 17040 11305 17049 11339
rect 17049 11305 17083 11339
rect 17083 11305 17092 11339
rect 17040 11296 17092 11305
rect 21548 11296 21600 11348
rect 4344 11228 4396 11280
rect 4712 11271 4764 11280
rect 4712 11237 4721 11271
rect 4721 11237 4755 11271
rect 4755 11237 4764 11271
rect 4712 11228 4764 11237
rect 9220 11228 9272 11280
rect 16120 11228 16172 11280
rect 17132 11228 17184 11280
rect 17868 11271 17920 11280
rect 17868 11237 17880 11271
rect 17880 11237 17920 11271
rect 17868 11228 17920 11237
rect 22376 11228 22428 11280
rect 25136 11296 25188 11348
rect 25780 11339 25832 11348
rect 25780 11305 25789 11339
rect 25789 11305 25823 11339
rect 25823 11305 25832 11339
rect 25780 11296 25832 11305
rect 26332 11296 26384 11348
rect 28356 11296 28408 11348
rect 29092 11296 29144 11348
rect 29828 11296 29880 11348
rect 35900 11296 35952 11348
rect 6184 11160 6236 11212
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 12348 11160 12400 11212
rect 22192 11160 22244 11212
rect 22652 11160 22704 11212
rect 22928 11228 22980 11280
rect 25872 11228 25924 11280
rect 26976 11228 27028 11280
rect 28632 11228 28684 11280
rect 34428 11228 34480 11280
rect 35716 11228 35768 11280
rect 24124 11203 24176 11212
rect 24124 11169 24158 11203
rect 24158 11169 24176 11203
rect 24124 11160 24176 11169
rect 24676 11160 24728 11212
rect 27988 11160 28040 11212
rect 29184 11160 29236 11212
rect 30932 11203 30984 11212
rect 30932 11169 30941 11203
rect 30941 11169 30975 11203
rect 30975 11169 30984 11203
rect 30932 11160 30984 11169
rect 34704 11160 34756 11212
rect 36176 11203 36228 11212
rect 36176 11169 36185 11203
rect 36185 11169 36219 11203
rect 36219 11169 36228 11203
rect 36176 11160 36228 11169
rect 2688 11135 2740 11144
rect 2688 11101 2697 11135
rect 2697 11101 2731 11135
rect 2731 11101 2740 11135
rect 2688 11092 2740 11101
rect 3884 11092 3936 11144
rect 4344 11092 4396 11144
rect 4712 11092 4764 11144
rect 9588 11092 9640 11144
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 12164 11092 12216 11144
rect 16488 11135 16540 11144
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 16488 11092 16540 11101
rect 5816 11067 5868 11076
rect 5816 11033 5825 11067
rect 5825 11033 5859 11067
rect 5859 11033 5868 11067
rect 5816 11024 5868 11033
rect 9772 11067 9824 11076
rect 9772 11033 9781 11067
rect 9781 11033 9815 11067
rect 9815 11033 9824 11067
rect 9772 11024 9824 11033
rect 15200 11024 15252 11076
rect 16212 11024 16264 11076
rect 17316 11092 17368 11144
rect 21272 11092 21324 11144
rect 23756 11092 23808 11144
rect 25320 11092 25372 11144
rect 26516 11135 26568 11144
rect 26516 11101 26525 11135
rect 26525 11101 26559 11135
rect 26559 11101 26568 11135
rect 26516 11092 26568 11101
rect 27896 11067 27948 11076
rect 3148 10999 3200 11008
rect 3148 10965 3157 10999
rect 3157 10965 3191 10999
rect 3191 10965 3200 10999
rect 3148 10956 3200 10965
rect 7196 10956 7248 11008
rect 13636 10999 13688 11008
rect 13636 10965 13645 10999
rect 13645 10965 13679 10999
rect 13679 10965 13688 10999
rect 13636 10956 13688 10965
rect 16396 10956 16448 11008
rect 27896 11033 27905 11067
rect 27905 11033 27939 11067
rect 27939 11033 27948 11067
rect 27896 11024 27948 11033
rect 18696 10956 18748 11008
rect 20168 10956 20220 11008
rect 22468 10956 22520 11008
rect 23296 10999 23348 11008
rect 23296 10965 23305 10999
rect 23305 10965 23339 10999
rect 23339 10965 23348 10999
rect 23296 10956 23348 10965
rect 23848 10956 23900 11008
rect 28356 10956 28408 11008
rect 33048 11092 33100 11144
rect 33324 11135 33376 11144
rect 33324 11101 33333 11135
rect 33333 11101 33367 11135
rect 33367 11101 33376 11135
rect 33324 11092 33376 11101
rect 33508 11135 33560 11144
rect 33508 11101 33517 11135
rect 33517 11101 33551 11135
rect 33551 11101 33560 11135
rect 33508 11092 33560 11101
rect 35164 11135 35216 11144
rect 35164 11101 35173 11135
rect 35173 11101 35207 11135
rect 35207 11101 35216 11135
rect 35164 11092 35216 11101
rect 29000 11024 29052 11076
rect 30380 11067 30432 11076
rect 29368 10956 29420 11008
rect 30380 11033 30389 11067
rect 30389 11033 30423 11067
rect 30423 11033 30432 11067
rect 30380 11024 30432 11033
rect 32404 11024 32456 11076
rect 36360 11067 36412 11076
rect 36360 11033 36369 11067
rect 36369 11033 36403 11067
rect 36403 11033 36412 11067
rect 36360 11024 36412 11033
rect 33876 10999 33928 11008
rect 33876 10965 33885 10999
rect 33885 10965 33919 10999
rect 33919 10965 33928 10999
rect 33876 10956 33928 10965
rect 35900 10956 35952 11008
rect 36912 10956 36964 11008
rect 7648 10854 7700 10906
rect 7712 10854 7764 10906
rect 7776 10854 7828 10906
rect 7840 10854 7892 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 34315 10854 34367 10906
rect 34379 10854 34431 10906
rect 34443 10854 34495 10906
rect 34507 10854 34559 10906
rect 2504 10795 2556 10804
rect 2504 10761 2513 10795
rect 2513 10761 2547 10795
rect 2547 10761 2556 10795
rect 2504 10752 2556 10761
rect 3608 10752 3660 10804
rect 5724 10795 5776 10804
rect 5724 10761 5733 10795
rect 5733 10761 5767 10795
rect 5767 10761 5776 10795
rect 5724 10752 5776 10761
rect 9220 10752 9272 10804
rect 10324 10752 10376 10804
rect 12348 10752 12400 10804
rect 12532 10795 12584 10804
rect 12532 10761 12541 10795
rect 12541 10761 12575 10795
rect 12575 10761 12584 10795
rect 12532 10752 12584 10761
rect 16396 10752 16448 10804
rect 16488 10752 16540 10804
rect 17868 10752 17920 10804
rect 18696 10795 18748 10804
rect 18696 10761 18705 10795
rect 18705 10761 18739 10795
rect 18739 10761 18748 10795
rect 18696 10752 18748 10761
rect 21732 10752 21784 10804
rect 25964 10752 26016 10804
rect 26148 10752 26200 10804
rect 30656 10795 30708 10804
rect 30656 10761 30665 10795
rect 30665 10761 30699 10795
rect 30699 10761 30708 10795
rect 30656 10752 30708 10761
rect 33324 10795 33376 10804
rect 33324 10761 33333 10795
rect 33333 10761 33367 10795
rect 33367 10761 33376 10795
rect 33324 10752 33376 10761
rect 34796 10752 34848 10804
rect 36544 10795 36596 10804
rect 6920 10727 6972 10736
rect 6920 10693 6929 10727
rect 6929 10693 6963 10727
rect 6963 10693 6972 10727
rect 6920 10684 6972 10693
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 3792 10616 3844 10668
rect 4344 10616 4396 10668
rect 6184 10616 6236 10668
rect 12164 10616 12216 10668
rect 2964 10523 3016 10532
rect 2964 10489 2973 10523
rect 2973 10489 3007 10523
rect 3007 10489 3016 10523
rect 2964 10480 3016 10489
rect 3148 10480 3200 10532
rect 3240 10412 3292 10464
rect 3608 10412 3660 10464
rect 4712 10412 4764 10464
rect 5448 10455 5500 10464
rect 5448 10421 5457 10455
rect 5457 10421 5491 10455
rect 5491 10421 5500 10455
rect 5448 10412 5500 10421
rect 6184 10455 6236 10464
rect 6184 10421 6193 10455
rect 6193 10421 6227 10455
rect 6227 10421 6236 10455
rect 6184 10412 6236 10421
rect 6368 10412 6420 10464
rect 7196 10523 7248 10532
rect 7196 10489 7205 10523
rect 7205 10489 7239 10523
rect 7239 10489 7248 10523
rect 7196 10480 7248 10489
rect 10048 10548 10100 10600
rect 12808 10591 12860 10600
rect 12808 10557 12817 10591
rect 12817 10557 12851 10591
rect 12851 10557 12860 10591
rect 12808 10548 12860 10557
rect 16304 10616 16356 10668
rect 17500 10616 17552 10668
rect 14740 10548 14792 10600
rect 9496 10523 9548 10532
rect 9496 10489 9530 10523
rect 9530 10489 9548 10523
rect 13084 10523 13136 10532
rect 9496 10480 9548 10489
rect 13084 10489 13093 10523
rect 13093 10489 13127 10523
rect 13127 10489 13136 10523
rect 13084 10480 13136 10489
rect 13636 10480 13688 10532
rect 7012 10412 7064 10464
rect 8116 10412 8168 10464
rect 12164 10455 12216 10464
rect 12164 10421 12173 10455
rect 12173 10421 12207 10455
rect 12207 10421 12216 10455
rect 12164 10412 12216 10421
rect 12992 10455 13044 10464
rect 12992 10421 13001 10455
rect 13001 10421 13035 10455
rect 13035 10421 13044 10455
rect 12992 10412 13044 10421
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 17316 10412 17368 10464
rect 22100 10616 22152 10668
rect 26516 10684 26568 10736
rect 27160 10727 27212 10736
rect 27160 10693 27169 10727
rect 27169 10693 27203 10727
rect 27203 10693 27212 10727
rect 27160 10684 27212 10693
rect 32312 10727 32364 10736
rect 32312 10693 32321 10727
rect 32321 10693 32355 10727
rect 32355 10693 32364 10727
rect 32312 10684 32364 10693
rect 22376 10659 22428 10668
rect 22376 10625 22385 10659
rect 22385 10625 22419 10659
rect 22419 10625 22428 10659
rect 22376 10616 22428 10625
rect 22652 10616 22704 10668
rect 23848 10616 23900 10668
rect 33140 10616 33192 10668
rect 34704 10616 34756 10668
rect 23296 10548 23348 10600
rect 23664 10548 23716 10600
rect 23756 10548 23808 10600
rect 25136 10548 25188 10600
rect 25320 10548 25372 10600
rect 29368 10548 29420 10600
rect 32128 10591 32180 10600
rect 32128 10557 32137 10591
rect 32137 10557 32171 10591
rect 32171 10557 32180 10591
rect 32128 10548 32180 10557
rect 22284 10523 22336 10532
rect 22284 10489 22293 10523
rect 22293 10489 22327 10523
rect 22327 10489 22336 10523
rect 22284 10480 22336 10489
rect 25688 10480 25740 10532
rect 29092 10480 29144 10532
rect 31668 10480 31720 10532
rect 33600 10523 33652 10532
rect 33600 10489 33609 10523
rect 33609 10489 33643 10523
rect 33643 10489 33652 10523
rect 33600 10480 33652 10489
rect 36544 10761 36553 10795
rect 36553 10761 36587 10795
rect 36587 10761 36596 10795
rect 36544 10752 36596 10761
rect 35900 10616 35952 10668
rect 37096 10616 37148 10668
rect 35348 10480 35400 10532
rect 19524 10412 19576 10464
rect 21180 10412 21232 10464
rect 21272 10412 21324 10464
rect 23480 10412 23532 10464
rect 28356 10455 28408 10464
rect 28356 10421 28365 10455
rect 28365 10421 28399 10455
rect 28399 10421 28408 10455
rect 28356 10412 28408 10421
rect 28632 10455 28684 10464
rect 28632 10421 28641 10455
rect 28641 10421 28675 10455
rect 28675 10421 28684 10455
rect 28632 10412 28684 10421
rect 29184 10412 29236 10464
rect 30380 10412 30432 10464
rect 30932 10412 30984 10464
rect 32956 10412 33008 10464
rect 33324 10412 33376 10464
rect 33876 10412 33928 10464
rect 34336 10455 34388 10464
rect 34336 10421 34345 10455
rect 34345 10421 34379 10455
rect 34379 10421 34388 10455
rect 34336 10412 34388 10421
rect 35440 10455 35492 10464
rect 35440 10421 35449 10455
rect 35449 10421 35483 10455
rect 35483 10421 35492 10455
rect 35440 10412 35492 10421
rect 36176 10455 36228 10464
rect 36176 10421 36185 10455
rect 36185 10421 36219 10455
rect 36219 10421 36228 10455
rect 36176 10412 36228 10421
rect 36912 10412 36964 10464
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 27648 10310 27700 10362
rect 27712 10310 27764 10362
rect 27776 10310 27828 10362
rect 27840 10310 27892 10362
rect 2504 10251 2556 10260
rect 2504 10217 2513 10251
rect 2513 10217 2547 10251
rect 2547 10217 2556 10251
rect 2504 10208 2556 10217
rect 4344 10251 4396 10260
rect 4344 10217 4353 10251
rect 4353 10217 4387 10251
rect 4387 10217 4396 10251
rect 4344 10208 4396 10217
rect 5908 10251 5960 10260
rect 5908 10217 5917 10251
rect 5917 10217 5951 10251
rect 5951 10217 5960 10251
rect 5908 10208 5960 10217
rect 9680 10208 9732 10260
rect 10232 10251 10284 10260
rect 10232 10217 10241 10251
rect 10241 10217 10275 10251
rect 10275 10217 10284 10251
rect 10232 10208 10284 10217
rect 11336 10208 11388 10260
rect 12440 10208 12492 10260
rect 12992 10251 13044 10260
rect 12992 10217 13001 10251
rect 13001 10217 13035 10251
rect 13035 10217 13044 10251
rect 12992 10208 13044 10217
rect 16120 10251 16172 10260
rect 16120 10217 16129 10251
rect 16129 10217 16163 10251
rect 16163 10217 16172 10251
rect 16120 10208 16172 10217
rect 17868 10208 17920 10260
rect 22100 10208 22152 10260
rect 22652 10251 22704 10260
rect 22652 10217 22661 10251
rect 22661 10217 22695 10251
rect 22695 10217 22704 10251
rect 22652 10208 22704 10217
rect 24124 10251 24176 10260
rect 24124 10217 24133 10251
rect 24133 10217 24167 10251
rect 24167 10217 24176 10251
rect 24124 10208 24176 10217
rect 25228 10251 25280 10260
rect 25228 10217 25237 10251
rect 25237 10217 25271 10251
rect 25271 10217 25280 10251
rect 25228 10208 25280 10217
rect 26976 10251 27028 10260
rect 26976 10217 26985 10251
rect 26985 10217 27019 10251
rect 27019 10217 27028 10251
rect 26976 10208 27028 10217
rect 31760 10208 31812 10260
rect 36912 10208 36964 10260
rect 37096 10251 37148 10260
rect 37096 10217 37105 10251
rect 37105 10217 37139 10251
rect 37139 10217 37148 10251
rect 37096 10208 37148 10217
rect 2688 10140 2740 10192
rect 4528 10140 4580 10192
rect 7104 10072 7156 10124
rect 13084 10140 13136 10192
rect 13912 10140 13964 10192
rect 19340 10140 19392 10192
rect 21272 10140 21324 10192
rect 22008 10140 22060 10192
rect 22192 10140 22244 10192
rect 25688 10183 25740 10192
rect 25688 10149 25697 10183
rect 25697 10149 25731 10183
rect 25731 10149 25740 10183
rect 25688 10140 25740 10149
rect 27528 10140 27580 10192
rect 32956 10183 33008 10192
rect 32956 10149 32990 10183
rect 32990 10149 33008 10183
rect 32956 10140 33008 10149
rect 33048 10140 33100 10192
rect 35348 10140 35400 10192
rect 35532 10140 35584 10192
rect 9956 10072 10008 10124
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 2412 10004 2464 10013
rect 2044 9979 2096 9988
rect 2044 9945 2053 9979
rect 2053 9945 2087 9979
rect 2087 9945 2096 9979
rect 2044 9936 2096 9945
rect 3148 9868 3200 9920
rect 3884 9911 3936 9920
rect 3884 9877 3893 9911
rect 3893 9877 3927 9911
rect 3927 9877 3936 9911
rect 3884 9868 3936 9877
rect 9496 10004 9548 10056
rect 12072 10047 12124 10056
rect 10048 9936 10100 9988
rect 4712 9868 4764 9920
rect 6460 9911 6512 9920
rect 6460 9877 6469 9911
rect 6469 9877 6503 9911
rect 6503 9877 6512 9911
rect 6460 9868 6512 9877
rect 7012 9868 7064 9920
rect 8208 9868 8260 9920
rect 12072 10013 12081 10047
rect 12081 10013 12115 10047
rect 12115 10013 12124 10047
rect 12072 10004 12124 10013
rect 12808 10072 12860 10124
rect 14096 10072 14148 10124
rect 15108 10072 15160 10124
rect 16948 10072 17000 10124
rect 17592 10072 17644 10124
rect 21180 10115 21232 10124
rect 21180 10081 21189 10115
rect 21189 10081 21223 10115
rect 21223 10081 21232 10115
rect 21180 10072 21232 10081
rect 21824 10072 21876 10124
rect 21916 10072 21968 10124
rect 23756 10072 23808 10124
rect 24952 10072 25004 10124
rect 25320 10115 25372 10124
rect 12348 10004 12400 10056
rect 14188 10047 14240 10056
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 14188 10004 14240 10013
rect 15292 10004 15344 10056
rect 16396 10047 16448 10056
rect 16396 10013 16405 10047
rect 16405 10013 16439 10047
rect 16439 10013 16448 10047
rect 16396 10004 16448 10013
rect 19800 10047 19852 10056
rect 19800 10013 19809 10047
rect 19809 10013 19843 10047
rect 19843 10013 19852 10047
rect 19800 10004 19852 10013
rect 19892 10047 19944 10056
rect 19892 10013 19901 10047
rect 19901 10013 19935 10047
rect 19935 10013 19944 10047
rect 19892 10004 19944 10013
rect 12992 9936 13044 9988
rect 13544 9936 13596 9988
rect 20628 9936 20680 9988
rect 10968 9868 11020 9920
rect 19524 9868 19576 9920
rect 20444 9868 20496 9920
rect 21272 10047 21324 10056
rect 21272 10013 21281 10047
rect 21281 10013 21315 10047
rect 21315 10013 21324 10047
rect 23480 10047 23532 10056
rect 21272 10004 21324 10013
rect 23480 10013 23489 10047
rect 23489 10013 23523 10047
rect 23523 10013 23532 10047
rect 23480 10004 23532 10013
rect 25320 10081 25329 10115
rect 25329 10081 25363 10115
rect 25363 10081 25372 10115
rect 25320 10072 25372 10081
rect 26516 10047 26568 10056
rect 24216 9936 24268 9988
rect 26516 10013 26525 10047
rect 26525 10013 26559 10047
rect 26559 10013 26568 10047
rect 26516 10004 26568 10013
rect 28172 10047 28224 10056
rect 28172 10013 28181 10047
rect 28181 10013 28215 10047
rect 28215 10013 28224 10047
rect 28172 10004 28224 10013
rect 28356 10047 28408 10056
rect 28356 10013 28365 10047
rect 28365 10013 28399 10047
rect 28399 10013 28408 10047
rect 28356 10004 28408 10013
rect 28816 10004 28868 10056
rect 29736 10047 29788 10056
rect 29736 10013 29745 10047
rect 29745 10013 29779 10047
rect 29779 10013 29788 10047
rect 29736 10004 29788 10013
rect 35164 10047 35216 10056
rect 22652 9868 22704 9920
rect 24308 9868 24360 9920
rect 24768 9911 24820 9920
rect 24768 9877 24777 9911
rect 24777 9877 24811 9911
rect 24811 9877 24820 9911
rect 24768 9868 24820 9877
rect 27988 9868 28040 9920
rect 29184 9911 29236 9920
rect 29184 9877 29193 9911
rect 29193 9877 29227 9911
rect 29227 9877 29236 9911
rect 35164 10013 35173 10047
rect 35173 10013 35207 10047
rect 35207 10013 35216 10047
rect 35164 10004 35216 10013
rect 29184 9868 29236 9877
rect 30288 9868 30340 9920
rect 33784 9868 33836 9920
rect 35348 9868 35400 9920
rect 7648 9766 7700 9818
rect 7712 9766 7764 9818
rect 7776 9766 7828 9818
rect 7840 9766 7892 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 34315 9766 34367 9818
rect 34379 9766 34431 9818
rect 34443 9766 34495 9818
rect 34507 9766 34559 9818
rect 4528 9664 4580 9716
rect 5908 9664 5960 9716
rect 9956 9664 10008 9716
rect 14188 9664 14240 9716
rect 14740 9664 14792 9716
rect 15292 9664 15344 9716
rect 16396 9664 16448 9716
rect 17316 9664 17368 9716
rect 17592 9707 17644 9716
rect 17592 9673 17601 9707
rect 17601 9673 17635 9707
rect 17635 9673 17644 9707
rect 17592 9664 17644 9673
rect 19800 9664 19852 9716
rect 5540 9639 5592 9648
rect 5540 9605 5549 9639
rect 5549 9605 5583 9639
rect 5583 9605 5592 9639
rect 5540 9596 5592 9605
rect 10232 9596 10284 9648
rect 11980 9596 12032 9648
rect 13820 9639 13872 9648
rect 13820 9605 13829 9639
rect 13829 9605 13863 9639
rect 13863 9605 13872 9639
rect 13820 9596 13872 9605
rect 15016 9596 15068 9648
rect 18788 9639 18840 9648
rect 18788 9605 18797 9639
rect 18797 9605 18831 9639
rect 18831 9605 18840 9639
rect 18788 9596 18840 9605
rect 20352 9639 20404 9648
rect 20352 9605 20361 9639
rect 20361 9605 20395 9639
rect 20395 9605 20404 9639
rect 20352 9596 20404 9605
rect 21272 9664 21324 9716
rect 25136 9707 25188 9716
rect 23848 9639 23900 9648
rect 23848 9605 23857 9639
rect 23857 9605 23891 9639
rect 23891 9605 23900 9639
rect 23848 9596 23900 9605
rect 1860 9571 1912 9580
rect 1860 9537 1869 9571
rect 1869 9537 1903 9571
rect 1903 9537 1912 9571
rect 1860 9528 1912 9537
rect 2688 9528 2740 9580
rect 1584 9503 1636 9512
rect 1584 9469 1593 9503
rect 1593 9469 1627 9503
rect 1627 9469 1636 9503
rect 1584 9460 1636 9469
rect 2780 9460 2832 9512
rect 3884 9460 3936 9512
rect 4712 9460 4764 9512
rect 7104 9528 7156 9580
rect 11060 9528 11112 9580
rect 11428 9571 11480 9580
rect 11428 9537 11437 9571
rect 11437 9537 11471 9571
rect 11471 9537 11480 9571
rect 11428 9528 11480 9537
rect 8208 9460 8260 9512
rect 11244 9460 11296 9512
rect 12164 9503 12216 9512
rect 12164 9469 12173 9503
rect 12173 9469 12207 9503
rect 12207 9469 12216 9503
rect 12164 9460 12216 9469
rect 8116 9392 8168 9444
rect 11152 9435 11204 9444
rect 11152 9401 11161 9435
rect 11161 9401 11195 9435
rect 11195 9401 11204 9435
rect 11152 9392 11204 9401
rect 15108 9460 15160 9512
rect 15292 9503 15344 9512
rect 15292 9469 15301 9503
rect 15301 9469 15335 9503
rect 15335 9469 15344 9503
rect 15292 9460 15344 9469
rect 19524 9528 19576 9580
rect 19892 9528 19944 9580
rect 20076 9571 20128 9580
rect 20076 9537 20085 9571
rect 20085 9537 20119 9571
rect 20119 9537 20128 9571
rect 20076 9528 20128 9537
rect 22192 9528 22244 9580
rect 24676 9528 24728 9580
rect 25136 9673 25145 9707
rect 25145 9673 25179 9707
rect 25179 9673 25188 9707
rect 25136 9664 25188 9673
rect 25320 9664 25372 9716
rect 27160 9664 27212 9716
rect 27528 9596 27580 9648
rect 28540 9664 28592 9716
rect 29368 9596 29420 9648
rect 16764 9460 16816 9512
rect 20444 9460 20496 9512
rect 12716 9435 12768 9444
rect 12716 9401 12750 9435
rect 12750 9401 12768 9435
rect 12716 9392 12768 9401
rect 18880 9392 18932 9444
rect 20720 9392 20772 9444
rect 22008 9460 22060 9512
rect 25228 9460 25280 9512
rect 2688 9367 2740 9376
rect 2688 9333 2697 9367
rect 2697 9333 2731 9367
rect 2731 9333 2740 9367
rect 2688 9324 2740 9333
rect 6000 9367 6052 9376
rect 6000 9333 6009 9367
rect 6009 9333 6043 9367
rect 6043 9333 6052 9367
rect 6000 9324 6052 9333
rect 9036 9367 9088 9376
rect 9036 9333 9045 9367
rect 9045 9333 9079 9367
rect 9079 9333 9088 9367
rect 9036 9324 9088 9333
rect 10600 9367 10652 9376
rect 10600 9333 10609 9367
rect 10609 9333 10643 9367
rect 10643 9333 10652 9367
rect 10600 9324 10652 9333
rect 11428 9324 11480 9376
rect 16672 9367 16724 9376
rect 16672 9333 16681 9367
rect 16681 9333 16715 9367
rect 16715 9333 16724 9367
rect 16672 9324 16724 9333
rect 18328 9324 18380 9376
rect 19432 9324 19484 9376
rect 20076 9324 20128 9376
rect 23480 9392 23532 9444
rect 24308 9435 24360 9444
rect 24308 9401 24317 9435
rect 24317 9401 24351 9435
rect 24351 9401 24360 9435
rect 24308 9392 24360 9401
rect 25136 9392 25188 9444
rect 21272 9367 21324 9376
rect 21272 9333 21281 9367
rect 21281 9333 21315 9367
rect 21315 9333 21324 9367
rect 21272 9324 21324 9333
rect 21732 9367 21784 9376
rect 21732 9333 21741 9367
rect 21741 9333 21775 9367
rect 21775 9333 21784 9367
rect 22376 9367 22428 9376
rect 21732 9324 21784 9333
rect 22376 9333 22385 9367
rect 22385 9333 22419 9367
rect 22419 9333 22428 9367
rect 22376 9324 22428 9333
rect 24952 9324 25004 9376
rect 28908 9528 28960 9580
rect 29276 9528 29328 9580
rect 33048 9528 33100 9580
rect 25596 9503 25648 9512
rect 25596 9469 25630 9503
rect 25630 9469 25648 9503
rect 25596 9460 25648 9469
rect 26148 9460 26200 9512
rect 30288 9460 30340 9512
rect 32128 9503 32180 9512
rect 32128 9469 32137 9503
rect 32137 9469 32171 9503
rect 32171 9469 32180 9503
rect 32128 9460 32180 9469
rect 26608 9392 26660 9444
rect 28356 9392 28408 9444
rect 29092 9392 29144 9444
rect 28172 9324 28224 9376
rect 29184 9324 29236 9376
rect 32312 9367 32364 9376
rect 32312 9333 32321 9367
rect 32321 9333 32355 9367
rect 32355 9333 32364 9367
rect 32312 9324 32364 9333
rect 32772 9367 32824 9376
rect 32772 9333 32781 9367
rect 32781 9333 32815 9367
rect 32815 9333 32824 9367
rect 32772 9324 32824 9333
rect 33968 9596 34020 9648
rect 35164 9664 35216 9716
rect 34612 9596 34664 9648
rect 33784 9528 33836 9580
rect 37556 9571 37608 9580
rect 35532 9503 35584 9512
rect 35532 9469 35541 9503
rect 35541 9469 35575 9503
rect 35575 9469 35584 9503
rect 37556 9537 37565 9571
rect 37565 9537 37599 9571
rect 37599 9537 37608 9571
rect 37556 9528 37608 9537
rect 35532 9460 35584 9469
rect 33508 9392 33560 9444
rect 33876 9435 33928 9444
rect 33876 9401 33885 9435
rect 33885 9401 33919 9435
rect 33919 9401 33928 9435
rect 33876 9392 33928 9401
rect 35256 9435 35308 9444
rect 35256 9401 35265 9435
rect 35265 9401 35299 9435
rect 35299 9401 35308 9435
rect 35256 9392 35308 9401
rect 35440 9435 35492 9444
rect 35440 9401 35449 9435
rect 35449 9401 35483 9435
rect 35483 9401 35492 9435
rect 35440 9392 35492 9401
rect 33784 9367 33836 9376
rect 33784 9333 33793 9367
rect 33793 9333 33827 9367
rect 33827 9333 33836 9367
rect 33784 9324 33836 9333
rect 34428 9324 34480 9376
rect 34612 9367 34664 9376
rect 34612 9333 34621 9367
rect 34621 9333 34655 9367
rect 34655 9333 34664 9367
rect 34612 9324 34664 9333
rect 36912 9324 36964 9376
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 27648 9222 27700 9274
rect 27712 9222 27764 9274
rect 27776 9222 27828 9274
rect 27840 9222 27892 9274
rect 3976 9120 4028 9172
rect 4620 9163 4672 9172
rect 4620 9129 4629 9163
rect 4629 9129 4663 9163
rect 4663 9129 4672 9163
rect 4620 9120 4672 9129
rect 4988 9163 5040 9172
rect 4988 9129 4997 9163
rect 4997 9129 5031 9163
rect 5031 9129 5040 9163
rect 4988 9120 5040 9129
rect 8208 9163 8260 9172
rect 6092 9095 6144 9104
rect 6092 9061 6101 9095
rect 6101 9061 6135 9095
rect 6135 9061 6144 9095
rect 6092 9052 6144 9061
rect 7288 9052 7340 9104
rect 7472 9052 7524 9104
rect 8208 9129 8217 9163
rect 8217 9129 8251 9163
rect 8251 9129 8260 9163
rect 8208 9120 8260 9129
rect 9496 9163 9548 9172
rect 9496 9129 9505 9163
rect 9505 9129 9539 9163
rect 9539 9129 9548 9163
rect 9496 9120 9548 9129
rect 11336 9163 11388 9172
rect 11336 9129 11345 9163
rect 11345 9129 11379 9163
rect 11379 9129 11388 9163
rect 11336 9120 11388 9129
rect 14096 9163 14148 9172
rect 14096 9129 14105 9163
rect 14105 9129 14139 9163
rect 14139 9129 14148 9163
rect 14096 9120 14148 9129
rect 17592 9120 17644 9172
rect 19340 9120 19392 9172
rect 20352 9120 20404 9172
rect 10968 9052 11020 9104
rect 11428 9052 11480 9104
rect 11704 9095 11756 9104
rect 11704 9061 11727 9095
rect 11727 9061 11756 9095
rect 11704 9052 11756 9061
rect 19800 9095 19852 9104
rect 19800 9061 19809 9095
rect 19809 9061 19843 9095
rect 19843 9061 19852 9095
rect 19800 9052 19852 9061
rect 22192 9120 22244 9172
rect 25596 9163 25648 9172
rect 25596 9129 25605 9163
rect 25605 9129 25639 9163
rect 25639 9129 25648 9163
rect 25596 9120 25648 9129
rect 27160 9163 27212 9172
rect 27160 9129 27169 9163
rect 27169 9129 27203 9163
rect 27203 9129 27212 9163
rect 27160 9120 27212 9129
rect 27988 9120 28040 9172
rect 30932 9163 30984 9172
rect 30932 9129 30941 9163
rect 30941 9129 30975 9163
rect 30975 9129 30984 9163
rect 30932 9120 30984 9129
rect 35440 9120 35492 9172
rect 4620 8984 4672 9036
rect 6736 8984 6788 9036
rect 9036 8984 9088 9036
rect 10416 8984 10468 9036
rect 17132 8984 17184 9036
rect 19432 8984 19484 9036
rect 19984 8984 20036 9036
rect 21640 9052 21692 9104
rect 1952 8959 2004 8968
rect 1952 8925 1961 8959
rect 1961 8925 1995 8959
rect 1995 8925 2004 8959
rect 1952 8916 2004 8925
rect 2412 8959 2464 8968
rect 2412 8925 2421 8959
rect 2421 8925 2455 8959
rect 2455 8925 2464 8959
rect 2412 8916 2464 8925
rect 2688 8916 2740 8968
rect 4712 8916 4764 8968
rect 6092 8959 6144 8968
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 6552 8916 6604 8968
rect 7656 8959 7708 8968
rect 7656 8925 7665 8959
rect 7665 8925 7699 8959
rect 7699 8925 7708 8959
rect 7656 8916 7708 8925
rect 10508 8916 10560 8968
rect 11244 8916 11296 8968
rect 15108 8916 15160 8968
rect 20352 8916 20404 8968
rect 22192 8984 22244 9036
rect 24860 9052 24912 9104
rect 25228 9052 25280 9104
rect 26608 9052 26660 9104
rect 31852 9052 31904 9104
rect 26148 8984 26200 9036
rect 28724 8984 28776 9036
rect 29184 8984 29236 9036
rect 32956 9027 33008 9036
rect 32956 8993 32965 9027
rect 32965 8993 32999 9027
rect 32999 8993 33008 9027
rect 32956 8984 33008 8993
rect 33876 8984 33928 9036
rect 34428 9027 34480 9036
rect 34428 8993 34462 9027
rect 34462 8993 34480 9027
rect 34428 8984 34480 8993
rect 35900 8984 35952 9036
rect 23572 8959 23624 8968
rect 23572 8925 23581 8959
rect 23581 8925 23615 8959
rect 23615 8925 23624 8959
rect 23572 8916 23624 8925
rect 24308 8916 24360 8968
rect 25136 8959 25188 8968
rect 25136 8925 25145 8959
rect 25145 8925 25179 8959
rect 25179 8925 25188 8959
rect 25136 8916 25188 8925
rect 27252 8959 27304 8968
rect 27252 8925 27261 8959
rect 27261 8925 27295 8959
rect 27295 8925 27304 8959
rect 27252 8916 27304 8925
rect 29368 8916 29420 8968
rect 29552 8959 29604 8968
rect 29552 8925 29561 8959
rect 29561 8925 29595 8959
rect 29595 8925 29604 8959
rect 29552 8916 29604 8925
rect 33232 8959 33284 8968
rect 33232 8925 33241 8959
rect 33241 8925 33275 8959
rect 33275 8925 33284 8959
rect 33232 8916 33284 8925
rect 33968 8916 34020 8968
rect 36636 8959 36688 8968
rect 36636 8925 36645 8959
rect 36645 8925 36679 8959
rect 36679 8925 36688 8959
rect 36636 8916 36688 8925
rect 1492 8891 1544 8900
rect 1492 8857 1501 8891
rect 1501 8857 1535 8891
rect 1535 8857 1544 8891
rect 1492 8848 1544 8857
rect 3148 8848 3200 8900
rect 5724 8848 5776 8900
rect 6460 8848 6512 8900
rect 20812 8848 20864 8900
rect 23020 8891 23072 8900
rect 23020 8857 23029 8891
rect 23029 8857 23063 8891
rect 23063 8857 23072 8891
rect 23020 8848 23072 8857
rect 35532 8891 35584 8900
rect 35532 8857 35541 8891
rect 35541 8857 35575 8891
rect 35575 8857 35584 8891
rect 35532 8848 35584 8857
rect 1308 8780 1360 8832
rect 2964 8780 3016 8832
rect 4344 8780 4396 8832
rect 7472 8780 7524 8832
rect 9772 8823 9824 8832
rect 9772 8789 9781 8823
rect 9781 8789 9815 8823
rect 9815 8789 9824 8823
rect 9772 8780 9824 8789
rect 12164 8780 12216 8832
rect 13820 8780 13872 8832
rect 18880 8780 18932 8832
rect 20720 8780 20772 8832
rect 21640 8780 21692 8832
rect 21916 8823 21968 8832
rect 21916 8789 21925 8823
rect 21925 8789 21959 8823
rect 21959 8789 21968 8823
rect 21916 8780 21968 8789
rect 24216 8823 24268 8832
rect 24216 8789 24225 8823
rect 24225 8789 24259 8823
rect 24259 8789 24268 8823
rect 24216 8780 24268 8789
rect 26700 8823 26752 8832
rect 26700 8789 26709 8823
rect 26709 8789 26743 8823
rect 26743 8789 26752 8823
rect 26700 8780 26752 8789
rect 28908 8823 28960 8832
rect 28908 8789 28917 8823
rect 28917 8789 28951 8823
rect 28951 8789 28960 8823
rect 28908 8780 28960 8789
rect 29736 8780 29788 8832
rect 33140 8780 33192 8832
rect 33508 8780 33560 8832
rect 34060 8823 34112 8832
rect 34060 8789 34069 8823
rect 34069 8789 34103 8823
rect 34103 8789 34112 8823
rect 34060 8780 34112 8789
rect 7648 8678 7700 8730
rect 7712 8678 7764 8730
rect 7776 8678 7828 8730
rect 7840 8678 7892 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 34315 8678 34367 8730
rect 34379 8678 34431 8730
rect 34443 8678 34495 8730
rect 34507 8678 34559 8730
rect 1584 8551 1636 8560
rect 1584 8517 1593 8551
rect 1593 8517 1627 8551
rect 1627 8517 1636 8551
rect 1584 8508 1636 8517
rect 3884 8576 3936 8628
rect 4620 8619 4672 8628
rect 4620 8585 4629 8619
rect 4629 8585 4663 8619
rect 4663 8585 4672 8619
rect 4620 8576 4672 8585
rect 5080 8619 5132 8628
rect 5080 8585 5089 8619
rect 5089 8585 5123 8619
rect 5123 8585 5132 8619
rect 5080 8576 5132 8585
rect 6184 8576 6236 8628
rect 5264 8551 5316 8560
rect 5264 8517 5273 8551
rect 5273 8517 5307 8551
rect 5307 8517 5316 8551
rect 5264 8508 5316 8517
rect 6552 8576 6604 8628
rect 7012 8619 7064 8628
rect 7012 8585 7021 8619
rect 7021 8585 7055 8619
rect 7055 8585 7064 8619
rect 7012 8576 7064 8585
rect 8116 8576 8168 8628
rect 10968 8619 11020 8628
rect 7288 8508 7340 8560
rect 5724 8483 5776 8492
rect 5724 8449 5733 8483
rect 5733 8449 5767 8483
rect 5767 8449 5776 8483
rect 5724 8440 5776 8449
rect 8024 8440 8076 8492
rect 10968 8585 10977 8619
rect 10977 8585 11011 8619
rect 11011 8585 11020 8619
rect 10968 8576 11020 8585
rect 11244 8576 11296 8628
rect 11520 8576 11572 8628
rect 12072 8576 12124 8628
rect 14924 8576 14976 8628
rect 16764 8619 16816 8628
rect 16764 8585 16773 8619
rect 16773 8585 16807 8619
rect 16807 8585 16816 8619
rect 16764 8576 16816 8585
rect 18604 8576 18656 8628
rect 19064 8619 19116 8628
rect 19064 8585 19073 8619
rect 19073 8585 19107 8619
rect 19107 8585 19116 8619
rect 19064 8576 19116 8585
rect 19340 8619 19392 8628
rect 19340 8585 19349 8619
rect 19349 8585 19383 8619
rect 19383 8585 19392 8619
rect 19340 8576 19392 8585
rect 24308 8619 24360 8628
rect 24308 8585 24317 8619
rect 24317 8585 24351 8619
rect 24351 8585 24360 8619
rect 24308 8576 24360 8585
rect 24584 8576 24636 8628
rect 25136 8576 25188 8628
rect 26148 8619 26200 8628
rect 26148 8585 26157 8619
rect 26157 8585 26191 8619
rect 26191 8585 26200 8619
rect 26148 8576 26200 8585
rect 28908 8576 28960 8628
rect 29552 8576 29604 8628
rect 9956 8551 10008 8560
rect 9956 8517 9965 8551
rect 9965 8517 9999 8551
rect 9999 8517 10008 8551
rect 9956 8508 10008 8517
rect 11704 8508 11756 8560
rect 28724 8551 28776 8560
rect 28724 8517 28733 8551
rect 28733 8517 28767 8551
rect 28767 8517 28776 8551
rect 28724 8508 28776 8517
rect 29368 8551 29420 8560
rect 29368 8517 29377 8551
rect 29377 8517 29411 8551
rect 29411 8517 29420 8551
rect 29368 8508 29420 8517
rect 33876 8576 33928 8628
rect 35900 8619 35952 8628
rect 35900 8585 35909 8619
rect 35909 8585 35943 8619
rect 35943 8585 35952 8619
rect 35900 8576 35952 8585
rect 14464 8483 14516 8492
rect 1860 8236 1912 8288
rect 2688 8372 2740 8424
rect 6736 8372 6788 8424
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 14464 8449 14473 8483
rect 14473 8449 14507 8483
rect 14507 8449 14516 8483
rect 14464 8440 14516 8449
rect 15108 8440 15160 8492
rect 19524 8440 19576 8492
rect 19984 8440 20036 8492
rect 24216 8440 24268 8492
rect 26516 8483 26568 8492
rect 26516 8449 26525 8483
rect 26525 8449 26559 8483
rect 26559 8449 26568 8483
rect 26516 8440 26568 8449
rect 26608 8440 26660 8492
rect 28172 8483 28224 8492
rect 28172 8449 28181 8483
rect 28181 8449 28215 8483
rect 28215 8449 28224 8483
rect 28172 8440 28224 8449
rect 28816 8440 28868 8492
rect 29184 8440 29236 8492
rect 31300 8483 31352 8492
rect 31300 8449 31309 8483
rect 31309 8449 31343 8483
rect 31343 8449 31352 8483
rect 31300 8440 31352 8449
rect 11244 8372 11296 8424
rect 3148 8304 3200 8356
rect 5448 8304 5500 8356
rect 5724 8347 5776 8356
rect 5724 8313 5733 8347
rect 5733 8313 5767 8347
rect 5767 8313 5776 8347
rect 5724 8304 5776 8313
rect 5172 8236 5224 8288
rect 6368 8304 6420 8356
rect 9404 8304 9456 8356
rect 10508 8347 10560 8356
rect 10508 8313 10517 8347
rect 10517 8313 10551 8347
rect 10551 8313 10560 8347
rect 10508 8304 10560 8313
rect 14188 8347 14240 8356
rect 14188 8313 14197 8347
rect 14197 8313 14231 8347
rect 14231 8313 14240 8347
rect 14188 8304 14240 8313
rect 15200 8372 15252 8424
rect 19064 8372 19116 8424
rect 14648 8304 14700 8356
rect 15660 8347 15712 8356
rect 15660 8313 15694 8347
rect 15694 8313 15712 8347
rect 15660 8304 15712 8313
rect 18052 8347 18104 8356
rect 18052 8313 18061 8347
rect 18061 8313 18095 8347
rect 18095 8313 18104 8347
rect 18052 8304 18104 8313
rect 18604 8304 18656 8356
rect 20904 8372 20956 8424
rect 26148 8372 26200 8424
rect 27252 8372 27304 8424
rect 28908 8372 28960 8424
rect 34152 8508 34204 8560
rect 34060 8440 34112 8492
rect 35808 8440 35860 8492
rect 36820 8440 36872 8492
rect 20352 8347 20404 8356
rect 20352 8313 20361 8347
rect 20361 8313 20395 8347
rect 20395 8313 20404 8347
rect 20352 8304 20404 8313
rect 21456 8304 21508 8356
rect 23940 8304 23992 8356
rect 7472 8279 7524 8288
rect 7472 8245 7481 8279
rect 7481 8245 7515 8279
rect 7515 8245 7524 8279
rect 7472 8236 7524 8245
rect 12900 8236 12952 8288
rect 15108 8236 15160 8288
rect 17316 8279 17368 8288
rect 17316 8245 17325 8279
rect 17325 8245 17359 8279
rect 17359 8245 17368 8279
rect 17316 8236 17368 8245
rect 20904 8236 20956 8288
rect 22192 8279 22244 8288
rect 22192 8245 22201 8279
rect 22201 8245 22235 8279
rect 22235 8245 22244 8279
rect 22192 8236 22244 8245
rect 22928 8279 22980 8288
rect 22928 8245 22937 8279
rect 22937 8245 22971 8279
rect 22971 8245 22980 8279
rect 22928 8236 22980 8245
rect 23480 8236 23532 8288
rect 24308 8236 24360 8288
rect 26424 8304 26476 8356
rect 27068 8304 27120 8356
rect 28080 8304 28132 8356
rect 28264 8347 28316 8356
rect 28264 8313 28273 8347
rect 28273 8313 28307 8347
rect 28307 8313 28316 8347
rect 28264 8304 28316 8313
rect 29552 8304 29604 8356
rect 33048 8372 33100 8424
rect 33968 8372 34020 8424
rect 34428 8372 34480 8424
rect 36452 8415 36504 8424
rect 36452 8381 36461 8415
rect 36461 8381 36495 8415
rect 36495 8381 36504 8415
rect 36452 8372 36504 8381
rect 31852 8347 31904 8356
rect 31852 8313 31861 8347
rect 31861 8313 31895 8347
rect 31895 8313 31904 8347
rect 31852 8304 31904 8313
rect 32588 8347 32640 8356
rect 32588 8313 32622 8347
rect 32622 8313 32640 8347
rect 32588 8304 32640 8313
rect 33232 8304 33284 8356
rect 35440 8347 35492 8356
rect 26700 8236 26752 8288
rect 28356 8236 28408 8288
rect 30932 8279 30984 8288
rect 30932 8245 30941 8279
rect 30941 8245 30975 8279
rect 30975 8245 30984 8279
rect 30932 8236 30984 8245
rect 35440 8313 35449 8347
rect 35449 8313 35483 8347
rect 35483 8313 35492 8347
rect 35440 8304 35492 8313
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 27648 8134 27700 8186
rect 27712 8134 27764 8186
rect 27776 8134 27828 8186
rect 27840 8134 27892 8186
rect 2780 8032 2832 8084
rect 4252 8075 4304 8084
rect 4252 8041 4261 8075
rect 4261 8041 4295 8075
rect 4295 8041 4304 8075
rect 4252 8032 4304 8041
rect 5448 8032 5500 8084
rect 6092 8032 6144 8084
rect 2964 8007 3016 8016
rect 2964 7973 2973 8007
rect 2973 7973 3007 8007
rect 3007 7973 3016 8007
rect 2964 7964 3016 7973
rect 5172 8007 5224 8016
rect 5172 7973 5181 8007
rect 5181 7973 5215 8007
rect 5215 7973 5224 8007
rect 5172 7964 5224 7973
rect 6736 8007 6788 8016
rect 2412 7896 2464 7948
rect 4068 7939 4120 7948
rect 4068 7905 4077 7939
rect 4077 7905 4111 7939
rect 4111 7905 4120 7939
rect 4068 7896 4120 7905
rect 6736 7973 6745 8007
rect 6745 7973 6779 8007
rect 6779 7973 6788 8007
rect 6736 7964 6788 7973
rect 7012 7964 7064 8016
rect 7748 7964 7800 8016
rect 8208 8032 8260 8084
rect 9404 8075 9456 8084
rect 9404 8041 9413 8075
rect 9413 8041 9447 8075
rect 9447 8041 9456 8075
rect 9404 8032 9456 8041
rect 10232 8075 10284 8084
rect 10232 8041 10241 8075
rect 10241 8041 10275 8075
rect 10275 8041 10284 8075
rect 10232 8032 10284 8041
rect 15660 8032 15712 8084
rect 17132 8075 17184 8084
rect 17132 8041 17141 8075
rect 17141 8041 17175 8075
rect 17175 8041 17184 8075
rect 17132 8032 17184 8041
rect 18696 8075 18748 8084
rect 18696 8041 18705 8075
rect 18705 8041 18739 8075
rect 18739 8041 18748 8075
rect 18696 8032 18748 8041
rect 19984 8075 20036 8084
rect 19984 8041 19993 8075
rect 19993 8041 20027 8075
rect 20027 8041 20036 8075
rect 19984 8032 20036 8041
rect 20720 8032 20772 8084
rect 21456 8075 21508 8084
rect 21456 8041 21465 8075
rect 21465 8041 21499 8075
rect 21499 8041 21508 8075
rect 21456 8032 21508 8041
rect 21640 8032 21692 8084
rect 24768 8032 24820 8084
rect 26148 8075 26200 8084
rect 26148 8041 26157 8075
rect 26157 8041 26191 8075
rect 26191 8041 26200 8075
rect 26148 8032 26200 8041
rect 28172 8032 28224 8084
rect 30656 8075 30708 8084
rect 30656 8041 30665 8075
rect 30665 8041 30699 8075
rect 30699 8041 30708 8075
rect 30656 8032 30708 8041
rect 34888 8075 34940 8084
rect 34888 8041 34897 8075
rect 34897 8041 34931 8075
rect 34931 8041 34940 8075
rect 34888 8032 34940 8041
rect 35072 8032 35124 8084
rect 36452 8075 36504 8084
rect 36452 8041 36461 8075
rect 36461 8041 36495 8075
rect 36495 8041 36504 8075
rect 36452 8032 36504 8041
rect 36636 8032 36688 8084
rect 6920 7896 6972 7948
rect 3056 7871 3108 7880
rect 3056 7837 3065 7871
rect 3065 7837 3099 7871
rect 3099 7837 3108 7871
rect 3056 7828 3108 7837
rect 5264 7828 5316 7880
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 6184 7828 6236 7880
rect 7564 7871 7616 7880
rect 5356 7760 5408 7812
rect 7196 7760 7248 7812
rect 7564 7837 7573 7871
rect 7573 7837 7607 7871
rect 7607 7837 7616 7871
rect 7564 7828 7616 7837
rect 7472 7760 7524 7812
rect 7656 7760 7708 7812
rect 10784 7828 10836 7880
rect 12164 7964 12216 8016
rect 19800 7964 19852 8016
rect 25044 7964 25096 8016
rect 25320 8007 25372 8016
rect 25320 7973 25329 8007
rect 25329 7973 25363 8007
rect 25363 7973 25372 8007
rect 25320 7964 25372 7973
rect 11520 7939 11572 7948
rect 11520 7905 11529 7939
rect 11529 7905 11563 7939
rect 11563 7905 11572 7939
rect 11520 7896 11572 7905
rect 16764 7939 16816 7948
rect 16764 7905 16773 7939
rect 16773 7905 16807 7939
rect 16807 7905 16816 7939
rect 16764 7896 16816 7905
rect 17592 7939 17644 7948
rect 17592 7905 17626 7939
rect 17626 7905 17644 7939
rect 17592 7896 17644 7905
rect 20812 7896 20864 7948
rect 22192 7896 22244 7948
rect 23480 7896 23532 7948
rect 24952 7896 25004 7948
rect 16304 7871 16356 7880
rect 16304 7837 16313 7871
rect 16313 7837 16347 7871
rect 16347 7837 16356 7871
rect 16304 7828 16356 7837
rect 17316 7871 17368 7880
rect 17316 7837 17325 7871
rect 17325 7837 17359 7871
rect 17359 7837 17368 7871
rect 17316 7828 17368 7837
rect 21916 7828 21968 7880
rect 22100 7828 22152 7880
rect 25412 7871 25464 7880
rect 25412 7837 25421 7871
rect 25421 7837 25455 7871
rect 25455 7837 25464 7871
rect 25412 7828 25464 7837
rect 26976 7871 27028 7880
rect 26976 7837 26985 7871
rect 26985 7837 27019 7871
rect 27019 7837 27028 7871
rect 26976 7828 27028 7837
rect 11336 7803 11388 7812
rect 11336 7769 11345 7803
rect 11345 7769 11379 7803
rect 11379 7769 11388 7803
rect 11336 7760 11388 7769
rect 29092 7964 29144 8016
rect 33232 8007 33284 8016
rect 33232 7973 33266 8007
rect 33266 7973 33284 8007
rect 33232 7964 33284 7973
rect 35992 8007 36044 8016
rect 35992 7973 36001 8007
rect 36001 7973 36035 8007
rect 36035 7973 36044 8007
rect 35992 7964 36044 7973
rect 36084 7964 36136 8016
rect 28724 7939 28776 7948
rect 28724 7905 28733 7939
rect 28733 7905 28767 7939
rect 28767 7905 28776 7939
rect 28724 7896 28776 7905
rect 29460 7896 29512 7948
rect 33048 7896 33100 7948
rect 28080 7828 28132 7880
rect 32588 7760 32640 7812
rect 1860 7735 1912 7744
rect 1860 7701 1869 7735
rect 1869 7701 1903 7735
rect 1903 7701 1912 7735
rect 1860 7692 1912 7701
rect 2320 7692 2372 7744
rect 9772 7735 9824 7744
rect 9772 7701 9781 7735
rect 9781 7701 9815 7735
rect 9815 7701 9824 7735
rect 9772 7692 9824 7701
rect 10324 7692 10376 7744
rect 11152 7692 11204 7744
rect 12900 7735 12952 7744
rect 12900 7701 12909 7735
rect 12909 7701 12943 7735
rect 12943 7701 12952 7735
rect 12900 7692 12952 7701
rect 14188 7692 14240 7744
rect 14740 7692 14792 7744
rect 15844 7735 15896 7744
rect 15844 7701 15853 7735
rect 15853 7701 15887 7735
rect 15887 7701 15896 7735
rect 15844 7692 15896 7701
rect 19340 7735 19392 7744
rect 19340 7701 19349 7735
rect 19349 7701 19383 7735
rect 19383 7701 19392 7735
rect 19340 7692 19392 7701
rect 22928 7692 22980 7744
rect 23572 7692 23624 7744
rect 24308 7735 24360 7744
rect 24308 7701 24317 7735
rect 24317 7701 24351 7735
rect 24351 7701 24360 7735
rect 24308 7692 24360 7701
rect 26240 7692 26292 7744
rect 28264 7692 28316 7744
rect 30104 7735 30156 7744
rect 30104 7701 30113 7735
rect 30113 7701 30147 7735
rect 30147 7701 30156 7735
rect 30104 7692 30156 7701
rect 35440 7760 35492 7812
rect 33600 7692 33652 7744
rect 35256 7735 35308 7744
rect 35256 7701 35265 7735
rect 35265 7701 35299 7735
rect 35299 7701 35308 7735
rect 35256 7692 35308 7701
rect 36544 7692 36596 7744
rect 7648 7590 7700 7642
rect 7712 7590 7764 7642
rect 7776 7590 7828 7642
rect 7840 7590 7892 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 34315 7590 34367 7642
rect 34379 7590 34431 7642
rect 34443 7590 34495 7642
rect 34507 7590 34559 7642
rect 3148 7531 3200 7540
rect 3148 7497 3157 7531
rect 3157 7497 3191 7531
rect 3191 7497 3200 7531
rect 3148 7488 3200 7497
rect 4068 7488 4120 7540
rect 6184 7531 6236 7540
rect 6184 7497 6193 7531
rect 6193 7497 6227 7531
rect 6227 7497 6236 7531
rect 6184 7488 6236 7497
rect 6920 7488 6972 7540
rect 7472 7488 7524 7540
rect 10232 7488 10284 7540
rect 13820 7488 13872 7540
rect 16304 7488 16356 7540
rect 20812 7488 20864 7540
rect 23480 7531 23532 7540
rect 7012 7420 7064 7472
rect 7380 7420 7432 7472
rect 10692 7463 10744 7472
rect 10692 7429 10701 7463
rect 10701 7429 10735 7463
rect 10735 7429 10744 7463
rect 10692 7420 10744 7429
rect 11520 7420 11572 7472
rect 1492 7148 1544 7200
rect 1860 7284 1912 7336
rect 2412 7284 2464 7336
rect 2964 7216 3016 7268
rect 3976 7216 4028 7268
rect 3884 7148 3936 7200
rect 6736 7284 6788 7336
rect 8116 7284 8168 7336
rect 10784 7284 10836 7336
rect 15660 7420 15712 7472
rect 16212 7463 16264 7472
rect 16212 7429 16221 7463
rect 16221 7429 16255 7463
rect 16255 7429 16264 7463
rect 16212 7420 16264 7429
rect 17224 7420 17276 7472
rect 19616 7463 19668 7472
rect 19616 7429 19625 7463
rect 19625 7429 19659 7463
rect 19659 7429 19668 7463
rect 19616 7420 19668 7429
rect 16580 7395 16632 7404
rect 16580 7361 16589 7395
rect 16589 7361 16623 7395
rect 16623 7361 16632 7395
rect 16580 7352 16632 7361
rect 16764 7395 16816 7404
rect 16764 7361 16773 7395
rect 16773 7361 16807 7395
rect 16807 7361 16816 7395
rect 16764 7352 16816 7361
rect 19432 7395 19484 7404
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 20628 7352 20680 7404
rect 23480 7497 23489 7531
rect 23489 7497 23523 7531
rect 23523 7497 23532 7531
rect 23480 7488 23532 7497
rect 24584 7488 24636 7540
rect 25964 7531 26016 7540
rect 25964 7497 25973 7531
rect 25973 7497 26007 7531
rect 26007 7497 26016 7531
rect 28080 7531 28132 7540
rect 25964 7488 26016 7497
rect 28080 7497 28089 7531
rect 28089 7497 28123 7531
rect 28123 7497 28132 7531
rect 28080 7488 28132 7497
rect 28724 7531 28776 7540
rect 28724 7497 28733 7531
rect 28733 7497 28767 7531
rect 28767 7497 28776 7531
rect 28724 7488 28776 7497
rect 27160 7463 27212 7472
rect 27160 7429 27169 7463
rect 27169 7429 27203 7463
rect 27203 7429 27212 7463
rect 27160 7420 27212 7429
rect 33048 7488 33100 7540
rect 33232 7488 33284 7540
rect 33784 7488 33836 7540
rect 35900 7488 35952 7540
rect 34980 7463 35032 7472
rect 34980 7429 34989 7463
rect 34989 7429 35023 7463
rect 35023 7429 35032 7463
rect 34980 7420 35032 7429
rect 36084 7420 36136 7472
rect 21088 7395 21140 7404
rect 21088 7361 21097 7395
rect 21097 7361 21131 7395
rect 21131 7361 21140 7395
rect 21088 7352 21140 7361
rect 29000 7352 29052 7404
rect 32312 7395 32364 7404
rect 32312 7361 32321 7395
rect 32321 7361 32355 7395
rect 32355 7361 32364 7395
rect 32312 7352 32364 7361
rect 36544 7352 36596 7404
rect 15476 7327 15528 7336
rect 4712 7216 4764 7268
rect 7748 7259 7800 7268
rect 7748 7225 7782 7259
rect 7782 7225 7800 7259
rect 7748 7216 7800 7225
rect 10968 7259 11020 7268
rect 10968 7225 10977 7259
rect 10977 7225 11011 7259
rect 11011 7225 11020 7259
rect 10968 7216 11020 7225
rect 11152 7259 11204 7268
rect 11152 7225 11161 7259
rect 11161 7225 11195 7259
rect 11195 7225 11204 7259
rect 11152 7216 11204 7225
rect 5632 7191 5684 7200
rect 5632 7157 5641 7191
rect 5641 7157 5675 7191
rect 5675 7157 5684 7191
rect 5632 7148 5684 7157
rect 9588 7148 9640 7200
rect 10324 7148 10376 7200
rect 10416 7191 10468 7200
rect 10416 7157 10425 7191
rect 10425 7157 10459 7191
rect 10459 7157 10468 7191
rect 15476 7293 15485 7327
rect 15485 7293 15519 7327
rect 15519 7293 15528 7327
rect 15476 7284 15528 7293
rect 24584 7327 24636 7336
rect 24584 7293 24593 7327
rect 24593 7293 24627 7327
rect 24627 7293 24636 7327
rect 24584 7284 24636 7293
rect 24676 7284 24728 7336
rect 25412 7284 25464 7336
rect 30104 7284 30156 7336
rect 34888 7284 34940 7336
rect 35348 7284 35400 7336
rect 36636 7284 36688 7336
rect 11980 7216 12032 7268
rect 12900 7216 12952 7268
rect 16672 7259 16724 7268
rect 16672 7225 16681 7259
rect 16681 7225 16715 7259
rect 16715 7225 16724 7259
rect 16672 7216 16724 7225
rect 20168 7259 20220 7268
rect 10416 7148 10468 7157
rect 17316 7148 17368 7200
rect 18236 7148 18288 7200
rect 20168 7225 20177 7259
rect 20177 7225 20211 7259
rect 20211 7225 20220 7259
rect 20168 7216 20220 7225
rect 21180 7216 21232 7268
rect 22928 7216 22980 7268
rect 27252 7216 27304 7268
rect 27988 7216 28040 7268
rect 33048 7216 33100 7268
rect 35532 7259 35584 7268
rect 35532 7225 35541 7259
rect 35541 7225 35575 7259
rect 35575 7225 35584 7259
rect 35532 7216 35584 7225
rect 36452 7216 36504 7268
rect 37004 7259 37056 7268
rect 37004 7225 37013 7259
rect 37013 7225 37047 7259
rect 37047 7225 37056 7259
rect 37004 7216 37056 7225
rect 20628 7148 20680 7200
rect 22468 7191 22520 7200
rect 22468 7157 22477 7191
rect 22477 7157 22511 7191
rect 22511 7157 22520 7191
rect 22468 7148 22520 7157
rect 23112 7191 23164 7200
rect 23112 7157 23121 7191
rect 23121 7157 23155 7191
rect 23155 7157 23164 7191
rect 23112 7148 23164 7157
rect 24584 7148 24636 7200
rect 24768 7148 24820 7200
rect 26884 7191 26936 7200
rect 26884 7157 26893 7191
rect 26893 7157 26927 7191
rect 26927 7157 26936 7191
rect 26884 7148 26936 7157
rect 30656 7191 30708 7200
rect 30656 7157 30665 7191
rect 30665 7157 30699 7191
rect 30699 7157 30708 7191
rect 30656 7148 30708 7157
rect 33692 7148 33744 7200
rect 33968 7148 34020 7200
rect 34336 7191 34388 7200
rect 34336 7157 34345 7191
rect 34345 7157 34379 7191
rect 34379 7157 34388 7191
rect 34336 7148 34388 7157
rect 34704 7191 34756 7200
rect 34704 7157 34713 7191
rect 34713 7157 34747 7191
rect 34747 7157 34756 7191
rect 34704 7148 34756 7157
rect 35992 7148 36044 7200
rect 36636 7148 36688 7200
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 27648 7046 27700 7098
rect 27712 7046 27764 7098
rect 27776 7046 27828 7098
rect 27840 7046 27892 7098
rect 2412 6944 2464 6996
rect 3056 6944 3108 6996
rect 6736 6987 6788 6996
rect 6736 6953 6745 6987
rect 6745 6953 6779 6987
rect 6779 6953 6788 6987
rect 6736 6944 6788 6953
rect 10140 6944 10192 6996
rect 10692 6944 10744 6996
rect 11796 6944 11848 6996
rect 16764 6944 16816 6996
rect 17408 6944 17460 6996
rect 21180 6987 21232 6996
rect 21180 6953 21189 6987
rect 21189 6953 21223 6987
rect 21223 6953 21232 6987
rect 21180 6944 21232 6953
rect 23940 6944 23992 6996
rect 24676 6987 24728 6996
rect 24676 6953 24685 6987
rect 24685 6953 24719 6987
rect 24719 6953 24728 6987
rect 24676 6944 24728 6953
rect 25964 6987 26016 6996
rect 25964 6953 25973 6987
rect 25973 6953 26007 6987
rect 26007 6953 26016 6987
rect 25964 6944 26016 6953
rect 3332 6876 3384 6928
rect 3976 6876 4028 6928
rect 6276 6876 6328 6928
rect 7012 6876 7064 6928
rect 7564 6876 7616 6928
rect 9772 6876 9824 6928
rect 1492 6851 1544 6860
rect 1492 6817 1501 6851
rect 1501 6817 1535 6851
rect 1535 6817 1544 6851
rect 1492 6808 1544 6817
rect 1768 6851 1820 6860
rect 1768 6817 1802 6851
rect 1802 6817 1820 6851
rect 1768 6808 1820 6817
rect 3792 6808 3844 6860
rect 5080 6808 5132 6860
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 5816 6740 5868 6792
rect 5908 6740 5960 6792
rect 7748 6740 7800 6792
rect 10784 6808 10836 6860
rect 11060 6808 11112 6860
rect 12164 6808 12216 6860
rect 12992 6808 13044 6860
rect 21088 6876 21140 6928
rect 22100 6876 22152 6928
rect 16488 6808 16540 6860
rect 17408 6808 17460 6860
rect 23112 6876 23164 6928
rect 22376 6808 22428 6860
rect 24216 6851 24268 6860
rect 24216 6817 24225 6851
rect 24225 6817 24259 6851
rect 24259 6817 24268 6851
rect 24216 6808 24268 6817
rect 25228 6808 25280 6860
rect 27252 6944 27304 6996
rect 32312 6987 32364 6996
rect 32312 6953 32321 6987
rect 32321 6953 32355 6987
rect 32355 6953 32364 6987
rect 32312 6944 32364 6953
rect 33784 6987 33836 6996
rect 33784 6953 33793 6987
rect 33793 6953 33827 6987
rect 33827 6953 33836 6987
rect 33784 6944 33836 6953
rect 26792 6808 26844 6860
rect 27068 6808 27120 6860
rect 29092 6876 29144 6928
rect 29184 6808 29236 6860
rect 29368 6851 29420 6860
rect 29368 6817 29391 6851
rect 29391 6817 29420 6851
rect 30656 6876 30708 6928
rect 29368 6808 29420 6817
rect 33140 6808 33192 6860
rect 33600 6876 33652 6928
rect 34888 6919 34940 6928
rect 34888 6885 34897 6919
rect 34897 6885 34931 6919
rect 34931 6885 34940 6919
rect 34888 6876 34940 6885
rect 36084 6876 36136 6928
rect 36360 6876 36412 6928
rect 34060 6808 34112 6860
rect 34336 6808 34388 6860
rect 35532 6808 35584 6860
rect 9588 6740 9640 6792
rect 9864 6740 9916 6792
rect 11152 6740 11204 6792
rect 4160 6672 4212 6724
rect 5724 6672 5776 6724
rect 11980 6783 12032 6792
rect 11980 6749 11989 6783
rect 11989 6749 12023 6783
rect 12023 6749 12032 6783
rect 13360 6783 13412 6792
rect 11980 6740 12032 6749
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 15108 6740 15160 6792
rect 15660 6740 15712 6792
rect 18236 6783 18288 6792
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 25412 6783 25464 6792
rect 25412 6749 25421 6783
rect 25421 6749 25455 6783
rect 25455 6749 25464 6783
rect 25412 6740 25464 6749
rect 25504 6783 25556 6792
rect 25504 6749 25513 6783
rect 25513 6749 25547 6783
rect 25547 6749 25556 6783
rect 25504 6740 25556 6749
rect 27804 6740 27856 6792
rect 29000 6740 29052 6792
rect 33692 6740 33744 6792
rect 34152 6740 34204 6792
rect 35072 6740 35124 6792
rect 36360 6783 36412 6792
rect 36360 6749 36369 6783
rect 36369 6749 36403 6783
rect 36403 6749 36412 6783
rect 36360 6740 36412 6749
rect 11520 6672 11572 6724
rect 24952 6715 25004 6724
rect 24952 6681 24961 6715
rect 24961 6681 24995 6715
rect 24995 6681 25004 6715
rect 24952 6672 25004 6681
rect 30932 6672 30984 6724
rect 3884 6604 3936 6656
rect 5448 6647 5500 6656
rect 5448 6613 5457 6647
rect 5457 6613 5491 6647
rect 5491 6613 5500 6647
rect 5448 6604 5500 6613
rect 9680 6604 9732 6656
rect 11336 6604 11388 6656
rect 12624 6647 12676 6656
rect 12624 6613 12633 6647
rect 12633 6613 12667 6647
rect 12667 6613 12676 6647
rect 12624 6604 12676 6613
rect 15384 6604 15436 6656
rect 17592 6604 17644 6656
rect 18512 6604 18564 6656
rect 26608 6647 26660 6656
rect 26608 6613 26617 6647
rect 26617 6613 26651 6647
rect 26651 6613 26660 6647
rect 26608 6604 26660 6613
rect 27896 6647 27948 6656
rect 27896 6613 27905 6647
rect 27905 6613 27939 6647
rect 27939 6613 27948 6647
rect 27896 6604 27948 6613
rect 30472 6647 30524 6656
rect 30472 6613 30481 6647
rect 30481 6613 30515 6647
rect 30515 6613 30524 6647
rect 30472 6604 30524 6613
rect 33876 6604 33928 6656
rect 35256 6604 35308 6656
rect 35992 6647 36044 6656
rect 35992 6613 36001 6647
rect 36001 6613 36035 6647
rect 36035 6613 36044 6647
rect 35992 6604 36044 6613
rect 36544 6604 36596 6656
rect 7648 6502 7700 6554
rect 7712 6502 7764 6554
rect 7776 6502 7828 6554
rect 7840 6502 7892 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 34315 6502 34367 6554
rect 34379 6502 34431 6554
rect 34443 6502 34495 6554
rect 34507 6502 34559 6554
rect 1400 6400 1452 6452
rect 2596 6400 2648 6452
rect 3792 6400 3844 6452
rect 5080 6443 5132 6452
rect 5080 6409 5089 6443
rect 5089 6409 5123 6443
rect 5123 6409 5132 6443
rect 5080 6400 5132 6409
rect 6276 6443 6328 6452
rect 6276 6409 6285 6443
rect 6285 6409 6319 6443
rect 6319 6409 6328 6443
rect 6276 6400 6328 6409
rect 6644 6443 6696 6452
rect 6644 6409 6653 6443
rect 6653 6409 6687 6443
rect 6687 6409 6696 6443
rect 6644 6400 6696 6409
rect 7012 6400 7064 6452
rect 8116 6400 8168 6452
rect 9772 6400 9824 6452
rect 10140 6443 10192 6452
rect 10140 6409 10149 6443
rect 10149 6409 10183 6443
rect 10183 6409 10192 6443
rect 10140 6400 10192 6409
rect 11796 6443 11848 6452
rect 11796 6409 11805 6443
rect 11805 6409 11839 6443
rect 11839 6409 11848 6443
rect 11796 6400 11848 6409
rect 12164 6443 12216 6452
rect 12164 6409 12173 6443
rect 12173 6409 12207 6443
rect 12207 6409 12216 6443
rect 12164 6400 12216 6409
rect 13544 6400 13596 6452
rect 17408 6443 17460 6452
rect 17408 6409 17417 6443
rect 17417 6409 17451 6443
rect 17451 6409 17460 6443
rect 17408 6400 17460 6409
rect 18236 6400 18288 6452
rect 6000 6332 6052 6384
rect 11060 6332 11112 6384
rect 14004 6375 14056 6384
rect 14004 6341 14013 6375
rect 14013 6341 14047 6375
rect 14047 6341 14056 6375
rect 14004 6332 14056 6341
rect 18144 6375 18196 6384
rect 18144 6341 18153 6375
rect 18153 6341 18187 6375
rect 18187 6341 18196 6375
rect 18144 6332 18196 6341
rect 5448 6264 5500 6316
rect 3792 6196 3844 6248
rect 5816 6239 5868 6248
rect 5816 6205 5825 6239
rect 5825 6205 5859 6239
rect 5859 6205 5868 6239
rect 5816 6196 5868 6205
rect 6736 6196 6788 6248
rect 9864 6264 9916 6316
rect 10048 6264 10100 6316
rect 11520 6264 11572 6316
rect 12624 6307 12676 6316
rect 12624 6273 12633 6307
rect 12633 6273 12667 6307
rect 12667 6273 12676 6307
rect 12624 6264 12676 6273
rect 22100 6400 22152 6452
rect 22376 6400 22428 6452
rect 23112 6443 23164 6452
rect 23112 6409 23121 6443
rect 23121 6409 23155 6443
rect 23155 6409 23164 6443
rect 23112 6400 23164 6409
rect 23940 6443 23992 6452
rect 23940 6409 23949 6443
rect 23949 6409 23983 6443
rect 23983 6409 23992 6443
rect 23940 6400 23992 6409
rect 24124 6443 24176 6452
rect 24124 6409 24133 6443
rect 24133 6409 24167 6443
rect 24167 6409 24176 6443
rect 24124 6400 24176 6409
rect 25412 6400 25464 6452
rect 27068 6400 27120 6452
rect 28632 6400 28684 6452
rect 29000 6443 29052 6452
rect 29000 6409 29009 6443
rect 29009 6409 29043 6443
rect 29043 6409 29052 6443
rect 29000 6400 29052 6409
rect 33140 6400 33192 6452
rect 34060 6443 34112 6452
rect 34060 6409 34069 6443
rect 34069 6409 34103 6443
rect 34103 6409 34112 6443
rect 34060 6400 34112 6409
rect 36544 6400 36596 6452
rect 27804 6332 27856 6384
rect 30196 6332 30248 6384
rect 33600 6332 33652 6384
rect 10784 6196 10836 6248
rect 11428 6239 11480 6248
rect 11428 6205 11437 6239
rect 11437 6205 11471 6239
rect 11471 6205 11480 6239
rect 11428 6196 11480 6205
rect 15108 6239 15160 6248
rect 15108 6205 15117 6239
rect 15117 6205 15151 6239
rect 15151 6205 15160 6239
rect 15108 6196 15160 6205
rect 24492 6307 24544 6316
rect 24492 6273 24501 6307
rect 24501 6273 24535 6307
rect 24535 6273 24544 6307
rect 24492 6264 24544 6273
rect 24676 6307 24728 6316
rect 24676 6273 24685 6307
rect 24685 6273 24719 6307
rect 24719 6273 24728 6307
rect 24676 6264 24728 6273
rect 25228 6264 25280 6316
rect 29828 6307 29880 6316
rect 29828 6273 29837 6307
rect 29837 6273 29871 6307
rect 29871 6273 29880 6307
rect 29828 6264 29880 6273
rect 33232 6264 33284 6316
rect 34888 6264 34940 6316
rect 35072 6307 35124 6316
rect 35072 6273 35081 6307
rect 35081 6273 35115 6307
rect 35115 6273 35124 6307
rect 35072 6264 35124 6273
rect 15384 6239 15436 6248
rect 15384 6205 15407 6239
rect 15407 6205 15436 6239
rect 15384 6196 15436 6205
rect 24860 6196 24912 6248
rect 25688 6196 25740 6248
rect 29920 6239 29972 6248
rect 29920 6205 29929 6239
rect 29929 6205 29963 6239
rect 29963 6205 29972 6239
rect 29920 6196 29972 6205
rect 32312 6196 32364 6248
rect 34060 6196 34112 6248
rect 34612 6196 34664 6248
rect 35256 6239 35308 6248
rect 35256 6205 35265 6239
rect 35265 6205 35299 6239
rect 35299 6205 35308 6239
rect 35256 6196 35308 6205
rect 35532 6239 35584 6248
rect 35532 6205 35566 6239
rect 35566 6205 35584 6239
rect 35532 6196 35584 6205
rect 1768 6128 1820 6180
rect 3056 6128 3108 6180
rect 5724 6171 5776 6180
rect 5724 6137 5733 6171
rect 5733 6137 5767 6171
rect 5767 6137 5776 6171
rect 5724 6128 5776 6137
rect 7012 6128 7064 6180
rect 11336 6171 11388 6180
rect 11336 6137 11345 6171
rect 11345 6137 11379 6171
rect 11379 6137 11388 6171
rect 11336 6128 11388 6137
rect 12532 6128 12584 6180
rect 13544 6128 13596 6180
rect 18420 6171 18472 6180
rect 18420 6137 18429 6171
rect 18429 6137 18463 6171
rect 18463 6137 18472 6171
rect 18420 6128 18472 6137
rect 18604 6171 18656 6180
rect 18604 6137 18613 6171
rect 18613 6137 18647 6171
rect 18647 6137 18656 6171
rect 18604 6128 18656 6137
rect 18696 6171 18748 6180
rect 18696 6137 18705 6171
rect 18705 6137 18739 6171
rect 18739 6137 18748 6171
rect 18696 6128 18748 6137
rect 21732 6128 21784 6180
rect 24584 6171 24636 6180
rect 24584 6137 24593 6171
rect 24593 6137 24627 6171
rect 24627 6137 24636 6171
rect 24584 6128 24636 6137
rect 25964 6128 26016 6180
rect 28908 6128 28960 6180
rect 30748 6128 30800 6180
rect 3976 6103 4028 6112
rect 3976 6069 3985 6103
rect 3985 6069 4019 6103
rect 4019 6069 4028 6103
rect 3976 6060 4028 6069
rect 8024 6060 8076 6112
rect 16488 6103 16540 6112
rect 16488 6069 16497 6103
rect 16497 6069 16531 6103
rect 16531 6069 16540 6103
rect 16488 6060 16540 6069
rect 17684 6060 17736 6112
rect 26976 6103 27028 6112
rect 26976 6069 26985 6103
rect 26985 6069 27019 6103
rect 27019 6069 27028 6103
rect 26976 6060 27028 6069
rect 29736 6060 29788 6112
rect 32128 6060 32180 6112
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 27648 5958 27700 6010
rect 27712 5958 27764 6010
rect 27776 5958 27828 6010
rect 27840 5958 27892 6010
rect 4436 5856 4488 5908
rect 5908 5856 5960 5908
rect 6092 5899 6144 5908
rect 6092 5865 6101 5899
rect 6101 5865 6135 5899
rect 6135 5865 6144 5899
rect 6092 5856 6144 5865
rect 7104 5856 7156 5908
rect 10048 5899 10100 5908
rect 10048 5865 10057 5899
rect 10057 5865 10091 5899
rect 10091 5865 10100 5899
rect 10048 5856 10100 5865
rect 11336 5856 11388 5908
rect 12440 5899 12492 5908
rect 12440 5865 12449 5899
rect 12449 5865 12483 5899
rect 12483 5865 12492 5899
rect 12992 5899 13044 5908
rect 12440 5856 12492 5865
rect 12992 5865 13001 5899
rect 13001 5865 13035 5899
rect 13035 5865 13044 5899
rect 12992 5856 13044 5865
rect 13360 5899 13412 5908
rect 13360 5865 13369 5899
rect 13369 5865 13403 5899
rect 13403 5865 13412 5899
rect 13360 5856 13412 5865
rect 15660 5856 15712 5908
rect 16672 5899 16724 5908
rect 16672 5865 16681 5899
rect 16681 5865 16715 5899
rect 16715 5865 16724 5899
rect 16672 5856 16724 5865
rect 17316 5856 17368 5908
rect 21640 5899 21692 5908
rect 21640 5865 21649 5899
rect 21649 5865 21683 5899
rect 21683 5865 21692 5899
rect 21640 5856 21692 5865
rect 22376 5899 22428 5908
rect 22376 5865 22385 5899
rect 22385 5865 22419 5899
rect 22419 5865 22428 5899
rect 22376 5856 22428 5865
rect 25504 5856 25556 5908
rect 26792 5899 26844 5908
rect 26792 5865 26801 5899
rect 26801 5865 26835 5899
rect 26835 5865 26844 5899
rect 26792 5856 26844 5865
rect 27436 5899 27488 5908
rect 27436 5865 27445 5899
rect 27445 5865 27479 5899
rect 27479 5865 27488 5899
rect 27436 5856 27488 5865
rect 29828 5899 29880 5908
rect 29828 5865 29837 5899
rect 29837 5865 29871 5899
rect 29871 5865 29880 5899
rect 29828 5856 29880 5865
rect 30380 5856 30432 5908
rect 33140 5899 33192 5908
rect 33140 5865 33149 5899
rect 33149 5865 33183 5899
rect 33183 5865 33192 5899
rect 33140 5856 33192 5865
rect 33876 5856 33928 5908
rect 35532 5899 35584 5908
rect 35532 5865 35541 5899
rect 35541 5865 35575 5899
rect 35575 5865 35584 5899
rect 35532 5856 35584 5865
rect 36084 5899 36136 5908
rect 36084 5865 36093 5899
rect 36093 5865 36127 5899
rect 36127 5865 36136 5899
rect 36084 5856 36136 5865
rect 2872 5788 2924 5840
rect 3976 5788 4028 5840
rect 4988 5788 5040 5840
rect 8024 5788 8076 5840
rect 10140 5788 10192 5840
rect 10784 5831 10836 5840
rect 10784 5797 10793 5831
rect 10793 5797 10827 5831
rect 10827 5797 10836 5831
rect 12256 5831 12308 5840
rect 10784 5788 10836 5797
rect 12256 5797 12265 5831
rect 12265 5797 12299 5831
rect 12299 5797 12308 5831
rect 12256 5788 12308 5797
rect 12532 5831 12584 5840
rect 12532 5797 12541 5831
rect 12541 5797 12575 5831
rect 12575 5797 12584 5831
rect 14004 5831 14056 5840
rect 12532 5788 12584 5797
rect 14004 5797 14013 5831
rect 14013 5797 14047 5831
rect 14047 5797 14056 5831
rect 14004 5788 14056 5797
rect 14188 5831 14240 5840
rect 14188 5797 14197 5831
rect 14197 5797 14231 5831
rect 14231 5797 14240 5831
rect 14188 5788 14240 5797
rect 2412 5720 2464 5772
rect 4068 5763 4120 5772
rect 2136 5652 2188 5704
rect 3056 5652 3108 5704
rect 4068 5729 4077 5763
rect 4077 5729 4111 5763
rect 4111 5729 4120 5763
rect 4068 5720 4120 5729
rect 5632 5720 5684 5772
rect 7012 5720 7064 5772
rect 10508 5763 10560 5772
rect 10508 5729 10517 5763
rect 10517 5729 10551 5763
rect 10551 5729 10560 5763
rect 10508 5720 10560 5729
rect 11980 5720 12032 5772
rect 13820 5720 13872 5772
rect 15108 5788 15160 5840
rect 16764 5831 16816 5840
rect 16764 5797 16773 5831
rect 16773 5797 16807 5831
rect 16807 5797 16816 5831
rect 18052 5831 18104 5840
rect 16764 5788 16816 5797
rect 18052 5797 18061 5831
rect 18061 5797 18095 5831
rect 18095 5797 18104 5831
rect 18052 5788 18104 5797
rect 18236 5831 18288 5840
rect 18236 5797 18245 5831
rect 18245 5797 18279 5831
rect 18279 5797 18288 5831
rect 18236 5788 18288 5797
rect 21732 5831 21784 5840
rect 21732 5797 21741 5831
rect 21741 5797 21775 5831
rect 21775 5797 21784 5831
rect 21732 5788 21784 5797
rect 22468 5788 22520 5840
rect 21456 5720 21508 5772
rect 4528 5652 4580 5704
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 6736 5652 6788 5704
rect 16396 5652 16448 5704
rect 16856 5652 16908 5704
rect 19800 5695 19852 5704
rect 6828 5584 6880 5636
rect 13728 5627 13780 5636
rect 13728 5593 13737 5627
rect 13737 5593 13771 5627
rect 13771 5593 13780 5627
rect 13728 5584 13780 5593
rect 1768 5516 1820 5568
rect 2136 5559 2188 5568
rect 2136 5525 2145 5559
rect 2145 5525 2179 5559
rect 2179 5525 2188 5559
rect 2136 5516 2188 5525
rect 2688 5516 2740 5568
rect 3148 5516 3200 5568
rect 4896 5516 4948 5568
rect 9496 5516 9548 5568
rect 10232 5559 10284 5568
rect 10232 5525 10241 5559
rect 10241 5525 10275 5559
rect 10275 5525 10284 5559
rect 10232 5516 10284 5525
rect 16212 5559 16264 5568
rect 16212 5525 16221 5559
rect 16221 5525 16255 5559
rect 16255 5525 16264 5559
rect 16212 5516 16264 5525
rect 16580 5516 16632 5568
rect 19800 5661 19809 5695
rect 19809 5661 19843 5695
rect 19843 5661 19852 5695
rect 19800 5652 19852 5661
rect 20812 5652 20864 5704
rect 21824 5720 21876 5772
rect 22008 5720 22060 5772
rect 23112 5788 23164 5840
rect 29184 5788 29236 5840
rect 29368 5788 29420 5840
rect 33048 5788 33100 5840
rect 33232 5831 33284 5840
rect 33232 5797 33241 5831
rect 33241 5797 33275 5831
rect 33275 5797 33284 5831
rect 33232 5788 33284 5797
rect 33692 5831 33744 5840
rect 33692 5797 33701 5831
rect 33701 5797 33735 5831
rect 33735 5797 33744 5831
rect 33692 5788 33744 5797
rect 34152 5788 34204 5840
rect 22928 5763 22980 5772
rect 22928 5729 22962 5763
rect 22962 5729 22980 5763
rect 22928 5720 22980 5729
rect 26976 5720 27028 5772
rect 27712 5720 27764 5772
rect 28448 5720 28500 5772
rect 24860 5652 24912 5704
rect 27436 5695 27488 5704
rect 27436 5661 27445 5695
rect 27445 5661 27479 5695
rect 27479 5661 27488 5695
rect 27436 5652 27488 5661
rect 28172 5652 28224 5704
rect 29000 5652 29052 5704
rect 30748 5720 30800 5772
rect 30472 5695 30524 5704
rect 30472 5661 30481 5695
rect 30481 5661 30515 5695
rect 30515 5661 30524 5695
rect 30472 5652 30524 5661
rect 34060 5652 34112 5704
rect 20720 5584 20772 5636
rect 26056 5627 26108 5636
rect 26056 5593 26065 5627
rect 26065 5593 26099 5627
rect 26099 5593 26108 5627
rect 26056 5584 26108 5593
rect 31852 5584 31904 5636
rect 35900 5584 35952 5636
rect 36360 5584 36412 5636
rect 18696 5559 18748 5568
rect 18696 5525 18705 5559
rect 18705 5525 18739 5559
rect 18739 5525 18748 5559
rect 18696 5516 18748 5525
rect 24308 5516 24360 5568
rect 25688 5559 25740 5568
rect 25688 5525 25697 5559
rect 25697 5525 25731 5559
rect 25731 5525 25740 5559
rect 25688 5516 25740 5525
rect 26148 5516 26200 5568
rect 30104 5559 30156 5568
rect 30104 5525 30113 5559
rect 30113 5525 30147 5559
rect 30147 5525 30156 5559
rect 30104 5516 30156 5525
rect 7648 5414 7700 5466
rect 7712 5414 7764 5466
rect 7776 5414 7828 5466
rect 7840 5414 7892 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 34315 5414 34367 5466
rect 34379 5414 34431 5466
rect 34443 5414 34495 5466
rect 34507 5414 34559 5466
rect 1676 5312 1728 5364
rect 2228 5312 2280 5364
rect 2412 5312 2464 5364
rect 2872 5355 2924 5364
rect 2872 5321 2881 5355
rect 2881 5321 2915 5355
rect 2915 5321 2924 5355
rect 2872 5312 2924 5321
rect 4344 5312 4396 5364
rect 5632 5355 5684 5364
rect 5632 5321 5641 5355
rect 5641 5321 5675 5355
rect 5675 5321 5684 5355
rect 5632 5312 5684 5321
rect 6552 5355 6604 5364
rect 6552 5321 6561 5355
rect 6561 5321 6595 5355
rect 6595 5321 6604 5355
rect 10876 5355 10928 5364
rect 6552 5312 6604 5321
rect 6736 5244 6788 5296
rect 7380 5287 7432 5296
rect 7380 5253 7389 5287
rect 7389 5253 7423 5287
rect 7423 5253 7432 5287
rect 7380 5244 7432 5253
rect 4988 5219 5040 5228
rect 4988 5185 4997 5219
rect 4997 5185 5031 5219
rect 5031 5185 5040 5219
rect 4988 5176 5040 5185
rect 10876 5321 10885 5355
rect 10885 5321 10919 5355
rect 10919 5321 10928 5355
rect 10876 5312 10928 5321
rect 12256 5312 12308 5364
rect 12532 5312 12584 5364
rect 13728 5355 13780 5364
rect 13728 5321 13737 5355
rect 13737 5321 13771 5355
rect 13771 5321 13780 5355
rect 13728 5312 13780 5321
rect 14188 5312 14240 5364
rect 16764 5312 16816 5364
rect 17408 5355 17460 5364
rect 17408 5321 17417 5355
rect 17417 5321 17451 5355
rect 17451 5321 17460 5355
rect 17408 5312 17460 5321
rect 17776 5355 17828 5364
rect 17776 5321 17785 5355
rect 17785 5321 17819 5355
rect 17819 5321 17828 5355
rect 17776 5312 17828 5321
rect 19524 5355 19576 5364
rect 19524 5321 19533 5355
rect 19533 5321 19567 5355
rect 19567 5321 19576 5355
rect 19524 5312 19576 5321
rect 20812 5355 20864 5364
rect 20812 5321 20821 5355
rect 20821 5321 20855 5355
rect 20855 5321 20864 5355
rect 20812 5312 20864 5321
rect 21548 5312 21600 5364
rect 22468 5312 22520 5364
rect 23112 5312 23164 5364
rect 23204 5312 23256 5364
rect 9404 5244 9456 5296
rect 10784 5244 10836 5296
rect 14004 5244 14056 5296
rect 16396 5244 16448 5296
rect 11428 5219 11480 5228
rect 11428 5185 11437 5219
rect 11437 5185 11471 5219
rect 11471 5185 11480 5219
rect 11428 5176 11480 5185
rect 13360 5176 13412 5228
rect 15844 5176 15896 5228
rect 17316 5176 17368 5228
rect 18144 5287 18196 5296
rect 18144 5253 18153 5287
rect 18153 5253 18187 5287
rect 18187 5253 18196 5287
rect 18144 5244 18196 5253
rect 20352 5244 20404 5296
rect 21180 5244 21232 5296
rect 21364 5287 21416 5296
rect 21364 5253 21373 5287
rect 21373 5253 21407 5287
rect 21407 5253 21416 5287
rect 21364 5244 21416 5253
rect 21824 5244 21876 5296
rect 24492 5312 24544 5364
rect 25596 5355 25648 5364
rect 25596 5321 25605 5355
rect 25605 5321 25639 5355
rect 25639 5321 25648 5355
rect 25596 5312 25648 5321
rect 26608 5355 26660 5364
rect 26608 5321 26617 5355
rect 26617 5321 26651 5355
rect 26651 5321 26660 5355
rect 26608 5312 26660 5321
rect 27344 5312 27396 5364
rect 28172 5355 28224 5364
rect 28172 5321 28181 5355
rect 28181 5321 28215 5355
rect 28215 5321 28224 5355
rect 28172 5312 28224 5321
rect 30380 5312 30432 5364
rect 30932 5355 30984 5364
rect 30932 5321 30941 5355
rect 30941 5321 30975 5355
rect 30975 5321 30984 5355
rect 30932 5312 30984 5321
rect 33048 5312 33100 5364
rect 35624 5355 35676 5364
rect 35624 5321 35633 5355
rect 35633 5321 35667 5355
rect 35667 5321 35676 5355
rect 35624 5312 35676 5321
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 24216 5219 24268 5228
rect 24216 5185 24225 5219
rect 24225 5185 24259 5219
rect 24259 5185 24268 5219
rect 24216 5176 24268 5185
rect 24768 5176 24820 5228
rect 26056 5219 26108 5228
rect 26056 5185 26065 5219
rect 26065 5185 26099 5219
rect 26099 5185 26108 5219
rect 26056 5176 26108 5185
rect 1676 5108 1728 5160
rect 3148 5151 3200 5160
rect 3148 5117 3157 5151
rect 3157 5117 3191 5151
rect 3191 5117 3200 5151
rect 3148 5108 3200 5117
rect 4160 5151 4212 5160
rect 4160 5117 4169 5151
rect 4169 5117 4203 5151
rect 4203 5117 4212 5151
rect 4160 5108 4212 5117
rect 5080 5108 5132 5160
rect 3424 5083 3476 5092
rect 3424 5049 3433 5083
rect 3433 5049 3467 5083
rect 3467 5049 3476 5083
rect 3424 5040 3476 5049
rect 3884 5040 3936 5092
rect 7932 5083 7984 5092
rect 7932 5049 7941 5083
rect 7941 5049 7975 5083
rect 7975 5049 7984 5083
rect 11060 5108 11112 5160
rect 19800 5108 19852 5160
rect 20260 5108 20312 5160
rect 21456 5108 21508 5160
rect 30288 5244 30340 5296
rect 27712 5219 27764 5228
rect 27712 5185 27721 5219
rect 27721 5185 27755 5219
rect 27755 5185 27764 5219
rect 27712 5176 27764 5185
rect 29920 5176 29972 5228
rect 32128 5176 32180 5228
rect 7932 5040 7984 5049
rect 8944 5040 8996 5092
rect 3148 4972 3200 5024
rect 3516 4972 3568 5024
rect 4896 5015 4948 5024
rect 4896 4981 4905 5015
rect 4905 4981 4939 5015
rect 4939 4981 4948 5015
rect 4896 4972 4948 4981
rect 6828 4972 6880 5024
rect 7288 4972 7340 5024
rect 8760 5015 8812 5024
rect 8760 4981 8769 5015
rect 8769 4981 8803 5015
rect 8803 4981 8812 5015
rect 9588 5040 9640 5092
rect 16212 5083 16264 5092
rect 16212 5049 16221 5083
rect 16221 5049 16255 5083
rect 16255 5049 16264 5083
rect 16212 5040 16264 5049
rect 18604 5083 18656 5092
rect 8760 4972 8812 4981
rect 10876 4972 10928 5024
rect 16120 4972 16172 5024
rect 18604 5049 18613 5083
rect 18613 5049 18647 5083
rect 18647 5049 18656 5083
rect 18604 5040 18656 5049
rect 18696 5083 18748 5092
rect 18696 5049 18705 5083
rect 18705 5049 18739 5083
rect 18739 5049 18748 5083
rect 21916 5083 21968 5092
rect 18696 5040 18748 5049
rect 21916 5049 21925 5083
rect 21925 5049 21959 5083
rect 21959 5049 21968 5083
rect 21916 5040 21968 5049
rect 24308 5083 24360 5092
rect 24308 5049 24317 5083
rect 24317 5049 24351 5083
rect 24351 5049 24360 5083
rect 24308 5040 24360 5049
rect 25872 5040 25924 5092
rect 28632 5108 28684 5160
rect 29000 5108 29052 5160
rect 19524 4972 19576 5024
rect 20444 4972 20496 5024
rect 21824 5015 21876 5024
rect 21824 4981 21833 5015
rect 21833 4981 21867 5015
rect 21867 4981 21876 5015
rect 21824 4972 21876 4981
rect 23112 5015 23164 5024
rect 23112 4981 23121 5015
rect 23121 4981 23155 5015
rect 23155 4981 23164 5015
rect 23112 4972 23164 4981
rect 24124 4972 24176 5024
rect 27344 5040 27396 5092
rect 28448 5083 28500 5092
rect 28448 5049 28457 5083
rect 28457 5049 28491 5083
rect 28491 5049 28500 5083
rect 28448 5040 28500 5049
rect 29920 5083 29972 5092
rect 29920 5049 29929 5083
rect 29929 5049 29963 5083
rect 29963 5049 29972 5083
rect 29920 5040 29972 5049
rect 30104 5083 30156 5092
rect 30104 5049 30113 5083
rect 30113 5049 30147 5083
rect 30147 5049 30156 5083
rect 30104 5040 30156 5049
rect 34060 5108 34112 5160
rect 35440 5151 35492 5160
rect 35440 5117 35449 5151
rect 35449 5117 35483 5151
rect 35483 5117 35492 5151
rect 35440 5108 35492 5117
rect 34152 5040 34204 5092
rect 28540 4972 28592 5024
rect 30472 4972 30524 5024
rect 33692 5015 33744 5024
rect 33692 4981 33701 5015
rect 33701 4981 33735 5015
rect 33735 4981 33744 5015
rect 33692 4972 33744 4981
rect 34060 4972 34112 5024
rect 34980 4972 35032 5024
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 27648 4870 27700 4922
rect 27712 4870 27764 4922
rect 27776 4870 27828 4922
rect 27840 4870 27892 4922
rect 1676 4811 1728 4820
rect 1676 4777 1685 4811
rect 1685 4777 1719 4811
rect 1719 4777 1728 4811
rect 1676 4768 1728 4777
rect 2136 4811 2188 4820
rect 2136 4777 2145 4811
rect 2145 4777 2179 4811
rect 2179 4777 2188 4811
rect 2136 4768 2188 4777
rect 2780 4768 2832 4820
rect 3884 4811 3936 4820
rect 3884 4777 3893 4811
rect 3893 4777 3927 4811
rect 3927 4777 3936 4811
rect 3884 4768 3936 4777
rect 5724 4768 5776 4820
rect 7196 4768 7248 4820
rect 8208 4768 8260 4820
rect 10232 4768 10284 4820
rect 10876 4811 10928 4820
rect 10876 4777 10885 4811
rect 10885 4777 10919 4811
rect 10919 4777 10928 4811
rect 10876 4768 10928 4777
rect 11060 4768 11112 4820
rect 12348 4768 12400 4820
rect 16120 4768 16172 4820
rect 16396 4811 16448 4820
rect 16396 4777 16405 4811
rect 16405 4777 16439 4811
rect 16439 4777 16448 4811
rect 16396 4768 16448 4777
rect 17868 4768 17920 4820
rect 18604 4768 18656 4820
rect 20076 4768 20128 4820
rect 21824 4768 21876 4820
rect 23204 4768 23256 4820
rect 2964 4700 3016 4752
rect 7104 4700 7156 4752
rect 7472 4700 7524 4752
rect 18696 4700 18748 4752
rect 3424 4675 3476 4684
rect 3424 4641 3433 4675
rect 3433 4641 3467 4675
rect 3467 4641 3476 4675
rect 3424 4632 3476 4641
rect 4712 4632 4764 4684
rect 12532 4632 12584 4684
rect 15200 4632 15252 4684
rect 15844 4632 15896 4684
rect 2872 4607 2924 4616
rect 2872 4573 2881 4607
rect 2881 4573 2915 4607
rect 2915 4573 2924 4607
rect 2872 4564 2924 4573
rect 2412 4539 2464 4548
rect 2412 4505 2421 4539
rect 2421 4505 2455 4539
rect 2455 4505 2464 4539
rect 2412 4496 2464 4505
rect 2136 4428 2188 4480
rect 3056 4428 3108 4480
rect 3884 4564 3936 4616
rect 7932 4564 7984 4616
rect 10140 4607 10192 4616
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 16396 4607 16448 4616
rect 16396 4573 16405 4607
rect 16405 4573 16439 4607
rect 16439 4573 16448 4607
rect 16396 4564 16448 4573
rect 19800 4607 19852 4616
rect 19800 4573 19809 4607
rect 19809 4573 19843 4607
rect 19843 4573 19852 4607
rect 19800 4564 19852 4573
rect 20260 4564 20312 4616
rect 22928 4700 22980 4752
rect 25872 4811 25924 4820
rect 25872 4777 25881 4811
rect 25881 4777 25915 4811
rect 25915 4777 25924 4811
rect 25872 4768 25924 4777
rect 28632 4811 28684 4820
rect 28632 4777 28641 4811
rect 28641 4777 28675 4811
rect 28675 4777 28684 4811
rect 28632 4768 28684 4777
rect 29828 4768 29880 4820
rect 30196 4768 30248 4820
rect 30564 4768 30616 4820
rect 30748 4811 30800 4820
rect 30748 4777 30757 4811
rect 30757 4777 30791 4811
rect 30791 4777 30800 4811
rect 30748 4768 30800 4777
rect 32128 4768 32180 4820
rect 25320 4743 25372 4752
rect 25320 4709 25329 4743
rect 25329 4709 25363 4743
rect 25363 4709 25372 4743
rect 25320 4700 25372 4709
rect 21180 4632 21232 4684
rect 23112 4675 23164 4684
rect 23112 4641 23121 4675
rect 23121 4641 23155 4675
rect 23155 4641 23164 4675
rect 25136 4675 25188 4684
rect 23112 4632 23164 4641
rect 25136 4641 25145 4675
rect 25145 4641 25179 4675
rect 25179 4641 25188 4675
rect 25136 4632 25188 4641
rect 6644 4471 6696 4480
rect 6644 4437 6653 4471
rect 6653 4437 6687 4471
rect 6687 4437 6696 4471
rect 15752 4496 15804 4548
rect 20720 4496 20772 4548
rect 25780 4700 25832 4752
rect 27528 4743 27580 4752
rect 27528 4709 27562 4743
rect 27562 4709 27580 4743
rect 27528 4700 27580 4709
rect 30380 4743 30432 4752
rect 30380 4709 30389 4743
rect 30389 4709 30423 4743
rect 30423 4709 30432 4743
rect 30380 4700 30432 4709
rect 27344 4632 27396 4684
rect 33140 4768 33192 4820
rect 33416 4811 33468 4820
rect 33416 4777 33425 4811
rect 33425 4777 33459 4811
rect 33459 4777 33468 4811
rect 33416 4768 33468 4777
rect 33232 4743 33284 4752
rect 33232 4709 33241 4743
rect 33241 4709 33275 4743
rect 33275 4709 33284 4743
rect 33232 4700 33284 4709
rect 26240 4564 26292 4616
rect 26792 4564 26844 4616
rect 30288 4607 30340 4616
rect 30288 4573 30297 4607
rect 30297 4573 30331 4607
rect 30331 4573 30340 4607
rect 30288 4564 30340 4573
rect 24124 4496 24176 4548
rect 29644 4496 29696 4548
rect 32956 4539 33008 4548
rect 32956 4505 32965 4539
rect 32965 4505 32999 4539
rect 32999 4505 33008 4539
rect 32956 4496 33008 4505
rect 6644 4428 6696 4437
rect 7288 4471 7340 4480
rect 7288 4437 7297 4471
rect 7297 4437 7331 4471
rect 7331 4437 7340 4471
rect 7288 4428 7340 4437
rect 8944 4471 8996 4480
rect 8944 4437 8953 4471
rect 8953 4437 8987 4471
rect 8987 4437 8996 4471
rect 8944 4428 8996 4437
rect 10508 4471 10560 4480
rect 10508 4437 10517 4471
rect 10517 4437 10551 4471
rect 10551 4437 10560 4471
rect 10508 4428 10560 4437
rect 20260 4471 20312 4480
rect 20260 4437 20269 4471
rect 20269 4437 20303 4471
rect 20303 4437 20312 4471
rect 20260 4428 20312 4437
rect 20812 4428 20864 4480
rect 21916 4471 21968 4480
rect 21916 4437 21925 4471
rect 21925 4437 21959 4471
rect 21959 4437 21968 4471
rect 21916 4428 21968 4437
rect 24308 4471 24360 4480
rect 24308 4437 24317 4471
rect 24317 4437 24351 4471
rect 24351 4437 24360 4471
rect 24308 4428 24360 4437
rect 24860 4471 24912 4480
rect 24860 4437 24869 4471
rect 24869 4437 24903 4471
rect 24903 4437 24912 4471
rect 24860 4428 24912 4437
rect 29184 4471 29236 4480
rect 29184 4437 29193 4471
rect 29193 4437 29227 4471
rect 29227 4437 29236 4471
rect 29184 4428 29236 4437
rect 31116 4471 31168 4480
rect 31116 4437 31125 4471
rect 31125 4437 31159 4471
rect 31159 4437 31168 4471
rect 31116 4428 31168 4437
rect 7648 4326 7700 4378
rect 7712 4326 7764 4378
rect 7776 4326 7828 4378
rect 7840 4326 7892 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 34315 4326 34367 4378
rect 34379 4326 34431 4378
rect 34443 4326 34495 4378
rect 34507 4326 34559 4378
rect 2872 4224 2924 4276
rect 3608 4224 3660 4276
rect 6644 4267 6696 4276
rect 6644 4233 6653 4267
rect 6653 4233 6687 4267
rect 6687 4233 6696 4267
rect 6644 4224 6696 4233
rect 7196 4267 7248 4276
rect 7196 4233 7205 4267
rect 7205 4233 7239 4267
rect 7239 4233 7248 4267
rect 7196 4224 7248 4233
rect 7472 4224 7524 4276
rect 15844 4267 15896 4276
rect 15844 4233 15853 4267
rect 15853 4233 15887 4267
rect 15887 4233 15896 4267
rect 15844 4224 15896 4233
rect 16304 4267 16356 4276
rect 16304 4233 16313 4267
rect 16313 4233 16347 4267
rect 16347 4233 16356 4267
rect 16304 4224 16356 4233
rect 20076 4224 20128 4276
rect 21456 4224 21508 4276
rect 25780 4224 25832 4276
rect 26792 4267 26844 4276
rect 26792 4233 26801 4267
rect 26801 4233 26835 4267
rect 26835 4233 26844 4267
rect 26792 4224 26844 4233
rect 29184 4224 29236 4276
rect 29920 4267 29972 4276
rect 29920 4233 29929 4267
rect 29929 4233 29963 4267
rect 29963 4233 29972 4267
rect 29920 4224 29972 4233
rect 31116 4224 31168 4276
rect 33140 4224 33192 4276
rect 33416 4224 33468 4276
rect 2412 4088 2464 4140
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 3056 4131 3108 4140
rect 3056 4097 3065 4131
rect 3065 4097 3099 4131
rect 3099 4097 3108 4131
rect 3056 4088 3108 4097
rect 4620 4088 4672 4140
rect 6000 4131 6052 4140
rect 6000 4097 6009 4131
rect 6009 4097 6043 4131
rect 6043 4097 6052 4131
rect 6000 4088 6052 4097
rect 10508 4156 10560 4208
rect 19340 4199 19392 4208
rect 19340 4165 19349 4199
rect 19349 4165 19383 4199
rect 19383 4165 19392 4199
rect 19340 4156 19392 4165
rect 19800 4156 19852 4208
rect 22836 4199 22888 4208
rect 22836 4165 22845 4199
rect 22845 4165 22879 4199
rect 22879 4165 22888 4199
rect 22836 4156 22888 4165
rect 23204 4199 23256 4208
rect 23204 4165 23213 4199
rect 23213 4165 23247 4199
rect 23247 4165 23256 4199
rect 23204 4156 23256 4165
rect 25320 4156 25372 4208
rect 26700 4156 26752 4208
rect 16580 4131 16632 4140
rect 2780 4020 2832 4072
rect 6092 4020 6144 4072
rect 7288 4020 7340 4072
rect 2044 3952 2096 4004
rect 2872 3952 2924 4004
rect 3792 3952 3844 4004
rect 4528 3995 4580 4004
rect 4528 3961 4537 3995
rect 4537 3961 4571 3995
rect 4571 3961 4580 3995
rect 4528 3952 4580 3961
rect 2780 3884 2832 3936
rect 3700 3884 3752 3936
rect 7380 3952 7432 4004
rect 16580 4097 16589 4131
rect 16589 4097 16623 4131
rect 16623 4097 16632 4131
rect 16580 4088 16632 4097
rect 20260 4088 20312 4140
rect 25136 4131 25188 4140
rect 9496 4063 9548 4072
rect 9496 4029 9505 4063
rect 9505 4029 9539 4063
rect 9539 4029 9548 4063
rect 9496 4020 9548 4029
rect 25136 4097 25145 4131
rect 25145 4097 25179 4131
rect 25179 4097 25188 4131
rect 25136 4088 25188 4097
rect 27528 4088 27580 4140
rect 30472 4156 30524 4208
rect 30564 4088 30616 4140
rect 33232 4156 33284 4208
rect 21088 4063 21140 4072
rect 21088 4029 21122 4063
rect 21122 4029 21140 4063
rect 9220 3995 9272 4004
rect 9220 3961 9229 3995
rect 9229 3961 9263 3995
rect 9263 3961 9272 3995
rect 9220 3952 9272 3961
rect 9404 3995 9456 4004
rect 9404 3961 9413 3995
rect 9413 3961 9447 3995
rect 9447 3961 9456 3995
rect 9404 3952 9456 3961
rect 21088 4020 21140 4029
rect 24032 4063 24084 4072
rect 24032 4029 24041 4063
rect 24041 4029 24075 4063
rect 24075 4029 24084 4063
rect 24032 4020 24084 4029
rect 22008 3952 22060 4004
rect 24860 4020 24912 4072
rect 30748 4020 30800 4072
rect 24308 3995 24360 4004
rect 24308 3961 24317 3995
rect 24317 3961 24351 3995
rect 24351 3961 24360 3995
rect 24308 3952 24360 3961
rect 25044 3952 25096 4004
rect 27344 3952 27396 4004
rect 30196 3995 30248 4004
rect 30196 3961 30205 3995
rect 30205 3961 30239 3995
rect 30239 3961 30248 3995
rect 30196 3952 30248 3961
rect 4712 3884 4764 3936
rect 8668 3927 8720 3936
rect 8668 3893 8677 3927
rect 8677 3893 8711 3927
rect 8711 3893 8720 3927
rect 8668 3884 8720 3893
rect 21916 3884 21968 3936
rect 29644 3927 29696 3936
rect 29644 3893 29653 3927
rect 29653 3893 29687 3927
rect 29687 3893 29696 3927
rect 29644 3884 29696 3893
rect 30564 3884 30616 3936
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 27648 3782 27700 3834
rect 27712 3782 27764 3834
rect 27776 3782 27828 3834
rect 27840 3782 27892 3834
rect 2504 3680 2556 3732
rect 3056 3680 3108 3732
rect 3608 3723 3660 3732
rect 3608 3689 3617 3723
rect 3617 3689 3651 3723
rect 3651 3689 3660 3723
rect 3608 3680 3660 3689
rect 7104 3680 7156 3732
rect 7288 3680 7340 3732
rect 9404 3680 9456 3732
rect 20352 3723 20404 3732
rect 20352 3689 20361 3723
rect 20361 3689 20395 3723
rect 20395 3689 20404 3723
rect 20352 3680 20404 3689
rect 20720 3723 20772 3732
rect 20720 3689 20729 3723
rect 20729 3689 20763 3723
rect 20763 3689 20772 3723
rect 20720 3680 20772 3689
rect 21088 3723 21140 3732
rect 21088 3689 21097 3723
rect 21097 3689 21131 3723
rect 21131 3689 21140 3723
rect 21088 3680 21140 3689
rect 24032 3680 24084 3732
rect 24584 3680 24636 3732
rect 24860 3680 24912 3732
rect 27528 3680 27580 3732
rect 29000 3680 29052 3732
rect 30196 3680 30248 3732
rect 30380 3680 30432 3732
rect 1952 3612 2004 3664
rect 2412 3655 2464 3664
rect 2412 3621 2421 3655
rect 2421 3621 2455 3655
rect 2455 3621 2464 3655
rect 2412 3612 2464 3621
rect 9496 3612 9548 3664
rect 24768 3655 24820 3664
rect 24768 3621 24777 3655
rect 24777 3621 24811 3655
rect 24811 3621 24820 3655
rect 24768 3612 24820 3621
rect 25780 3612 25832 3664
rect 30748 3612 30800 3664
rect 2964 3544 3016 3596
rect 21916 3587 21968 3596
rect 21916 3553 21950 3587
rect 21950 3553 21968 3587
rect 21916 3544 21968 3553
rect 2320 3519 2372 3528
rect 2320 3485 2329 3519
rect 2329 3485 2363 3519
rect 2363 3485 2372 3519
rect 2320 3476 2372 3485
rect 2412 3476 2464 3528
rect 24676 3519 24728 3528
rect 1860 3408 1912 3460
rect 2872 3408 2924 3460
rect 9588 3408 9640 3460
rect 24676 3485 24685 3519
rect 24685 3485 24719 3519
rect 24719 3485 24728 3519
rect 24676 3476 24728 3485
rect 24216 3451 24268 3460
rect 24216 3417 24225 3451
rect 24225 3417 24259 3451
rect 24259 3417 24268 3451
rect 24216 3408 24268 3417
rect 3516 3340 3568 3392
rect 3884 3340 3936 3392
rect 4160 3340 4212 3392
rect 4712 3383 4764 3392
rect 4712 3349 4721 3383
rect 4721 3349 4755 3383
rect 4755 3349 4764 3383
rect 4712 3340 4764 3349
rect 21640 3340 21692 3392
rect 22008 3340 22060 3392
rect 23020 3383 23072 3392
rect 23020 3349 23029 3383
rect 23029 3349 23063 3383
rect 23063 3349 23072 3383
rect 23020 3340 23072 3349
rect 27344 3383 27396 3392
rect 27344 3349 27353 3383
rect 27353 3349 27387 3383
rect 27387 3349 27396 3383
rect 27344 3340 27396 3349
rect 7648 3238 7700 3290
rect 7712 3238 7764 3290
rect 7776 3238 7828 3290
rect 7840 3238 7892 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 34315 3238 34367 3290
rect 34379 3238 34431 3290
rect 34443 3238 34495 3290
rect 34507 3238 34559 3290
rect 2504 3136 2556 3188
rect 2964 3179 3016 3188
rect 2964 3145 2973 3179
rect 2973 3145 3007 3179
rect 3007 3145 3016 3179
rect 2964 3136 3016 3145
rect 1768 3000 1820 3052
rect 2412 3000 2464 3052
rect 2964 3000 3016 3052
rect 6552 3136 6604 3188
rect 21640 3179 21692 3188
rect 21640 3145 21649 3179
rect 21649 3145 21683 3179
rect 21683 3145 21692 3179
rect 21640 3136 21692 3145
rect 21916 3136 21968 3188
rect 24676 3136 24728 3188
rect 24768 3136 24820 3188
rect 20536 3111 20588 3120
rect 20536 3077 20545 3111
rect 20545 3077 20579 3111
rect 20579 3077 20588 3111
rect 20536 3068 20588 3077
rect 5264 3043 5316 3052
rect 5264 3009 5273 3043
rect 5273 3009 5307 3043
rect 5307 3009 5316 3043
rect 5264 3000 5316 3009
rect 23020 3000 23072 3052
rect 24584 3000 24636 3052
rect 20812 2975 20864 2984
rect 20812 2941 20821 2975
rect 20821 2941 20855 2975
rect 20855 2941 20864 2975
rect 20812 2932 20864 2941
rect 3516 2907 3568 2916
rect 3516 2873 3525 2907
rect 3525 2873 3559 2907
rect 3559 2873 3568 2907
rect 3516 2864 3568 2873
rect 4620 2864 4672 2916
rect 4988 2864 5040 2916
rect 20628 2864 20680 2916
rect 21364 2864 21416 2916
rect 2688 2839 2740 2848
rect 2688 2805 2697 2839
rect 2697 2805 2731 2839
rect 2731 2805 2740 2839
rect 2688 2796 2740 2805
rect 6828 2796 6880 2848
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 27648 2694 27700 2746
rect 27712 2694 27764 2746
rect 27776 2694 27828 2746
rect 27840 2694 27892 2746
rect 1952 2635 2004 2644
rect 1952 2601 1961 2635
rect 1961 2601 1995 2635
rect 1995 2601 2004 2635
rect 1952 2592 2004 2601
rect 2320 2635 2372 2644
rect 2320 2601 2329 2635
rect 2329 2601 2363 2635
rect 2363 2601 2372 2635
rect 2320 2592 2372 2601
rect 2964 2635 3016 2644
rect 2964 2601 2973 2635
rect 2973 2601 3007 2635
rect 3007 2601 3016 2635
rect 2964 2592 3016 2601
rect 4712 2592 4764 2644
rect 20628 2592 20680 2644
rect 4344 2499 4396 2508
rect 4344 2465 4378 2499
rect 4378 2465 4396 2499
rect 4344 2456 4396 2465
rect 4068 2431 4120 2440
rect 4068 2397 4077 2431
rect 4077 2397 4111 2431
rect 4111 2397 4120 2431
rect 4068 2388 4120 2397
rect 7648 2150 7700 2202
rect 7712 2150 7764 2202
rect 7776 2150 7828 2202
rect 7840 2150 7892 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 34315 2150 34367 2202
rect 34379 2150 34431 2202
rect 34443 2150 34495 2202
rect 34507 2150 34559 2202
<< metal2 >>
rect 1214 15520 1270 16000
rect 3054 15872 3110 15881
rect 3054 15807 3110 15816
rect 1228 12850 1256 15520
rect 3068 13870 3096 15807
rect 3698 15520 3754 16000
rect 6182 15520 6238 16000
rect 8666 15520 8722 16000
rect 11150 15520 11206 16000
rect 13634 15520 13690 16000
rect 16210 15520 16266 16000
rect 18694 15520 18750 16000
rect 21178 15520 21234 16000
rect 23662 15520 23718 16000
rect 26146 15520 26202 16000
rect 28722 15520 28778 16000
rect 31206 15520 31262 16000
rect 33690 15520 33746 16000
rect 36174 15520 36230 16000
rect 36726 15872 36782 15881
rect 36726 15807 36782 15816
rect 3422 15464 3478 15473
rect 3422 15399 3478 15408
rect 3330 15056 3386 15065
rect 3330 14991 3386 15000
rect 3344 13938 3372 14991
rect 3436 14074 3464 15399
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2136 13456 2188 13462
rect 2792 13433 2820 13466
rect 2136 13398 2188 13404
rect 2778 13424 2834 13433
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1216 12844 1268 12850
rect 1216 12786 1268 12792
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1400 12640 1452 12646
rect 1400 12582 1452 12588
rect 1412 10674 1440 12582
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1398 10160 1454 10169
rect 1398 10095 1454 10104
rect 1308 8832 1360 8838
rect 1308 8774 1360 8780
rect 1320 513 1348 8774
rect 1412 6458 1440 10095
rect 1504 8906 1532 12718
rect 1584 11824 1636 11830
rect 1582 11792 1584 11801
rect 1636 11792 1638 11801
rect 1582 11727 1638 11736
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1596 11150 1624 11630
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1688 9738 1716 13126
rect 1858 11112 1914 11121
rect 1858 11047 1914 11056
rect 1596 9710 1716 9738
rect 1596 9518 1624 9710
rect 1674 9616 1730 9625
rect 1872 9586 1900 11047
rect 2056 9994 2084 13262
rect 2148 11082 2176 13398
rect 2778 13359 2834 13368
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2332 12170 2360 13262
rect 2412 12912 2464 12918
rect 2412 12854 2464 12860
rect 2320 12164 2372 12170
rect 2320 12106 2372 12112
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2240 11354 2268 12038
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2332 11257 2360 12106
rect 2318 11248 2374 11257
rect 2318 11183 2374 11192
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 2044 9988 2096 9994
rect 2044 9930 2096 9936
rect 2332 9874 2360 11086
rect 2424 10062 2452 12854
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2504 12368 2556 12374
rect 2504 12310 2556 12316
rect 2516 11218 2544 12310
rect 2884 12238 2912 12650
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3424 12300 3476 12306
rect 3424 12242 3476 12248
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 3436 11665 3464 12242
rect 3528 12238 3556 12582
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3422 11656 3478 11665
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 3148 11620 3200 11626
rect 3422 11591 3478 11600
rect 3148 11562 3200 11568
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2516 10810 2544 11154
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2502 10296 2558 10305
rect 2502 10231 2504 10240
rect 2556 10231 2558 10240
rect 2504 10202 2556 10208
rect 2412 10056 2464 10062
rect 2410 10024 2412 10033
rect 2464 10024 2466 10033
rect 2410 9959 2466 9968
rect 2332 9846 2544 9874
rect 1674 9551 1730 9560
rect 1860 9580 1912 9586
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1492 8900 1544 8906
rect 1492 8842 1544 8848
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 1596 8265 1624 8502
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 6866 1532 7142
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1688 5370 1716 9551
rect 1860 9522 1912 9528
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1872 7750 1900 8230
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1872 7342 1900 7686
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1964 7154 1992 8910
rect 2424 7954 2452 8910
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 1872 7126 1992 7154
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1780 6186 1808 6802
rect 1768 6180 1820 6186
rect 1768 6122 1820 6128
rect 1780 5574 1808 6122
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 1688 4826 1716 5102
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1780 3058 1808 5510
rect 1872 3466 1900 7126
rect 2042 6624 2098 6633
rect 2042 6559 2098 6568
rect 2056 4010 2084 6559
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 2148 5574 2176 5646
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2148 4826 2176 5510
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 2148 4486 2176 4762
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 2240 4185 2268 5306
rect 2226 4176 2282 4185
rect 2226 4111 2282 4120
rect 2044 4004 2096 4010
rect 2044 3946 2096 3952
rect 1952 3664 2004 3670
rect 1952 3606 2004 3612
rect 1860 3460 1912 3466
rect 1860 3402 1912 3408
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1964 2650 1992 3606
rect 2332 3534 2360 7686
rect 2424 7342 2452 7890
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2424 7002 2452 7278
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2424 5370 2452 5714
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2410 4992 2466 5001
rect 2410 4927 2466 4936
rect 2424 4554 2452 4927
rect 2516 4729 2544 9846
rect 2608 7585 2636 11562
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2700 10198 2728 11086
rect 3160 11014 3188 11562
rect 3436 11558 3464 11591
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10538 3188 10950
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 3148 10532 3200 10538
rect 3148 10474 3200 10480
rect 2688 10192 2740 10198
rect 2688 10134 2740 10140
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2700 9382 2728 9522
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2700 8974 2728 9318
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2700 8430 2728 8910
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2792 8090 2820 9454
rect 2976 8838 3004 10474
rect 3160 9926 3188 10474
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3160 8906 3188 9862
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2976 8265 3004 8774
rect 3160 8362 3188 8842
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 2962 8256 3018 8265
rect 2962 8191 3018 8200
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 2594 7576 2650 7585
rect 2594 7511 2650 7520
rect 2608 6458 2636 7511
rect 2976 7274 3004 7958
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 3068 7002 3096 7822
rect 3160 7546 3188 8298
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3252 7177 3280 10406
rect 3238 7168 3294 7177
rect 3238 7103 3294 7112
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 3068 6186 3096 6938
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2700 4808 2728 5510
rect 2884 5370 2912 5782
rect 3068 5710 3096 6122
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 3160 5166 3188 5510
rect 3148 5160 3200 5166
rect 3146 5128 3148 5137
rect 3200 5128 3202 5137
rect 3146 5063 3202 5072
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 2780 4820 2832 4826
rect 2700 4780 2780 4808
rect 2780 4762 2832 4768
rect 2964 4752 3016 4758
rect 2502 4720 2558 4729
rect 2964 4694 3016 4700
rect 2502 4655 2558 4664
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2412 4548 2464 4554
rect 2412 4490 2464 4496
rect 2884 4282 2912 4558
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2424 3670 2452 4082
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2792 3942 2820 4014
rect 2884 4010 2912 4082
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2412 3664 2464 3670
rect 2412 3606 2464 3612
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2332 2650 2360 3470
rect 2424 3058 2452 3470
rect 2516 3194 2544 3674
rect 2884 3466 2912 3946
rect 2976 3602 3004 4694
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 3068 4146 3096 4422
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 3068 3738 3096 4082
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2976 3194 3004 3538
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 1306 504 1362 513
rect 1306 439 1362 448
rect 2700 241 2728 2790
rect 2976 2650 3004 2994
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3160 1737 3188 4966
rect 3146 1728 3202 1737
rect 3146 1663 3202 1672
rect 3252 1329 3280 7103
rect 3344 6934 3372 11494
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 3436 6746 3464 11494
rect 3528 7041 3556 11698
rect 3620 10810 3648 12038
rect 3712 11121 3740 15520
rect 4434 14648 4490 14657
rect 4434 14583 4490 14592
rect 4066 14240 4122 14249
rect 4066 14175 4122 14184
rect 4080 14006 4108 14175
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 4342 13832 4398 13841
rect 4342 13767 4398 13776
rect 4356 13530 4384 13767
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4158 13016 4214 13025
rect 4158 12951 4214 12960
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4080 12617 4108 12786
rect 4066 12608 4122 12617
rect 4066 12543 4122 12552
rect 4172 12442 4200 12951
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 4250 12200 4306 12209
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 3804 11354 3832 11766
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3896 11150 3924 12174
rect 4250 12135 4252 12144
rect 4304 12135 4306 12144
rect 4252 12106 4304 12112
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4356 11150 4384 11222
rect 3884 11144 3936 11150
rect 3698 11112 3754 11121
rect 3884 11086 3936 11092
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 3698 11047 3754 11056
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3698 10432 3754 10441
rect 3514 7032 3570 7041
rect 3514 6967 3570 6976
rect 3344 6718 3464 6746
rect 3344 4570 3372 6718
rect 3514 5264 3570 5273
rect 3514 5199 3570 5208
rect 3424 5092 3476 5098
rect 3424 5034 3476 5040
rect 3436 4690 3464 5034
rect 3528 5030 3556 5199
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3620 4593 3648 10406
rect 3698 10367 3754 10376
rect 3712 5409 3740 10367
rect 3804 6905 3832 10610
rect 3896 9926 3924 11086
rect 3974 10976 4030 10985
rect 3974 10911 4030 10920
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3896 9518 3924 9862
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3896 8634 3924 9454
rect 3988 9178 4016 10911
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4066 10568 4122 10577
rect 4066 10503 4122 10512
rect 4080 9625 4108 10503
rect 4356 10266 4384 10610
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 4066 9616 4122 9625
rect 4066 9551 4122 9560
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 4250 8936 4306 8945
rect 4250 8871 4306 8880
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 4158 8528 4214 8537
rect 4158 8463 4214 8472
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 4080 7546 4108 7890
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3976 7268 4028 7274
rect 3976 7210 4028 7216
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3988 7154 4016 7210
rect 3790 6896 3846 6905
rect 3790 6831 3792 6840
rect 3844 6831 3846 6840
rect 3792 6802 3844 6808
rect 3804 6458 3832 6802
rect 3896 6662 3924 7142
rect 3988 7126 4108 7154
rect 3974 7032 4030 7041
rect 3974 6967 4030 6976
rect 3988 6934 4016 6967
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3896 6338 3924 6598
rect 3804 6310 3924 6338
rect 3804 6254 3832 6310
rect 3792 6248 3844 6254
rect 3988 6202 4016 6870
rect 3792 6190 3844 6196
rect 3698 5400 3754 5409
rect 3698 5335 3754 5344
rect 3804 4604 3832 6190
rect 3896 6174 4016 6202
rect 3896 5250 3924 6174
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5846 4016 6054
rect 3976 5840 4028 5846
rect 3976 5782 4028 5788
rect 4080 5778 4108 7126
rect 4172 6730 4200 8463
rect 4264 8090 4292 8871
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4080 5658 4108 5714
rect 4080 5630 4200 5658
rect 3896 5222 4108 5250
rect 3884 5092 3936 5098
rect 3884 5034 3936 5040
rect 3896 4826 3924 5034
rect 4080 4978 4108 5222
rect 4172 5166 4200 5630
rect 4356 5370 4384 8774
rect 4448 5914 4476 14583
rect 4620 13456 4672 13462
rect 4620 13398 4672 13404
rect 4632 12986 4660 13398
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5184 12986 5212 13330
rect 4620 12980 4672 12986
rect 5172 12980 5224 12986
rect 4620 12922 4672 12928
rect 5092 12940 5172 12968
rect 4526 11928 4582 11937
rect 4526 11863 4582 11872
rect 4540 11762 4568 11863
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4632 10305 4660 11766
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4724 11286 4752 11562
rect 4802 11520 4858 11529
rect 4802 11455 4858 11464
rect 4712 11280 4764 11286
rect 4712 11222 4764 11228
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4724 10470 4752 11086
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4618 10296 4674 10305
rect 4618 10231 4674 10240
rect 4528 10192 4580 10198
rect 4528 10134 4580 10140
rect 4540 9722 4568 10134
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4526 9208 4582 9217
rect 4632 9178 4660 10231
rect 4724 10169 4752 10406
rect 4710 10160 4766 10169
rect 4710 10095 4766 10104
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4724 9518 4752 9862
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4526 9143 4582 9152
rect 4620 9172 4672 9178
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4540 5710 4568 9143
rect 4620 9114 4672 9120
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4632 8673 4660 8978
rect 4724 8974 4752 9454
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4618 8664 4674 8673
rect 4618 8599 4620 8608
rect 4672 8599 4674 8608
rect 4620 8570 4672 8576
rect 4816 7449 4844 11455
rect 4894 11112 4950 11121
rect 4894 11047 4950 11056
rect 4908 7857 4936 11047
rect 4986 10024 5042 10033
rect 4986 9959 5042 9968
rect 5000 9178 5028 9959
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5092 8634 5120 12940
rect 5172 12922 5224 12928
rect 6196 12850 6224 15520
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5170 12336 5226 12345
rect 5170 12271 5172 12280
rect 5224 12271 5226 12280
rect 5172 12242 5224 12248
rect 5184 11898 5212 12242
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 8022 5212 8230
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5276 7886 5304 8502
rect 5264 7880 5316 7886
rect 4894 7848 4950 7857
rect 5264 7822 5316 7828
rect 5368 7818 5396 12718
rect 5644 11898 5672 12786
rect 6472 12442 6500 13942
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7024 12986 7052 13874
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7116 13258 7144 13806
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 7208 12442 7236 14010
rect 8024 13388 8076 13394
rect 8024 13330 8076 13336
rect 7622 13084 7918 13104
rect 7678 13082 7702 13084
rect 7758 13082 7782 13084
rect 7838 13082 7862 13084
rect 7700 13030 7702 13082
rect 7764 13030 7776 13082
rect 7838 13030 7840 13082
rect 7678 13028 7702 13030
rect 7758 13028 7782 13030
rect 7838 13028 7862 13030
rect 7622 13008 7918 13028
rect 8036 12918 8064 13330
rect 8024 12912 8076 12918
rect 8024 12854 8076 12860
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 6196 11642 6224 12242
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6274 11792 6330 11801
rect 6274 11727 6276 11736
rect 6328 11727 6330 11736
rect 6276 11698 6328 11704
rect 6840 11694 6868 12038
rect 6828 11688 6880 11694
rect 6196 11614 6316 11642
rect 6828 11630 6880 11636
rect 6288 11558 6316 11614
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 5722 11384 5778 11393
rect 5722 11319 5778 11328
rect 5736 10810 5764 11319
rect 5906 11248 5962 11257
rect 5906 11183 5962 11192
rect 6184 11212 6236 11218
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5448 10464 5500 10470
rect 5446 10432 5448 10441
rect 5500 10432 5502 10441
rect 5446 10367 5502 10376
rect 5540 9648 5592 9654
rect 5538 9616 5540 9625
rect 5592 9616 5594 9625
rect 5538 9551 5594 9560
rect 5828 9353 5856 11018
rect 5920 10266 5948 11183
rect 6184 11154 6236 11160
rect 6196 10674 6224 11154
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6196 10470 6224 10610
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6196 10305 6224 10406
rect 6182 10296 6238 10305
rect 5908 10260 5960 10266
rect 6182 10231 6238 10240
rect 5908 10202 5960 10208
rect 5920 9722 5948 10202
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 6000 9376 6052 9382
rect 5814 9344 5870 9353
rect 6000 9318 6052 9324
rect 5814 9279 5870 9288
rect 6012 8945 6040 9318
rect 6092 9104 6144 9110
rect 6090 9072 6092 9081
rect 6144 9072 6146 9081
rect 6146 9030 6224 9058
rect 6090 9007 6146 9016
rect 6092 8968 6144 8974
rect 5998 8936 6054 8945
rect 5724 8900 5776 8906
rect 6092 8910 6144 8916
rect 5998 8871 6054 8880
rect 5724 8842 5776 8848
rect 5736 8498 5764 8842
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5722 8392 5778 8401
rect 5448 8356 5500 8362
rect 5722 8327 5724 8336
rect 5448 8298 5500 8304
rect 5776 8327 5778 8336
rect 5724 8298 5776 8304
rect 5460 8090 5488 8298
rect 6104 8090 6132 8910
rect 6196 8634 6224 9030
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 5908 7880 5960 7886
rect 6184 7880 6236 7886
rect 5908 7822 5960 7828
rect 6182 7848 6184 7857
rect 6236 7848 6238 7857
rect 4894 7783 4950 7792
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 4802 7440 4858 7449
rect 4802 7375 4858 7384
rect 5920 7313 5948 7822
rect 6182 7783 6238 7792
rect 6196 7546 6224 7783
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 5906 7304 5962 7313
rect 4712 7268 4764 7274
rect 5906 7239 5962 7248
rect 4712 7210 4764 7216
rect 4724 6798 4752 7210
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 5092 6458 5120 6802
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5460 6322 5488 6598
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 4988 5840 5040 5846
rect 4988 5782 5040 5788
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4908 5030 4936 5510
rect 5000 5234 5028 5782
rect 5644 5778 5672 7142
rect 6288 6934 6316 11494
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6380 8537 6408 10406
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6472 8906 6500 9862
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6460 8900 6512 8906
rect 6460 8842 6512 8848
rect 6564 8634 6592 8910
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6366 8528 6422 8537
rect 6366 8463 6422 8472
rect 6380 8362 6408 8463
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6276 6928 6328 6934
rect 6276 6870 6328 6876
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5736 6186 5764 6666
rect 5828 6361 5856 6734
rect 5814 6352 5870 6361
rect 5814 6287 5870 6296
rect 5828 6254 5856 6287
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5644 5370 5672 5714
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4896 5024 4948 5030
rect 4894 4992 4896 5001
rect 5092 5001 5120 5102
rect 4948 4992 4950 5001
rect 4080 4950 4200 4978
rect 4066 4856 4122 4865
rect 3884 4820 3936 4826
rect 4066 4791 4122 4800
rect 3884 4762 3936 4768
rect 3884 4616 3936 4622
rect 3606 4584 3662 4593
rect 3344 4542 3556 4570
rect 3528 4434 3556 4542
rect 3804 4576 3884 4604
rect 3884 4558 3936 4564
rect 3606 4519 3662 4528
rect 3528 4406 3740 4434
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3620 3738 3648 4218
rect 3712 3942 3740 4406
rect 3792 4004 3844 4010
rect 3792 3946 3844 3952
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3528 2922 3556 3334
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3238 1320 3294 1329
rect 3238 1255 3294 1264
rect 3804 921 3832 3946
rect 3896 3398 3924 4558
rect 4080 4185 4108 4791
rect 4066 4176 4122 4185
rect 4066 4111 4122 4120
rect 3974 3904 4030 3913
rect 3974 3839 4030 3848
rect 3884 3392 3936 3398
rect 3988 3369 4016 3839
rect 4172 3482 4200 4950
rect 4894 4927 4950 4936
rect 5078 4992 5134 5001
rect 5078 4927 5134 4936
rect 5736 4826 5764 6122
rect 5920 5914 5948 6734
rect 6288 6497 6316 6870
rect 6274 6488 6330 6497
rect 6274 6423 6276 6432
rect 6328 6423 6330 6432
rect 6276 6394 6328 6400
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 6012 5710 6040 6326
rect 6090 5944 6146 5953
rect 6090 5879 6092 5888
rect 6144 5879 6146 5888
rect 6092 5850 6144 5856
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4526 4040 4582 4049
rect 4526 3975 4528 3984
rect 4580 3975 4582 3984
rect 4528 3946 4580 3952
rect 4632 3777 4660 4082
rect 4724 3942 4752 4626
rect 6012 4146 6040 5646
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 6104 4078 6132 5850
rect 6564 5370 6592 8570
rect 6748 8430 6776 8978
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6748 8022 6776 8366
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6748 7002 6776 7278
rect 6736 6996 6788 7002
rect 6736 6938 6788 6944
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6656 6225 6684 6394
rect 6748 6254 6776 6938
rect 6736 6248 6788 6254
rect 6642 6216 6698 6225
rect 6736 6190 6788 6196
rect 6642 6151 6698 6160
rect 6748 5710 6776 6190
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4618 3768 4674 3777
rect 4618 3703 4674 3712
rect 4080 3454 4200 3482
rect 3884 3334 3936 3340
rect 3974 3360 4030 3369
rect 3974 3295 4030 3304
rect 4080 3210 4108 3454
rect 4724 3398 4752 3878
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 3896 3182 4108 3210
rect 3896 2145 3924 3182
rect 4068 2440 4120 2446
rect 4172 2428 4200 3334
rect 4620 2916 4672 2922
rect 4724 2904 4752 3334
rect 6564 3194 6592 5306
rect 6748 5302 6776 5646
rect 6840 5642 6868 11630
rect 7392 11558 7420 12242
rect 7622 11996 7918 12016
rect 7678 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7700 11942 7702 11994
rect 7764 11942 7776 11994
rect 7838 11942 7840 11994
rect 7678 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7622 11920 7918 11940
rect 8680 11762 8708 15520
rect 11164 12850 11192 15520
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 9586 12200 9642 12209
rect 9586 12135 9642 12144
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 9140 11694 9168 11725
rect 9128 11688 9180 11694
rect 9126 11656 9128 11665
rect 9180 11656 9182 11665
rect 9126 11591 9182 11600
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 8024 11552 8076 11558
rect 8944 11552 8996 11558
rect 8024 11494 8076 11500
rect 8942 11520 8944 11529
rect 8996 11520 8998 11529
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6932 7954 6960 10678
rect 7208 10538 7236 10950
rect 7622 10908 7918 10928
rect 7678 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7700 10854 7702 10906
rect 7764 10854 7776 10906
rect 7838 10854 7840 10906
rect 7678 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7622 10832 7918 10852
rect 8036 10713 8064 11494
rect 8942 11455 8998 11464
rect 9140 11354 9168 11591
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9232 11286 9260 11766
rect 9508 11762 9536 12038
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 8114 10840 8170 10849
rect 9232 10810 9260 11222
rect 8114 10775 8170 10784
rect 9220 10804 9272 10810
rect 8022 10704 8078 10713
rect 8022 10639 8078 10648
rect 8128 10577 8156 10775
rect 9220 10746 9272 10752
rect 8114 10568 8170 10577
rect 7196 10532 7248 10538
rect 9508 10538 9536 11698
rect 9600 11626 9628 12135
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9770 11112 9826 11121
rect 8114 10503 8170 10512
rect 9496 10532 9548 10538
rect 7196 10474 7248 10480
rect 9496 10474 9548 10480
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7024 9926 7052 10406
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 7024 8634 7052 9862
rect 7116 9586 7144 10066
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7102 8664 7158 8673
rect 7012 8628 7064 8634
rect 7102 8599 7158 8608
rect 7012 8570 7064 8576
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6656 4282 6684 4422
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 5262 3088 5318 3097
rect 5262 3023 5264 3032
rect 5316 3023 5318 3032
rect 5264 2994 5316 3000
rect 4672 2876 4752 2904
rect 4620 2858 4672 2864
rect 4724 2650 4752 2876
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4342 2544 4398 2553
rect 4342 2479 4344 2488
rect 4396 2479 4398 2488
rect 4344 2450 4396 2456
rect 4120 2400 4200 2428
rect 4068 2382 4120 2388
rect 3882 2136 3938 2145
rect 3882 2071 3938 2080
rect 3790 912 3846 921
rect 3790 847 3846 856
rect 5000 480 5028 2858
rect 6840 2854 6868 4966
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6932 2689 6960 7482
rect 7024 7478 7052 7958
rect 7012 7472 7064 7478
rect 7012 7414 7064 7420
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 7024 6458 7052 6870
rect 7116 6769 7144 8599
rect 7208 7818 7236 10474
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8298 10432 8354 10441
rect 7470 10024 7526 10033
rect 7470 9959 7526 9968
rect 7484 9110 7512 9959
rect 7622 9820 7918 9840
rect 7678 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7700 9766 7702 9818
rect 7764 9766 7776 9818
rect 7838 9766 7840 9818
rect 7678 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7622 9744 7918 9764
rect 8128 9450 8156 10406
rect 8298 10367 8354 10376
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8220 9518 8248 9862
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 7654 9344 7710 9353
rect 7654 9279 7710 9288
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 7300 8566 7328 9046
rect 7668 8974 7696 9279
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7102 6760 7158 6769
rect 7102 6695 7158 6704
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 7024 5778 7052 6122
rect 7116 5914 7144 6695
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 7300 5030 7328 8502
rect 7484 8294 7512 8774
rect 7622 8732 7918 8752
rect 7678 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7700 8678 7702 8730
rect 7764 8678 7776 8730
rect 7838 8678 7840 8730
rect 7678 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7622 8656 7918 8676
rect 8022 8664 8078 8673
rect 8128 8634 8156 9386
rect 8220 9178 8248 9454
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8022 8599 8078 8608
rect 8116 8628 8168 8634
rect 8036 8498 8064 8599
rect 8116 8570 8168 8576
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7576 7886 7604 8366
rect 7746 8120 7802 8129
rect 7746 8055 7802 8064
rect 7760 8022 7788 8055
rect 7748 8016 7800 8022
rect 7654 7984 7710 7993
rect 7748 7958 7800 7964
rect 7654 7919 7710 7928
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7668 7818 7696 7919
rect 7472 7812 7524 7818
rect 7472 7754 7524 7760
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7484 7546 7512 7754
rect 7622 7644 7918 7664
rect 7678 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7700 7590 7702 7642
rect 7764 7590 7776 7642
rect 7838 7590 7840 7642
rect 7678 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7622 7568 7918 7588
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7392 5386 7420 7414
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7576 6769 7604 6870
rect 7760 6798 7788 7210
rect 7748 6792 7800 6798
rect 7562 6760 7618 6769
rect 7748 6734 7800 6740
rect 7562 6695 7618 6704
rect 8036 6610 8064 8434
rect 8128 7342 8156 8570
rect 8220 8090 8248 9114
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8206 7576 8262 7585
rect 8206 7511 8262 7520
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8114 7032 8170 7041
rect 8220 7018 8248 7511
rect 8312 7041 8340 10367
rect 9508 10062 9536 10474
rect 9600 10248 9628 11086
rect 9770 11047 9772 11056
rect 9824 11047 9826 11056
rect 9772 11018 9824 11024
rect 9680 10260 9732 10266
rect 9600 10220 9680 10248
rect 9680 10202 9732 10208
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9048 9042 9076 9318
rect 9508 9178 9536 9998
rect 9876 9897 9904 11562
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10060 10606 10088 11154
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10336 10810 10364 11086
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10230 10704 10286 10713
rect 10230 10639 10286 10648
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9862 9888 9918 9897
rect 9862 9823 9918 9832
rect 9968 9722 9996 10066
rect 10060 9994 10088 10542
rect 10138 10296 10194 10305
rect 10244 10266 10272 10639
rect 10138 10231 10194 10240
rect 10232 10260 10284 10266
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 10152 8786 10180 10231
rect 10232 10202 10284 10208
rect 10244 9654 10272 10202
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10612 9217 10640 9318
rect 10598 9208 10654 9217
rect 10598 9143 10654 9152
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10230 8800 10286 8809
rect 9784 8401 9812 8774
rect 10152 8758 10230 8786
rect 10230 8735 10286 8744
rect 9956 8560 10008 8566
rect 9954 8528 9956 8537
rect 10008 8528 10010 8537
rect 9954 8463 10010 8472
rect 9770 8392 9826 8401
rect 9404 8356 9456 8362
rect 9770 8327 9826 8336
rect 9404 8298 9456 8304
rect 9416 8090 9444 8298
rect 10244 8090 10272 8735
rect 10428 8129 10456 8978
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10520 8362 10548 8910
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10414 8120 10470 8129
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 10232 8084 10284 8090
rect 10414 8055 10470 8064
rect 10232 8026 10284 8032
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 8942 7304 8998 7313
rect 8942 7239 8998 7248
rect 8170 6990 8248 7018
rect 8298 7032 8354 7041
rect 8114 6967 8170 6976
rect 8298 6967 8354 6976
rect 8956 6866 8984 7239
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 9600 6798 9628 7142
rect 9784 6934 9812 7686
rect 10244 7546 10272 8026
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10336 7206 10364 7686
rect 10324 7200 10376 7206
rect 10416 7200 10468 7206
rect 10324 7142 10376 7148
rect 10414 7168 10416 7177
rect 10468 7168 10470 7177
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9680 6656 9732 6662
rect 8036 6582 8248 6610
rect 9680 6598 9732 6604
rect 7622 6556 7918 6576
rect 7678 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7700 6502 7702 6554
rect 7764 6502 7776 6554
rect 7838 6502 7840 6554
rect 7678 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7622 6480 7918 6500
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 8036 5846 8064 6054
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 7622 5468 7918 5488
rect 7678 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7700 5414 7702 5466
rect 7764 5414 7776 5466
rect 7838 5414 7840 5466
rect 7678 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7622 5392 7918 5412
rect 7392 5358 7512 5386
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 7116 3777 7144 4694
rect 7208 4282 7236 4762
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7208 4049 7236 4218
rect 7300 4078 7328 4422
rect 7288 4072 7340 4078
rect 7194 4040 7250 4049
rect 7288 4014 7340 4020
rect 7194 3975 7250 3984
rect 7102 3768 7158 3777
rect 7300 3738 7328 4014
rect 7392 4010 7420 5238
rect 7484 4758 7512 5358
rect 8036 5352 8064 5782
rect 8128 5409 8156 6394
rect 7944 5324 8064 5352
rect 8114 5400 8170 5409
rect 8114 5335 8170 5344
rect 7944 5098 7972 5324
rect 7932 5092 7984 5098
rect 7932 5034 7984 5040
rect 7472 4752 7524 4758
rect 7472 4694 7524 4700
rect 7944 4622 7972 5034
rect 8220 4826 8248 6582
rect 9692 5953 9720 6598
rect 9784 6458 9812 6870
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9954 6760 10010 6769
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9876 6361 9904 6734
rect 9954 6695 10010 6704
rect 9862 6352 9918 6361
rect 9862 6287 9864 6296
rect 9916 6287 9918 6296
rect 9864 6258 9916 6264
rect 9876 6227 9904 6258
rect 9678 5944 9734 5953
rect 9678 5879 9734 5888
rect 9968 5817 9996 6695
rect 10152 6458 10180 6938
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10060 5914 10088 6258
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10140 5840 10192 5846
rect 9954 5808 10010 5817
rect 10336 5817 10364 7142
rect 10414 7103 10470 7112
rect 10520 6769 10548 8298
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10692 7472 10744 7478
rect 10692 7414 10744 7420
rect 10704 7002 10732 7414
rect 10796 7342 10824 7822
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10796 6866 10824 7278
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10506 6760 10562 6769
rect 10506 6695 10562 6704
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10796 5846 10824 6190
rect 10784 5840 10836 5846
rect 10140 5782 10192 5788
rect 10322 5808 10378 5817
rect 9954 5743 10010 5752
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9404 5296 9456 5302
rect 8758 5264 8814 5273
rect 9404 5238 9456 5244
rect 8758 5199 8814 5208
rect 8772 5030 8800 5199
rect 8942 5128 8998 5137
rect 8942 5063 8944 5072
rect 8996 5063 8998 5072
rect 8944 5034 8996 5040
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 7932 4616 7984 4622
rect 7470 4584 7526 4593
rect 7932 4558 7984 4564
rect 7470 4519 7526 4528
rect 7484 4282 7512 4519
rect 8956 4486 8984 5034
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 7622 4380 7918 4400
rect 7678 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7700 4326 7702 4378
rect 7764 4326 7776 4378
rect 7838 4326 7840 4378
rect 7678 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7622 4304 7918 4324
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 8956 4185 8984 4422
rect 8942 4176 8998 4185
rect 8942 4111 8998 4120
rect 9218 4040 9274 4049
rect 7380 4004 7432 4010
rect 9416 4010 9444 5238
rect 9508 4865 9536 5510
rect 9586 5128 9642 5137
rect 9586 5063 9588 5072
rect 9640 5063 9642 5072
rect 9588 5034 9640 5040
rect 9494 4856 9550 4865
rect 9494 4791 9550 4800
rect 9508 4078 9536 4791
rect 10152 4622 10180 5782
rect 10784 5782 10836 5788
rect 10322 5743 10378 5752
rect 10508 5772 10560 5778
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10244 4826 10272 5510
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10140 4616 10192 4622
rect 10138 4584 10140 4593
rect 10192 4584 10194 4593
rect 10138 4519 10194 4528
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9218 3975 9220 3984
rect 7380 3946 7432 3952
rect 9272 3975 9274 3984
rect 9404 4004 9456 4010
rect 9220 3946 9272 3952
rect 9404 3946 9456 3952
rect 8668 3936 8720 3942
rect 8666 3904 8668 3913
rect 8720 3904 8722 3913
rect 8666 3839 8722 3848
rect 9416 3738 9444 3946
rect 7102 3703 7104 3712
rect 7156 3703 7158 3712
rect 7288 3732 7340 3738
rect 7104 3674 7156 3680
rect 7288 3674 7340 3680
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 7116 3643 7144 3674
rect 9508 3670 9536 4014
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 9588 3460 9640 3466
rect 9640 3420 9720 3448
rect 9588 3402 9640 3408
rect 9692 3369 9720 3420
rect 9678 3360 9734 3369
rect 7622 3292 7918 3312
rect 9678 3295 9734 3304
rect 7678 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7700 3238 7702 3290
rect 7764 3238 7776 3290
rect 7838 3238 7840 3290
rect 7678 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7622 3216 7918 3236
rect 10336 2961 10364 5743
rect 10508 5714 10560 5720
rect 10520 4486 10548 5714
rect 10796 5302 10824 5782
rect 10888 5370 10916 12582
rect 12072 12368 12124 12374
rect 12072 12310 12124 12316
rect 12084 11898 12112 12310
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 12084 10577 12112 11834
rect 12360 11370 12388 12242
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12268 11354 12388 11370
rect 12268 11348 12400 11354
rect 12268 11342 12348 11348
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12176 10674 12204 11086
rect 12268 10985 12296 11342
rect 12348 11290 12400 11296
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12254 10976 12310 10985
rect 12254 10911 12310 10920
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 12070 10568 12126 10577
rect 11992 10526 12070 10554
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10980 9738 11008 9862
rect 10980 9710 11100 9738
rect 11072 9586 11100 9710
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11244 9512 11296 9518
rect 11150 9480 11206 9489
rect 11244 9454 11296 9460
rect 11150 9415 11152 9424
rect 11204 9415 11206 9424
rect 11152 9386 11204 9392
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10980 8945 11008 9046
rect 11256 8974 11284 9454
rect 11348 9178 11376 10202
rect 11992 10033 12020 10526
rect 12070 10503 12126 10512
rect 12176 10470 12204 10610
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12072 10056 12124 10062
rect 11978 10024 12034 10033
rect 12072 9998 12124 10004
rect 11978 9959 12034 9968
rect 11980 9648 12032 9654
rect 11426 9616 11482 9625
rect 12084 9636 12112 9998
rect 12032 9608 12112 9636
rect 11980 9590 12032 9596
rect 11426 9551 11428 9560
rect 11480 9551 11482 9560
rect 11428 9522 11480 9528
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11440 9110 11468 9318
rect 11428 9104 11480 9110
rect 11426 9072 11428 9081
rect 11704 9104 11756 9110
rect 11480 9072 11482 9081
rect 11704 9046 11756 9052
rect 11426 9007 11482 9016
rect 11440 8981 11468 9007
rect 11244 8968 11296 8974
rect 10966 8936 11022 8945
rect 11244 8910 11296 8916
rect 10966 8871 11022 8880
rect 10980 8634 11008 8871
rect 11256 8634 11284 8910
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11256 8430 11284 8570
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11532 7954 11560 8570
rect 11716 8566 11744 9046
rect 12084 8634 12112 9608
rect 12176 9518 12204 10406
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12268 9353 12296 10911
rect 12360 10810 12388 11154
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12360 10062 12388 10746
rect 12452 10266 12480 11766
rect 12544 10810 12572 12582
rect 13648 12374 13676 15520
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13740 12782 13768 13126
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 14924 12912 14976 12918
rect 14924 12854 14976 12860
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12728 11626 12756 12174
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12716 11620 12768 11626
rect 12716 11562 12768 11568
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12728 9450 12756 11562
rect 12806 11112 12862 11121
rect 12806 11047 12862 11056
rect 12820 10606 12848 11047
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12820 10130 12848 10542
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12254 9344 12310 9353
rect 12254 9279 12310 9288
rect 12728 8945 12756 9386
rect 12530 8936 12586 8945
rect 12530 8871 12586 8880
rect 12714 8936 12770 8945
rect 12714 8871 12770 8880
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11794 8256 11850 8265
rect 11794 8191 11850 8200
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11334 7848 11390 7857
rect 11334 7783 11336 7792
rect 11388 7783 11390 7792
rect 11336 7754 11388 7760
rect 11152 7744 11204 7750
rect 10966 7712 11022 7721
rect 11152 7686 11204 7692
rect 10966 7647 11022 7656
rect 10980 7274 11008 7647
rect 11164 7274 11192 7686
rect 11532 7478 11560 7890
rect 11520 7472 11572 7478
rect 11520 7414 11572 7420
rect 11808 7313 11836 8191
rect 12176 8022 12204 8774
rect 12544 8537 12572 8871
rect 12912 8673 12940 11698
rect 13004 11626 13032 12038
rect 13542 11656 13598 11665
rect 12992 11620 13044 11626
rect 13542 11591 13598 11600
rect 12992 11562 13044 11568
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13004 10266 13032 10406
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 13004 9994 13032 10202
rect 13096 10198 13124 10474
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 12992 9988 13044 9994
rect 12992 9930 13044 9936
rect 13464 9625 13492 11494
rect 13556 9994 13584 11591
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13648 10538 13676 10950
rect 13636 10532 13688 10538
rect 13636 10474 13688 10480
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 13450 9616 13506 9625
rect 13450 9551 13506 9560
rect 12990 9208 13046 9217
rect 12990 9143 13046 9152
rect 12898 8664 12954 8673
rect 12898 8599 12954 8608
rect 12530 8528 12586 8537
rect 12530 8463 12586 8472
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 12912 7750 12940 8230
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 11794 7304 11850 7313
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 11152 7268 11204 7274
rect 12912 7274 12940 7686
rect 11794 7239 11850 7248
rect 11980 7268 12032 7274
rect 11152 7210 11204 7216
rect 10966 6896 11022 6905
rect 11022 6866 11100 6882
rect 11022 6860 11112 6866
rect 11022 6854 11060 6860
rect 10966 6831 11022 6840
rect 11060 6802 11112 6808
rect 11164 6798 11192 7210
rect 11808 7002 11836 7239
rect 11980 7210 12032 7216
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10784 5296 10836 5302
rect 10784 5238 10836 5244
rect 11072 5166 11100 6326
rect 11348 6186 11376 6598
rect 11426 6352 11482 6361
rect 11532 6322 11560 6666
rect 11808 6458 11836 6938
rect 11992 6798 12020 7210
rect 12438 6896 12494 6905
rect 12164 6860 12216 6866
rect 13004 6866 13032 9143
rect 12438 6831 12494 6840
rect 12992 6860 13044 6866
rect 12164 6802 12216 6808
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11426 6287 11482 6296
rect 11520 6316 11572 6322
rect 11440 6254 11468 6287
rect 11520 6258 11572 6264
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 11348 5914 11376 6122
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11992 5778 12020 6734
rect 12176 6497 12204 6802
rect 12254 6760 12310 6769
rect 12254 6695 12310 6704
rect 12162 6488 12218 6497
rect 12162 6423 12164 6432
rect 12216 6423 12218 6432
rect 12164 6394 12216 6400
rect 12176 6363 12204 6394
rect 12268 5846 12296 6695
rect 12452 5914 12480 6831
rect 12992 6802 13044 6808
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12636 6322 12664 6598
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12440 5908 12492 5914
rect 12360 5868 12440 5896
rect 12256 5840 12308 5846
rect 12256 5782 12308 5788
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11426 5536 11482 5545
rect 11426 5471 11482 5480
rect 11440 5234 11468 5471
rect 12268 5370 12296 5782
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10888 4826 10916 4966
rect 11072 4826 11100 5102
rect 12360 4826 12388 5868
rect 12440 5850 12492 5856
rect 12544 5846 12572 6122
rect 13004 5914 13032 6802
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13372 5914 13400 6734
rect 13556 6458 13584 6734
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 13556 6186 13584 6394
rect 13544 6180 13596 6186
rect 13544 6122 13596 6128
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12544 5370 12572 5782
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12544 4865 12572 5306
rect 13372 5234 13400 5850
rect 13740 5642 13768 12718
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 14844 12306 14872 12854
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 13924 11898 13952 12242
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14289 10288 14585 10308
rect 13912 10192 13964 10198
rect 13912 10134 13964 10140
rect 14186 10160 14242 10169
rect 13820 9648 13872 9654
rect 13818 9616 13820 9625
rect 13872 9616 13874 9625
rect 13818 9551 13874 9560
rect 13924 9466 13952 10134
rect 14096 10124 14148 10130
rect 14186 10095 14242 10104
rect 14096 10066 14148 10072
rect 14002 9616 14058 9625
rect 14002 9551 14058 9560
rect 13832 9438 13952 9466
rect 13832 8838 13860 9438
rect 14016 9217 14044 9551
rect 14002 9208 14058 9217
rect 14108 9178 14136 10066
rect 14200 10062 14228 10095
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14200 9722 14228 9998
rect 14752 9722 14780 10542
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14740 9716 14792 9722
rect 14740 9658 14792 9664
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 14002 9143 14058 9152
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 13820 8832 13872 8838
rect 13818 8800 13820 8809
rect 13872 8800 13874 8809
rect 13818 8735 13874 8744
rect 14278 8800 14334 8809
rect 14278 8735 14334 8744
rect 13832 7546 13860 8735
rect 14292 8537 14320 8735
rect 14936 8634 14964 12854
rect 16224 12850 16252 15520
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 16960 12782 16988 13126
rect 17040 12912 17092 12918
rect 17040 12854 17092 12860
rect 16948 12776 17000 12782
rect 15028 12714 15424 12730
rect 16948 12718 17000 12724
rect 15028 12708 15436 12714
rect 15028 12702 15384 12708
rect 15028 12646 15056 12702
rect 15384 12650 15436 12656
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15028 9654 15056 12582
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 15120 11626 15148 12038
rect 15198 11792 15254 11801
rect 15198 11727 15254 11736
rect 15384 11756 15436 11762
rect 15108 11620 15160 11626
rect 15108 11562 15160 11568
rect 15120 10130 15148 11562
rect 15212 11558 15240 11727
rect 15384 11698 15436 11704
rect 15200 11552 15252 11558
rect 15396 11529 15424 11698
rect 15200 11494 15252 11500
rect 15382 11520 15438 11529
rect 15212 11082 15240 11494
rect 15382 11455 15438 11464
rect 15396 11257 15424 11455
rect 15382 11248 15438 11257
rect 15382 11183 15438 11192
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15212 9761 15240 11018
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15198 9752 15254 9761
rect 15304 9722 15332 9998
rect 15198 9687 15254 9696
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 15304 9518 15332 9658
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15120 8974 15148 9454
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 14278 8528 14334 8537
rect 14278 8463 14334 8472
rect 14462 8528 14518 8537
rect 15120 8498 15148 8910
rect 15396 8537 15424 10406
rect 15382 8528 15438 8537
rect 14462 8463 14464 8472
rect 14516 8463 14518 8472
rect 15108 8492 15160 8498
rect 14464 8434 14516 8440
rect 15382 8463 15438 8472
rect 15108 8434 15160 8440
rect 14188 8356 14240 8362
rect 14188 8298 14240 8304
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14200 7750 14228 8298
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 14660 7313 14688 8298
rect 15120 8294 15148 8434
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 15658 8392 15714 8401
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14646 7304 14702 7313
rect 14646 7239 14702 7248
rect 14289 7100 14585 7120
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14289 7024 14585 7044
rect 14660 6497 14688 7239
rect 14646 6488 14702 6497
rect 14646 6423 14702 6432
rect 14004 6384 14056 6390
rect 14002 6352 14004 6361
rect 14752 6361 14780 7686
rect 15120 6798 15148 8230
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 14056 6352 14058 6361
rect 14002 6287 14058 6296
rect 14738 6352 14794 6361
rect 14738 6287 14794 6296
rect 14002 6216 14058 6225
rect 14002 6151 14058 6160
rect 14016 5846 14044 6151
rect 14752 6089 14780 6287
rect 15120 6254 15148 6734
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 14738 6080 14794 6089
rect 14289 6012 14585 6032
rect 14738 6015 14794 6024
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 14188 5840 14240 5846
rect 14188 5782 14240 5788
rect 15108 5840 15160 5846
rect 15212 5828 15240 8366
rect 15658 8327 15660 8336
rect 15712 8327 15714 8336
rect 15660 8298 15712 8304
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15672 7721 15700 8026
rect 15658 7712 15714 7721
rect 15658 7647 15714 7656
rect 15474 7576 15530 7585
rect 15474 7511 15530 7520
rect 15488 7342 15516 7511
rect 15672 7478 15700 7647
rect 15660 7472 15712 7478
rect 15660 7414 15712 7420
rect 15476 7336 15528 7342
rect 15476 7278 15528 7284
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15396 6254 15424 6598
rect 15384 6248 15436 6254
rect 15384 6190 15436 6196
rect 15672 5914 15700 6734
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15160 5800 15240 5828
rect 15108 5782 15160 5788
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 13832 5522 13860 5714
rect 13740 5494 13860 5522
rect 13740 5370 13768 5494
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 14016 5302 14044 5782
rect 14200 5370 14228 5782
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14004 5296 14056 5302
rect 14004 5238 14056 5244
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 14289 4924 14585 4944
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 12530 4856 12586 4865
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 12348 4820 12400 4826
rect 14289 4848 14585 4868
rect 12530 4791 12586 4800
rect 12348 4762 12400 4768
rect 12544 4690 12572 4791
rect 15212 4690 15240 5800
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15764 4554 15792 12582
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15948 11354 15976 11698
rect 16040 11665 16068 12038
rect 16026 11656 16082 11665
rect 16026 11591 16082 11600
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 16132 11286 16160 12106
rect 16210 12064 16266 12073
rect 16210 11999 16266 12008
rect 16120 11280 16172 11286
rect 16120 11222 16172 11228
rect 16132 10266 16160 11222
rect 16224 11082 16252 11999
rect 16488 11824 16540 11830
rect 16488 11766 16540 11772
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 16212 11076 16264 11082
rect 16212 11018 16264 11024
rect 16316 10674 16344 11630
rect 16500 11150 16528 11766
rect 16960 11665 16988 12718
rect 17052 12374 17080 12854
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 16946 11656 17002 11665
rect 16946 11591 17002 11600
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16408 10810 16436 10950
rect 16500 10810 16528 11086
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16960 10130 16988 11591
rect 17052 11354 17080 12310
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17144 11626 17172 12174
rect 17880 11694 17908 13330
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17972 12073 18000 12242
rect 17958 12064 18014 12073
rect 17958 11999 18014 12008
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17132 11620 17184 11626
rect 17132 11562 17184 11568
rect 17500 11620 17552 11626
rect 17500 11562 17552 11568
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 17144 11286 17172 11562
rect 17132 11280 17184 11286
rect 17132 11222 17184 11228
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17328 10470 17356 11086
rect 17512 10674 17540 11562
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 17880 10810 17908 11222
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16408 9722 16436 9998
rect 17328 9722 17356 10406
rect 17880 10266 17908 10746
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17604 9722 17632 10066
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16684 8945 16712 9318
rect 16670 8936 16726 8945
rect 16670 8871 16726 8880
rect 16776 8634 16804 9454
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 17144 8537 17172 8978
rect 17130 8528 17186 8537
rect 17130 8463 17186 8472
rect 17144 8090 17172 8463
rect 17328 8294 17356 9658
rect 17604 9178 17632 9658
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 17316 8288 17368 8294
rect 17314 8256 17316 8265
rect 17368 8256 17370 8265
rect 17314 8191 17370 8200
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16304 7880 16356 7886
rect 16302 7848 16304 7857
rect 16356 7848 16358 7857
rect 16302 7783 16358 7792
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15856 5234 15884 7686
rect 16316 7546 16344 7783
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16212 7472 16264 7478
rect 16212 7414 16264 7420
rect 16578 7440 16634 7449
rect 16224 7041 16252 7414
rect 16776 7410 16804 7890
rect 17328 7886 17356 8191
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17038 7712 17094 7721
rect 17038 7647 17094 7656
rect 16578 7375 16580 7384
rect 16632 7375 16634 7384
rect 16764 7404 16816 7410
rect 16580 7346 16632 7352
rect 16764 7346 16816 7352
rect 16670 7304 16726 7313
rect 16670 7239 16672 7248
rect 16724 7239 16726 7248
rect 16672 7210 16724 7216
rect 16210 7032 16266 7041
rect 16776 7002 16804 7346
rect 16210 6967 16266 6976
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16500 6118 16528 6802
rect 16670 6488 16726 6497
rect 16670 6423 16726 6432
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16212 5568 16264 5574
rect 16212 5510 16264 5516
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 16224 5098 16252 5510
rect 16408 5302 16436 5646
rect 16500 5545 16528 6054
rect 16684 5914 16712 6423
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16776 5846 16804 6938
rect 17052 6769 17080 7647
rect 17224 7472 17276 7478
rect 17224 7414 17276 7420
rect 17038 6760 17094 6769
rect 17038 6695 17094 6704
rect 16854 6080 16910 6089
rect 16854 6015 16910 6024
rect 16764 5840 16816 5846
rect 16764 5782 16816 5788
rect 16580 5568 16632 5574
rect 16486 5536 16542 5545
rect 16580 5510 16632 5516
rect 16486 5471 16542 5480
rect 16396 5296 16448 5302
rect 16396 5238 16448 5244
rect 16212 5092 16264 5098
rect 16212 5034 16264 5040
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16132 4826 16160 4966
rect 16394 4856 16450 4865
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16316 4800 16394 4808
rect 16316 4780 16396 4800
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15752 4548 15804 4554
rect 15752 4490 15804 4496
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 10520 4214 10548 4422
rect 15856 4282 15884 4626
rect 16316 4282 16344 4780
rect 16448 4791 16450 4800
rect 16396 4762 16448 4768
rect 16592 4706 16620 5510
rect 16776 5370 16804 5782
rect 16868 5710 16896 6015
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16408 4678 16620 4706
rect 16408 4622 16436 4678
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 16304 4276 16356 4282
rect 16304 4218 16356 4224
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 16592 4146 16620 4678
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 10322 2952 10378 2961
rect 10322 2887 10378 2896
rect 14289 2748 14585 2768
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 6918 2680 6974 2689
rect 14289 2672 14585 2692
rect 6918 2615 6974 2624
rect 14922 2544 14978 2553
rect 14922 2479 14978 2488
rect 7622 2204 7918 2224
rect 7678 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7700 2150 7702 2202
rect 7764 2150 7776 2202
rect 7838 2150 7840 2202
rect 7678 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7622 2128 7918 2148
rect 14936 480 14964 2479
rect 17236 1465 17264 7414
rect 17328 7206 17356 7822
rect 17316 7200 17368 7206
rect 17316 7142 17368 7148
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17420 6866 17448 6938
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17420 6458 17448 6802
rect 17604 6662 17632 7890
rect 17592 6656 17644 6662
rect 17592 6598 17644 6604
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17328 5817 17356 5850
rect 17314 5808 17370 5817
rect 17314 5743 17370 5752
rect 17328 5234 17356 5743
rect 17406 5672 17462 5681
rect 17406 5607 17462 5616
rect 17420 5370 17448 5607
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17696 3641 17724 6054
rect 18064 5846 18092 8298
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18248 6798 18276 7142
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18248 6458 18276 6734
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18144 6384 18196 6390
rect 18144 6326 18196 6332
rect 18234 6352 18290 6361
rect 18156 6225 18184 6326
rect 18234 6287 18290 6296
rect 18142 6216 18198 6225
rect 18142 6151 18198 6160
rect 18248 5846 18276 6287
rect 18052 5840 18104 5846
rect 18052 5782 18104 5788
rect 18236 5840 18288 5846
rect 18236 5782 18288 5788
rect 17774 5400 17830 5409
rect 17774 5335 17776 5344
rect 17828 5335 17830 5344
rect 17776 5306 17828 5312
rect 17868 4820 17920 4826
rect 18064 4808 18092 5782
rect 18248 5681 18276 5782
rect 18234 5672 18290 5681
rect 18234 5607 18290 5616
rect 18144 5296 18196 5302
rect 18144 5238 18196 5244
rect 18156 4865 18184 5238
rect 17920 4780 18092 4808
rect 18142 4856 18198 4865
rect 18142 4791 18198 4800
rect 17868 4762 17920 4768
rect 18340 4049 18368 9318
rect 18432 6186 18460 12786
rect 18708 12374 18736 15520
rect 21192 13954 21220 15520
rect 20732 13926 21220 13954
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19536 11898 19564 12242
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 18602 11792 18658 11801
rect 18602 11727 18658 11736
rect 18616 11626 18644 11727
rect 18694 11656 18750 11665
rect 18604 11620 18656 11626
rect 18694 11591 18696 11600
rect 18604 11562 18656 11568
rect 18748 11591 18750 11600
rect 18696 11562 18748 11568
rect 19982 11248 20038 11257
rect 19982 11183 20038 11192
rect 18696 11008 18748 11014
rect 18602 10976 18658 10985
rect 18696 10950 18748 10956
rect 18602 10911 18658 10920
rect 18616 9217 18644 10911
rect 18708 10810 18736 10950
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 19524 10464 19576 10470
rect 19062 10432 19118 10441
rect 19524 10406 19576 10412
rect 19062 10367 19118 10376
rect 18786 10024 18842 10033
rect 18786 9959 18842 9968
rect 18800 9654 18828 9959
rect 18788 9648 18840 9654
rect 18788 9590 18840 9596
rect 18880 9444 18932 9450
rect 18880 9386 18932 9392
rect 18602 9208 18658 9217
rect 18602 9143 18658 9152
rect 18616 8634 18644 9143
rect 18892 8838 18920 9386
rect 19076 8945 19104 10367
rect 19430 10296 19486 10305
rect 19430 10231 19486 10240
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 19352 9178 19380 10134
rect 19444 9382 19472 10231
rect 19536 9926 19564 10406
rect 19800 10056 19852 10062
rect 19800 9998 19852 10004
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19536 9586 19564 9862
rect 19812 9722 19840 9998
rect 19800 9716 19852 9722
rect 19800 9658 19852 9664
rect 19904 9586 19932 9998
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19062 8936 19118 8945
rect 19062 8871 19118 8880
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18616 8362 18644 8570
rect 18694 8392 18750 8401
rect 18604 8356 18656 8362
rect 18694 8327 18750 8336
rect 18604 8298 18656 8304
rect 18708 8090 18736 8327
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18602 7032 18658 7041
rect 18602 6967 18658 6976
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18420 6180 18472 6186
rect 18420 6122 18472 6128
rect 18524 6066 18552 6598
rect 18616 6186 18644 6967
rect 18892 6905 18920 8774
rect 19076 8634 19104 8871
rect 19352 8634 19380 9114
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19076 8430 19104 8570
rect 19444 8514 19472 8978
rect 19352 8486 19472 8514
rect 19536 8498 19564 9522
rect 19800 9104 19852 9110
rect 19800 9046 19852 9052
rect 19812 8809 19840 9046
rect 19996 9042 20024 11183
rect 20168 11008 20220 11014
rect 20168 10950 20220 10956
rect 20180 9897 20208 10950
rect 20456 10010 20484 12650
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20548 12442 20576 12582
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 20628 12368 20680 12374
rect 20732 12356 20760 13926
rect 23572 13728 23624 13734
rect 23572 13670 23624 13676
rect 22468 13388 22520 13394
rect 22468 13330 22520 13336
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 21548 12912 21600 12918
rect 21548 12854 21600 12860
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20680 12328 20760 12356
rect 20628 12310 20680 12316
rect 20824 10577 20852 12582
rect 21560 12306 21588 12854
rect 22376 12776 22428 12782
rect 22376 12718 22428 12724
rect 22192 12708 22244 12714
rect 22192 12650 22244 12656
rect 22204 12442 22232 12650
rect 22192 12436 22244 12442
rect 22192 12378 22244 12384
rect 21732 12368 21784 12374
rect 21732 12310 21784 12316
rect 21548 12300 21600 12306
rect 21548 12242 21600 12248
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 21284 11762 21312 12038
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 21456 11620 21508 11626
rect 21456 11562 21508 11568
rect 21468 11393 21496 11562
rect 21454 11384 21510 11393
rect 21560 11354 21588 12242
rect 21744 12102 21772 12310
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21732 12096 21784 12102
rect 21732 12038 21784 12044
rect 21744 11830 21772 12038
rect 21836 11898 21864 12174
rect 21824 11892 21876 11898
rect 21824 11834 21876 11840
rect 21732 11824 21784 11830
rect 21732 11766 21784 11772
rect 21836 11626 21864 11834
rect 21824 11620 21876 11626
rect 21824 11562 21876 11568
rect 22204 11558 22232 12378
rect 22388 11762 22416 12718
rect 22480 12646 22508 13330
rect 22664 12782 22692 13330
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22848 12986 22876 13262
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 23584 12850 23612 13670
rect 23676 12850 23704 15520
rect 25412 13864 25464 13870
rect 25412 13806 25464 13812
rect 24032 13524 24084 13530
rect 24032 13466 24084 13472
rect 24044 13297 24072 13466
rect 25424 13326 25452 13806
rect 26160 13530 26188 15520
rect 27622 13628 27918 13648
rect 27678 13626 27702 13628
rect 27758 13626 27782 13628
rect 27838 13626 27862 13628
rect 27700 13574 27702 13626
rect 27764 13574 27776 13626
rect 27838 13574 27840 13626
rect 27678 13572 27702 13574
rect 27758 13572 27782 13574
rect 27838 13572 27862 13574
rect 27622 13552 27918 13572
rect 26148 13524 26200 13530
rect 26148 13466 26200 13472
rect 28540 13524 28592 13530
rect 28540 13466 28592 13472
rect 25504 13456 25556 13462
rect 25504 13398 25556 13404
rect 26608 13456 26660 13462
rect 26608 13398 26660 13404
rect 25412 13320 25464 13326
rect 24030 13288 24086 13297
rect 25412 13262 25464 13268
rect 24030 13223 24086 13232
rect 24584 13252 24636 13258
rect 24584 13194 24636 13200
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 24030 13016 24086 13025
rect 24030 12951 24086 12960
rect 24044 12918 24072 12951
rect 24032 12912 24084 12918
rect 24032 12854 24084 12860
rect 23572 12844 23624 12850
rect 23572 12786 23624 12792
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22468 12640 22520 12646
rect 22468 12582 22520 12588
rect 23020 12640 23072 12646
rect 23020 12582 23072 12588
rect 22928 12300 22980 12306
rect 22928 12242 22980 12248
rect 22940 12209 22968 12242
rect 22926 12200 22982 12209
rect 22926 12135 22982 12144
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22940 11694 22968 12135
rect 22928 11688 22980 11694
rect 22926 11656 22928 11665
rect 22980 11656 22982 11665
rect 22376 11620 22428 11626
rect 22926 11591 22982 11600
rect 22376 11562 22428 11568
rect 21732 11552 21784 11558
rect 21732 11494 21784 11500
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 21454 11319 21510 11328
rect 21548 11348 21600 11354
rect 21548 11290 21600 11296
rect 21272 11144 21324 11150
rect 21272 11086 21324 11092
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 20810 10568 20866 10577
rect 20810 10503 20866 10512
rect 21284 10470 21312 11086
rect 21744 10810 21772 11494
rect 22204 11218 22232 11494
rect 22388 11286 22416 11562
rect 22376 11280 22428 11286
rect 22376 11222 22428 11228
rect 22928 11280 22980 11286
rect 22928 11222 22980 11228
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 22190 10840 22246 10849
rect 21732 10804 21784 10810
rect 22190 10775 22246 10784
rect 21732 10746 21784 10752
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 21180 10464 21232 10470
rect 20626 10432 20682 10441
rect 21180 10406 21232 10412
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 20626 10367 20682 10376
rect 20456 9982 20576 10010
rect 20640 9994 20668 10367
rect 21192 10130 21220 10406
rect 21284 10198 21312 10406
rect 21836 10254 22048 10282
rect 22112 10266 22140 10610
rect 22204 10577 22232 10775
rect 22388 10674 22416 11222
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 22468 11008 22520 11014
rect 22468 10950 22520 10956
rect 22376 10668 22428 10674
rect 22376 10610 22428 10616
rect 22480 10577 22508 10950
rect 22664 10674 22692 11154
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22190 10568 22246 10577
rect 22466 10568 22522 10577
rect 22190 10503 22246 10512
rect 22284 10532 22336 10538
rect 22466 10503 22522 10512
rect 22284 10474 22336 10480
rect 22296 10441 22324 10474
rect 22282 10432 22338 10441
rect 22282 10367 22338 10376
rect 22664 10266 22692 10610
rect 21272 10192 21324 10198
rect 21272 10134 21324 10140
rect 21180 10124 21232 10130
rect 21180 10066 21232 10072
rect 21284 10062 21312 10134
rect 21836 10130 21864 10254
rect 22020 10198 22048 10254
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22008 10192 22060 10198
rect 22008 10134 22060 10140
rect 22192 10192 22244 10198
rect 22192 10134 22244 10140
rect 21824 10124 21876 10130
rect 21824 10066 21876 10072
rect 21916 10124 21968 10130
rect 21916 10066 21968 10072
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 20444 9920 20496 9926
rect 20166 9888 20222 9897
rect 20444 9862 20496 9868
rect 20548 9874 20576 9982
rect 20628 9988 20680 9994
rect 20628 9930 20680 9936
rect 20824 9880 21312 9908
rect 20824 9874 20852 9880
rect 20166 9823 20222 9832
rect 20074 9616 20130 9625
rect 20074 9551 20076 9560
rect 20128 9551 20130 9560
rect 20076 9522 20128 9528
rect 20088 9382 20116 9522
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19798 8800 19854 8809
rect 19798 8735 19854 8744
rect 19524 8492 19576 8498
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 19352 7750 19380 8486
rect 19524 8434 19576 8440
rect 19812 8022 19840 8735
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19996 8090 20024 8434
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19800 8016 19852 8022
rect 19800 7958 19852 7964
rect 19340 7744 19392 7750
rect 19338 7712 19340 7721
rect 19392 7712 19394 7721
rect 19338 7647 19394 7656
rect 19430 7576 19486 7585
rect 19430 7511 19486 7520
rect 19444 7410 19472 7511
rect 19616 7472 19668 7478
rect 19614 7440 19616 7449
rect 19668 7440 19670 7449
rect 20180 7426 20208 9823
rect 20352 9648 20404 9654
rect 20352 9590 20404 9596
rect 20364 9178 20392 9590
rect 20456 9518 20484 9862
rect 20548 9846 20852 9874
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20456 9058 20484 9454
rect 20364 9030 20484 9058
rect 20364 8974 20392 9030
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 20364 8362 20392 8910
rect 20352 8356 20404 8362
rect 20352 8298 20404 8304
rect 19432 7404 19484 7410
rect 19614 7375 19670 7384
rect 20088 7398 20208 7426
rect 20640 7410 20668 9846
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 21284 9722 21312 9880
rect 21272 9716 21324 9722
rect 21272 9658 21324 9664
rect 20720 9444 20772 9450
rect 20720 9386 20772 9392
rect 20732 8838 20760 9386
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21732 9376 21784 9382
rect 21732 9318 21784 9324
rect 21284 9081 21312 9318
rect 21640 9104 21692 9110
rect 21270 9072 21326 9081
rect 21640 9046 21692 9052
rect 21270 9007 21326 9016
rect 20812 8900 20864 8906
rect 20812 8842 20864 8848
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20732 8090 20760 8774
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20824 7954 20852 8842
rect 21652 8838 21680 9046
rect 21640 8832 21692 8838
rect 21640 8774 21692 8780
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 20904 8424 20956 8430
rect 20904 8366 20956 8372
rect 21454 8392 21510 8401
rect 20916 8294 20944 8366
rect 21454 8327 21456 8336
rect 21508 8327 21510 8336
rect 21456 8298 21508 8304
rect 20904 8288 20956 8294
rect 20902 8256 20904 8265
rect 20956 8256 20958 8265
rect 20902 8191 20958 8200
rect 20812 7948 20864 7954
rect 20812 7890 20864 7896
rect 20916 7834 20944 8191
rect 21468 8090 21496 8298
rect 21652 8090 21680 8774
rect 21744 8537 21772 9318
rect 21928 8838 21956 10066
rect 22204 9586 22232 10134
rect 22664 9926 22692 10202
rect 22652 9920 22704 9926
rect 22652 9862 22704 9868
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 21730 8528 21786 8537
rect 21730 8463 21786 8472
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 21640 8084 21692 8090
rect 21640 8026 21692 8032
rect 21928 7886 21956 8774
rect 22020 8537 22048 9454
rect 22204 9178 22232 9522
rect 22376 9376 22428 9382
rect 22376 9318 22428 9324
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22388 9081 22416 9318
rect 22940 9217 22968 11222
rect 22926 9208 22982 9217
rect 22848 9166 22926 9194
rect 22374 9072 22430 9081
rect 22192 9036 22244 9042
rect 22374 9007 22430 9016
rect 22192 8978 22244 8984
rect 22006 8528 22062 8537
rect 22006 8463 22062 8472
rect 22204 8294 22232 8978
rect 22192 8288 22244 8294
rect 22192 8230 22244 8236
rect 22204 7954 22232 8230
rect 22192 7948 22244 7954
rect 22192 7890 22244 7896
rect 20824 7806 20944 7834
rect 21916 7880 21968 7886
rect 21916 7822 21968 7828
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 20824 7546 20852 7806
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 21638 7576 21694 7585
rect 20812 7540 20864 7546
rect 21638 7511 21694 7520
rect 20812 7482 20864 7488
rect 20628 7404 20680 7410
rect 19432 7346 19484 7352
rect 18878 6896 18934 6905
rect 18878 6831 18934 6840
rect 18604 6180 18656 6186
rect 18604 6122 18656 6128
rect 18696 6180 18748 6186
rect 18696 6122 18748 6128
rect 18708 6066 18736 6122
rect 18524 6038 18736 6066
rect 18708 5574 18736 6038
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18510 5264 18566 5273
rect 18510 5199 18512 5208
rect 18564 5199 18566 5208
rect 18512 5170 18564 5176
rect 18602 5128 18658 5137
rect 18708 5098 18736 5510
rect 18786 5128 18842 5137
rect 18602 5063 18604 5072
rect 18656 5063 18658 5072
rect 18696 5092 18748 5098
rect 18604 5034 18656 5040
rect 18786 5063 18842 5072
rect 18696 5034 18748 5040
rect 18616 4826 18644 5034
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 18616 4729 18644 4762
rect 18708 4758 18736 5034
rect 18696 4752 18748 4758
rect 18602 4720 18658 4729
rect 18696 4694 18748 4700
rect 18602 4655 18658 4664
rect 18800 4321 18828 5063
rect 18786 4312 18842 4321
rect 18786 4247 18842 4256
rect 18326 4040 18382 4049
rect 18326 3975 18382 3984
rect 17682 3632 17738 3641
rect 17682 3567 17738 3576
rect 18892 2961 18920 6831
rect 19800 5704 19852 5710
rect 19800 5646 19852 5652
rect 19522 5400 19578 5409
rect 19522 5335 19524 5344
rect 19576 5335 19578 5344
rect 19524 5306 19576 5312
rect 19536 5030 19564 5306
rect 19812 5166 19840 5646
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 20088 4826 20116 7398
rect 20628 7346 20680 7352
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 20168 7268 20220 7274
rect 20168 7210 20220 7216
rect 20180 6905 20208 7210
rect 20628 7200 20680 7206
rect 20680 7148 20760 7154
rect 20628 7142 20760 7148
rect 20640 7126 20760 7142
rect 20166 6896 20222 6905
rect 20166 6831 20222 6840
rect 20732 5642 20760 7126
rect 21100 6934 21128 7346
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 21192 7002 21220 7210
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 21088 6928 21140 6934
rect 21088 6870 21140 6876
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 20810 6080 20866 6089
rect 20810 6015 20866 6024
rect 20824 5710 20852 6015
rect 21652 5914 21680 7511
rect 22112 6934 22140 7822
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 22100 6928 22152 6934
rect 22100 6870 22152 6876
rect 22374 6896 22430 6905
rect 22112 6458 22140 6870
rect 22374 6831 22376 6840
rect 22428 6831 22430 6840
rect 22376 6802 22428 6808
rect 22388 6458 22416 6802
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 22376 6452 22428 6458
rect 22376 6394 22428 6400
rect 21732 6180 21784 6186
rect 21732 6122 21784 6128
rect 21640 5908 21692 5914
rect 21560 5868 21640 5896
rect 21560 5817 21588 5868
rect 21640 5850 21692 5856
rect 21744 5846 21772 6122
rect 22388 5914 22416 6394
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 22480 5846 22508 7142
rect 21732 5840 21784 5846
rect 21546 5808 21602 5817
rect 21456 5772 21508 5778
rect 22468 5840 22520 5846
rect 21732 5782 21784 5788
rect 21822 5808 21878 5817
rect 21546 5743 21602 5752
rect 22468 5782 22520 5788
rect 21822 5743 21824 5752
rect 21456 5714 21508 5720
rect 20812 5704 20864 5710
rect 20812 5646 20864 5652
rect 20720 5636 20772 5642
rect 20720 5578 20772 5584
rect 20824 5370 20852 5646
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20352 5296 20404 5302
rect 20352 5238 20404 5244
rect 21180 5296 21232 5302
rect 21180 5238 21232 5244
rect 21364 5296 21416 5302
rect 21364 5238 21416 5244
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20076 4820 20128 4826
rect 20076 4762 20128 4768
rect 19798 4720 19854 4729
rect 19798 4655 19854 4664
rect 19812 4622 19840 4655
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19812 4214 19840 4558
rect 20088 4282 20116 4762
rect 20272 4622 20300 5102
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20272 4486 20300 4558
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 20076 4276 20128 4282
rect 20076 4218 20128 4224
rect 19340 4208 19392 4214
rect 19340 4150 19392 4156
rect 19800 4208 19852 4214
rect 19800 4150 19852 4156
rect 19352 3369 19380 4150
rect 20272 4146 20300 4422
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20364 3738 20392 5238
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20456 3641 20484 4966
rect 21192 4690 21220 5238
rect 21180 4684 21232 4690
rect 21180 4626 21232 4632
rect 20720 4548 20772 4554
rect 20720 4490 20772 4496
rect 20732 3738 20760 4490
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20442 3632 20498 3641
rect 20442 3567 20498 3576
rect 19338 3360 19394 3369
rect 19338 3295 19394 3304
rect 20536 3120 20588 3126
rect 20534 3088 20536 3097
rect 20588 3088 20590 3097
rect 20534 3023 20590 3032
rect 20824 2990 20852 4422
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 21088 4072 21140 4078
rect 21086 4040 21088 4049
rect 21140 4040 21142 4049
rect 21086 3975 21142 3984
rect 21100 3738 21128 3975
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 20812 2984 20864 2990
rect 18878 2952 18934 2961
rect 20812 2926 20864 2932
rect 21376 2922 21404 5238
rect 21468 5166 21496 5714
rect 21560 5370 21588 5743
rect 21876 5743 21878 5752
rect 22008 5772 22060 5778
rect 21824 5714 21876 5720
rect 22008 5714 22060 5720
rect 21548 5364 21600 5370
rect 21548 5306 21600 5312
rect 21824 5296 21876 5302
rect 21824 5238 21876 5244
rect 21456 5160 21508 5166
rect 21456 5102 21508 5108
rect 21468 4282 21496 5102
rect 21836 5030 21864 5238
rect 21916 5092 21968 5098
rect 21916 5034 21968 5040
rect 21824 5024 21876 5030
rect 21824 4966 21876 4972
rect 21836 4826 21864 4966
rect 21824 4820 21876 4826
rect 21824 4762 21876 4768
rect 21928 4486 21956 5034
rect 21916 4480 21968 4486
rect 21916 4422 21968 4428
rect 21456 4276 21508 4282
rect 21456 4218 21508 4224
rect 21928 3942 21956 4422
rect 22020 4010 22048 5714
rect 22480 5370 22508 5782
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22848 4740 22876 9166
rect 22926 9143 22982 9152
rect 23032 8906 23060 12582
rect 23296 12368 23348 12374
rect 23294 12336 23296 12345
rect 23348 12336 23350 12345
rect 23294 12271 23350 12280
rect 23308 11898 23336 12271
rect 23848 12232 23900 12238
rect 23848 12174 23900 12180
rect 23296 11892 23348 11898
rect 23348 11852 23428 11880
rect 23296 11834 23348 11840
rect 23296 11008 23348 11014
rect 23296 10950 23348 10956
rect 23308 10606 23336 10950
rect 23296 10600 23348 10606
rect 23296 10542 23348 10548
rect 23202 8936 23258 8945
rect 23020 8900 23072 8906
rect 23202 8871 23258 8880
rect 23020 8842 23072 8848
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 22940 7750 22968 8230
rect 22928 7744 22980 7750
rect 22928 7686 22980 7692
rect 22940 7274 22968 7686
rect 22928 7268 22980 7274
rect 22928 7210 22980 7216
rect 23112 7200 23164 7206
rect 23112 7142 23164 7148
rect 23124 6934 23152 7142
rect 23112 6928 23164 6934
rect 23112 6870 23164 6876
rect 23124 6458 23152 6870
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23124 5846 23152 6394
rect 23112 5840 23164 5846
rect 23112 5782 23164 5788
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 22940 5250 22968 5714
rect 23124 5370 23152 5782
rect 23216 5370 23244 8871
rect 23400 8265 23428 11852
rect 23756 11144 23808 11150
rect 23756 11086 23808 11092
rect 23768 10606 23796 11086
rect 23860 11014 23888 12174
rect 24044 11694 24072 12854
rect 24320 12782 24348 13126
rect 24596 12918 24624 13194
rect 24860 13184 24912 13190
rect 24860 13126 24912 13132
rect 25044 13184 25096 13190
rect 25044 13126 25096 13132
rect 25228 13184 25280 13190
rect 25228 13126 25280 13132
rect 24584 12912 24636 12918
rect 24584 12854 24636 12860
rect 24872 12832 24900 13126
rect 24952 12844 25004 12850
rect 24872 12804 24952 12832
rect 24952 12786 25004 12792
rect 24308 12776 24360 12782
rect 24308 12718 24360 12724
rect 25056 12714 25084 13126
rect 25044 12708 25096 12714
rect 25044 12650 25096 12656
rect 24952 12368 25004 12374
rect 24952 12310 25004 12316
rect 24584 12164 24636 12170
rect 24584 12106 24636 12112
rect 24400 12096 24452 12102
rect 24398 12064 24400 12073
rect 24452 12064 24454 12073
rect 24398 11999 24454 12008
rect 24032 11688 24084 11694
rect 24032 11630 24084 11636
rect 24412 11626 24440 11999
rect 24596 11762 24624 12106
rect 24964 11937 24992 12310
rect 24950 11928 25006 11937
rect 24950 11863 25006 11872
rect 24584 11756 24636 11762
rect 24584 11698 24636 11704
rect 24400 11620 24452 11626
rect 24400 11562 24452 11568
rect 24964 11558 24992 11863
rect 24952 11552 25004 11558
rect 24674 11520 24730 11529
rect 24952 11494 25004 11500
rect 24674 11455 24730 11464
rect 24688 11218 24716 11455
rect 24124 11212 24176 11218
rect 24124 11154 24176 11160
rect 24676 11212 24728 11218
rect 24676 11154 24728 11160
rect 23848 11008 23900 11014
rect 23848 10950 23900 10956
rect 23860 10674 23888 10950
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 23756 10600 23808 10606
rect 23756 10542 23808 10548
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 23492 10062 23520 10406
rect 23480 10056 23532 10062
rect 23478 10024 23480 10033
rect 23532 10024 23534 10033
rect 23478 9959 23534 9968
rect 23480 9444 23532 9450
rect 23480 9386 23532 9392
rect 23492 8294 23520 9386
rect 23572 8968 23624 8974
rect 23572 8910 23624 8916
rect 23480 8288 23532 8294
rect 23386 8256 23442 8265
rect 23480 8230 23532 8236
rect 23386 8191 23442 8200
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23492 7546 23520 7890
rect 23584 7750 23612 8910
rect 23572 7744 23624 7750
rect 23572 7686 23624 7692
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 23204 5364 23256 5370
rect 23204 5306 23256 5312
rect 22940 5222 23152 5250
rect 23124 5030 23152 5222
rect 23112 5024 23164 5030
rect 23112 4966 23164 4972
rect 22928 4752 22980 4758
rect 22848 4712 22928 4740
rect 22848 4214 22876 4712
rect 22928 4694 22980 4700
rect 23124 4690 23152 4966
rect 23216 4826 23244 5306
rect 23676 5137 23704 10542
rect 23768 10130 23796 10542
rect 24136 10266 24164 11154
rect 24124 10260 24176 10266
rect 24124 10202 24176 10208
rect 23756 10124 23808 10130
rect 23756 10066 23808 10072
rect 24216 9988 24268 9994
rect 24216 9930 24268 9936
rect 23848 9648 23900 9654
rect 23848 9590 23900 9596
rect 23860 9217 23888 9590
rect 24030 9480 24086 9489
rect 24030 9415 24086 9424
rect 23846 9208 23902 9217
rect 23846 9143 23902 9152
rect 23940 8356 23992 8362
rect 23940 8298 23992 8304
rect 23952 8129 23980 8298
rect 23938 8120 23994 8129
rect 23938 8055 23994 8064
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 23952 6458 23980 6938
rect 23940 6452 23992 6458
rect 23940 6394 23992 6400
rect 23662 5128 23718 5137
rect 23662 5063 23718 5072
rect 23204 4820 23256 4826
rect 23204 4762 23256 4768
rect 23112 4684 23164 4690
rect 23112 4626 23164 4632
rect 23216 4214 23244 4762
rect 22836 4208 22888 4214
rect 22836 4150 22888 4156
rect 23204 4208 23256 4214
rect 23204 4150 23256 4156
rect 24044 4078 24072 9415
rect 24228 8838 24256 9930
rect 24308 9920 24360 9926
rect 24308 9862 24360 9868
rect 24320 9761 24348 9862
rect 24306 9752 24362 9761
rect 24306 9687 24362 9696
rect 24320 9489 24348 9687
rect 24688 9586 24716 11154
rect 24964 10713 24992 11494
rect 25134 11384 25190 11393
rect 25134 11319 25136 11328
rect 25188 11319 25190 11328
rect 25136 11290 25188 11296
rect 24950 10704 25006 10713
rect 24950 10639 25006 10648
rect 25136 10600 25188 10606
rect 25136 10542 25188 10548
rect 24952 10124 25004 10130
rect 24952 10066 25004 10072
rect 24768 9920 24820 9926
rect 24768 9862 24820 9868
rect 24676 9580 24728 9586
rect 24676 9522 24728 9528
rect 24306 9480 24362 9489
rect 24306 9415 24308 9424
rect 24360 9415 24362 9424
rect 24308 9386 24360 9392
rect 24780 9092 24808 9862
rect 24964 9382 24992 10066
rect 25148 9722 25176 10542
rect 25240 10266 25268 13126
rect 25516 12986 25544 13398
rect 25688 13320 25740 13326
rect 25740 13280 25912 13308
rect 25688 13262 25740 13268
rect 25596 13184 25648 13190
rect 25596 13126 25648 13132
rect 25504 12980 25556 12986
rect 25504 12922 25556 12928
rect 25502 12336 25558 12345
rect 25502 12271 25504 12280
rect 25556 12271 25558 12280
rect 25504 12242 25556 12248
rect 25608 12170 25636 13126
rect 25884 12646 25912 13280
rect 25964 13252 26016 13258
rect 25964 13194 26016 13200
rect 26056 13252 26108 13258
rect 26056 13194 26108 13200
rect 25780 12640 25832 12646
rect 25780 12582 25832 12588
rect 25872 12640 25924 12646
rect 25872 12582 25924 12588
rect 25792 12374 25820 12582
rect 25780 12368 25832 12374
rect 25780 12310 25832 12316
rect 25596 12164 25648 12170
rect 25596 12106 25648 12112
rect 25688 12096 25740 12102
rect 25688 12038 25740 12044
rect 25320 11552 25372 11558
rect 25320 11494 25372 11500
rect 25332 11150 25360 11494
rect 25320 11144 25372 11150
rect 25700 11121 25728 12038
rect 25780 11620 25832 11626
rect 25780 11562 25832 11568
rect 25792 11354 25820 11562
rect 25780 11348 25832 11354
rect 25780 11290 25832 11296
rect 25884 11286 25912 12582
rect 25872 11280 25924 11286
rect 25872 11222 25924 11228
rect 25320 11086 25372 11092
rect 25686 11112 25742 11121
rect 25332 10606 25360 11086
rect 25686 11047 25742 11056
rect 25320 10600 25372 10606
rect 25320 10542 25372 10548
rect 25700 10538 25728 11047
rect 25976 10810 26004 13194
rect 26068 11257 26096 13194
rect 26620 13190 26648 13398
rect 27436 13320 27488 13326
rect 27066 13288 27122 13297
rect 27436 13262 27488 13268
rect 27988 13320 28040 13326
rect 27988 13262 28040 13268
rect 27066 13223 27122 13232
rect 27080 13190 27108 13223
rect 26608 13184 26660 13190
rect 26528 13144 26608 13172
rect 26238 13016 26294 13025
rect 26238 12951 26294 12960
rect 26252 12918 26280 12951
rect 26240 12912 26292 12918
rect 26240 12854 26292 12860
rect 26424 12708 26476 12714
rect 26424 12650 26476 12656
rect 26332 12436 26384 12442
rect 26332 12378 26384 12384
rect 26240 12368 26292 12374
rect 26240 12310 26292 12316
rect 26054 11248 26110 11257
rect 26054 11183 26110 11192
rect 25964 10804 26016 10810
rect 25964 10746 26016 10752
rect 26148 10804 26200 10810
rect 26148 10746 26200 10752
rect 25688 10532 25740 10538
rect 25688 10474 25740 10480
rect 25228 10260 25280 10266
rect 25228 10202 25280 10208
rect 25700 10198 25728 10474
rect 25688 10192 25740 10198
rect 25688 10134 25740 10140
rect 25320 10124 25372 10130
rect 25320 10066 25372 10072
rect 25332 9722 25360 10066
rect 25136 9716 25188 9722
rect 25136 9658 25188 9664
rect 25320 9716 25372 9722
rect 25320 9658 25372 9664
rect 25148 9450 25176 9658
rect 26160 9518 26188 10746
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25596 9512 25648 9518
rect 25596 9454 25648 9460
rect 26148 9512 26200 9518
rect 26148 9454 26200 9460
rect 25136 9444 25188 9450
rect 25136 9386 25188 9392
rect 24952 9376 25004 9382
rect 24952 9318 25004 9324
rect 24860 9104 24912 9110
rect 24780 9064 24860 9092
rect 24308 8968 24360 8974
rect 24308 8910 24360 8916
rect 24216 8832 24268 8838
rect 24216 8774 24268 8780
rect 24228 8498 24256 8774
rect 24320 8634 24348 8910
rect 24308 8628 24360 8634
rect 24308 8570 24360 8576
rect 24584 8628 24636 8634
rect 24584 8570 24636 8576
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 24228 8401 24256 8434
rect 24214 8392 24270 8401
rect 24214 8327 24270 8336
rect 24308 8288 24360 8294
rect 24308 8230 24360 8236
rect 24320 7750 24348 8230
rect 24308 7744 24360 7750
rect 24308 7686 24360 7692
rect 24214 7440 24270 7449
rect 24214 7375 24270 7384
rect 24228 6866 24256 7375
rect 24216 6860 24268 6866
rect 24216 6802 24268 6808
rect 24122 6624 24178 6633
rect 24122 6559 24178 6568
rect 24136 6458 24164 6559
rect 24124 6452 24176 6458
rect 24124 6394 24176 6400
rect 24320 5681 24348 7686
rect 24596 7546 24624 8570
rect 24780 8090 24808 9064
rect 24964 9081 24992 9318
rect 25240 9110 25268 9454
rect 25608 9178 25636 9454
rect 25596 9172 25648 9178
rect 25596 9114 25648 9120
rect 25228 9104 25280 9110
rect 24860 9046 24912 9052
rect 24950 9072 25006 9081
rect 25228 9046 25280 9052
rect 24950 9007 25006 9016
rect 26148 9036 26200 9042
rect 26148 8978 26200 8984
rect 25136 8968 25188 8974
rect 25136 8910 25188 8916
rect 25148 8634 25176 8910
rect 26160 8634 26188 8978
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 26148 8628 26200 8634
rect 26148 8570 26200 8576
rect 26148 8424 26200 8430
rect 26148 8366 26200 8372
rect 26160 8090 26188 8366
rect 24768 8084 24820 8090
rect 24768 8026 24820 8032
rect 26148 8084 26200 8090
rect 26148 8026 26200 8032
rect 25044 8016 25096 8022
rect 25044 7958 25096 7964
rect 25320 8016 25372 8022
rect 25320 7958 25372 7964
rect 24952 7948 25004 7954
rect 24952 7890 25004 7896
rect 24584 7540 24636 7546
rect 24584 7482 24636 7488
rect 24584 7336 24636 7342
rect 24584 7278 24636 7284
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 24596 7206 24624 7278
rect 24584 7200 24636 7206
rect 24584 7142 24636 7148
rect 24490 7032 24546 7041
rect 24688 7002 24716 7278
rect 24768 7200 24820 7206
rect 24820 7148 24900 7154
rect 24768 7142 24900 7148
rect 24780 7126 24900 7142
rect 24490 6967 24546 6976
rect 24676 6996 24728 7002
rect 24504 6322 24532 6967
rect 24676 6938 24728 6944
rect 24688 6322 24716 6938
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 24306 5672 24362 5681
rect 24306 5607 24362 5616
rect 24308 5568 24360 5574
rect 24308 5510 24360 5516
rect 24216 5228 24268 5234
rect 24216 5170 24268 5176
rect 24124 5024 24176 5030
rect 24124 4966 24176 4972
rect 24136 4554 24164 4966
rect 24124 4548 24176 4554
rect 24124 4490 24176 4496
rect 24032 4072 24084 4078
rect 24032 4014 24084 4020
rect 22008 4004 22060 4010
rect 22008 3946 22060 3952
rect 21916 3936 21968 3942
rect 21916 3878 21968 3884
rect 21928 3602 21956 3878
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 21640 3392 21692 3398
rect 21640 3334 21692 3340
rect 21652 3194 21680 3334
rect 21928 3194 21956 3538
rect 22020 3398 22048 3946
rect 24044 3738 24072 4014
rect 24032 3732 24084 3738
rect 24032 3674 24084 3680
rect 24228 3466 24256 5170
rect 24320 5098 24348 5510
rect 24504 5370 24532 6258
rect 24872 6254 24900 7126
rect 24964 6730 24992 7890
rect 24952 6724 25004 6730
rect 24952 6666 25004 6672
rect 24860 6248 24912 6254
rect 24582 6216 24638 6225
rect 24860 6190 24912 6196
rect 24582 6151 24584 6160
rect 24636 6151 24638 6160
rect 24584 6122 24636 6128
rect 24860 5704 24912 5710
rect 24674 5672 24730 5681
rect 24860 5646 24912 5652
rect 24674 5607 24730 5616
rect 24492 5364 24544 5370
rect 24492 5306 24544 5312
rect 24308 5092 24360 5098
rect 24308 5034 24360 5040
rect 24320 4486 24348 5034
rect 24308 4480 24360 4486
rect 24308 4422 24360 4428
rect 24320 4049 24348 4422
rect 24306 4040 24362 4049
rect 24306 3975 24308 3984
rect 24360 3975 24362 3984
rect 24308 3946 24360 3952
rect 24582 3768 24638 3777
rect 24582 3703 24584 3712
rect 24636 3703 24638 3712
rect 24584 3674 24636 3680
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 22008 3392 22060 3398
rect 23020 3392 23072 3398
rect 22008 3334 22060 3340
rect 23018 3360 23020 3369
rect 23072 3360 23074 3369
rect 23018 3295 23074 3304
rect 21640 3188 21692 3194
rect 21640 3130 21692 3136
rect 21916 3188 21968 3194
rect 21916 3130 21968 3136
rect 23032 3058 23060 3295
rect 24596 3058 24624 3674
rect 24688 3534 24716 5607
rect 24872 5250 24900 5646
rect 24780 5234 24900 5250
rect 24768 5228 24900 5234
rect 24820 5222 24900 5228
rect 24768 5170 24820 5176
rect 24860 4480 24912 4486
rect 24860 4422 24912 4428
rect 24872 4078 24900 4422
rect 24860 4072 24912 4078
rect 24860 4014 24912 4020
rect 24872 3738 24900 4014
rect 25056 4010 25084 7958
rect 25226 7848 25282 7857
rect 25226 7783 25282 7792
rect 25240 7177 25268 7783
rect 25332 7449 25360 7958
rect 25412 7880 25464 7886
rect 25412 7822 25464 7828
rect 25318 7440 25374 7449
rect 25318 7375 25374 7384
rect 25424 7342 25452 7822
rect 26252 7750 26280 12310
rect 26344 11354 26372 12378
rect 26436 12102 26464 12650
rect 26424 12096 26476 12102
rect 26424 12038 26476 12044
rect 26528 11898 26556 13144
rect 26608 13126 26660 13132
rect 26976 13184 27028 13190
rect 26976 13126 27028 13132
rect 27068 13184 27120 13190
rect 27068 13126 27120 13132
rect 26700 12776 26752 12782
rect 26620 12724 26700 12730
rect 26620 12718 26752 12724
rect 26620 12702 26740 12718
rect 26516 11892 26568 11898
rect 26516 11834 26568 11840
rect 26620 11801 26648 12702
rect 26988 12646 27016 13126
rect 26976 12640 27028 12646
rect 26976 12582 27028 12588
rect 27448 12238 27476 13262
rect 27804 12912 27856 12918
rect 27540 12860 27804 12866
rect 27540 12854 27856 12860
rect 27540 12838 27844 12854
rect 27540 12442 27568 12838
rect 27622 12540 27918 12560
rect 27678 12538 27702 12540
rect 27758 12538 27782 12540
rect 27838 12538 27862 12540
rect 27700 12486 27702 12538
rect 27764 12486 27776 12538
rect 27838 12486 27840 12538
rect 27678 12484 27702 12486
rect 27758 12484 27782 12486
rect 27838 12484 27862 12486
rect 27622 12464 27918 12484
rect 27528 12436 27580 12442
rect 27528 12378 27580 12384
rect 26976 12232 27028 12238
rect 27436 12232 27488 12238
rect 26976 12174 27028 12180
rect 27434 12200 27436 12209
rect 27488 12200 27490 12209
rect 26606 11792 26662 11801
rect 26606 11727 26662 11736
rect 26332 11348 26384 11354
rect 26332 11290 26384 11296
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 26528 10742 26556 11086
rect 26516 10736 26568 10742
rect 26516 10678 26568 10684
rect 26620 10146 26648 11727
rect 26988 11286 27016 12174
rect 27434 12135 27490 12144
rect 27448 12109 27476 12135
rect 27804 12096 27856 12102
rect 27802 12064 27804 12073
rect 27856 12064 27858 12073
rect 27802 11999 27858 12008
rect 27622 11452 27918 11472
rect 27678 11450 27702 11452
rect 27758 11450 27782 11452
rect 27838 11450 27862 11452
rect 27700 11398 27702 11450
rect 27764 11398 27776 11450
rect 27838 11398 27840 11450
rect 27678 11396 27702 11398
rect 27758 11396 27782 11398
rect 27838 11396 27862 11398
rect 27622 11376 27918 11396
rect 26976 11280 27028 11286
rect 26976 11222 27028 11228
rect 26790 10976 26846 10985
rect 26790 10911 26846 10920
rect 26436 10118 26648 10146
rect 26436 8362 26464 10118
rect 26516 10056 26568 10062
rect 26516 9998 26568 10004
rect 26528 8498 26556 9998
rect 26608 9444 26660 9450
rect 26608 9386 26660 9392
rect 26620 9110 26648 9386
rect 26608 9104 26660 9110
rect 26608 9046 26660 9052
rect 26620 8498 26648 9046
rect 26700 8832 26752 8838
rect 26700 8774 26752 8780
rect 26712 8537 26740 8774
rect 26698 8528 26754 8537
rect 26516 8492 26568 8498
rect 26516 8434 26568 8440
rect 26608 8492 26660 8498
rect 26698 8463 26754 8472
rect 26608 8434 26660 8440
rect 26424 8356 26476 8362
rect 26424 8298 26476 8304
rect 26700 8288 26752 8294
rect 26700 8230 26752 8236
rect 26240 7744 26292 7750
rect 26240 7686 26292 7692
rect 25964 7540 26016 7546
rect 25964 7482 26016 7488
rect 25412 7336 25464 7342
rect 25412 7278 25464 7284
rect 25226 7168 25282 7177
rect 25226 7103 25282 7112
rect 25240 6866 25268 7103
rect 25976 7002 26004 7482
rect 25964 6996 26016 7002
rect 25964 6938 26016 6944
rect 25228 6860 25280 6866
rect 25228 6802 25280 6808
rect 25240 6322 25268 6802
rect 25412 6792 25464 6798
rect 25412 6734 25464 6740
rect 25504 6792 25556 6798
rect 25504 6734 25556 6740
rect 25424 6497 25452 6734
rect 25410 6488 25466 6497
rect 25410 6423 25412 6432
rect 25464 6423 25466 6432
rect 25412 6394 25464 6400
rect 25228 6316 25280 6322
rect 25228 6258 25280 6264
rect 25424 5953 25452 6394
rect 25410 5944 25466 5953
rect 25516 5914 25544 6734
rect 25778 6488 25834 6497
rect 25778 6423 25834 6432
rect 25688 6248 25740 6254
rect 25688 6190 25740 6196
rect 25410 5879 25466 5888
rect 25504 5908 25556 5914
rect 25504 5850 25556 5856
rect 25700 5574 25728 6190
rect 25688 5568 25740 5574
rect 25594 5536 25650 5545
rect 25688 5510 25740 5516
rect 25594 5471 25650 5480
rect 25608 5370 25636 5471
rect 25596 5364 25648 5370
rect 25596 5306 25648 5312
rect 25318 4992 25374 5001
rect 25318 4927 25374 4936
rect 25332 4758 25360 4927
rect 25792 4758 25820 6423
rect 25976 6186 26004 6938
rect 26608 6656 26660 6662
rect 26608 6598 26660 6604
rect 26620 6225 26648 6598
rect 26606 6216 26662 6225
rect 25964 6180 26016 6186
rect 26606 6151 26662 6160
rect 25964 6122 26016 6128
rect 26056 5636 26108 5642
rect 26056 5578 26108 5584
rect 26068 5234 26096 5578
rect 26148 5568 26200 5574
rect 26200 5516 26280 5522
rect 26148 5510 26280 5516
rect 26160 5494 26280 5510
rect 26056 5228 26108 5234
rect 26056 5170 26108 5176
rect 25872 5092 25924 5098
rect 25872 5034 25924 5040
rect 25884 4826 25912 5034
rect 25872 4820 25924 4826
rect 25872 4762 25924 4768
rect 25320 4752 25372 4758
rect 25320 4694 25372 4700
rect 25780 4752 25832 4758
rect 25780 4694 25832 4700
rect 25136 4684 25188 4690
rect 25136 4626 25188 4632
rect 25148 4185 25176 4626
rect 25332 4214 25360 4694
rect 25792 4282 25820 4694
rect 26252 4622 26280 5494
rect 26608 5364 26660 5370
rect 26608 5306 26660 5312
rect 26240 4616 26292 4622
rect 26240 4558 26292 4564
rect 25780 4276 25832 4282
rect 25780 4218 25832 4224
rect 25320 4208 25372 4214
rect 25134 4176 25190 4185
rect 25134 4111 25136 4120
rect 25188 4111 25190 4120
rect 25318 4176 25320 4185
rect 25372 4176 25374 4185
rect 25318 4111 25374 4120
rect 25136 4082 25188 4088
rect 25044 4004 25096 4010
rect 25044 3946 25096 3952
rect 24860 3732 24912 3738
rect 24860 3674 24912 3680
rect 24768 3664 24820 3670
rect 24768 3606 24820 3612
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 24688 3194 24716 3470
rect 24780 3194 24808 3606
rect 24950 3360 25006 3369
rect 24950 3295 25006 3304
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24768 3188 24820 3194
rect 24768 3130 24820 3136
rect 23020 3052 23072 3058
rect 23020 2994 23072 3000
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 18878 2887 18934 2896
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 20640 2650 20668 2858
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 17222 1456 17278 1465
rect 17222 1391 17278 1400
rect 24964 480 24992 3295
rect 25148 1737 25176 4082
rect 25792 3670 25820 4218
rect 26620 3777 26648 5306
rect 26712 4214 26740 8230
rect 26804 6866 26832 10911
rect 26882 10704 26938 10713
rect 26882 10639 26938 10648
rect 26896 10305 26924 10639
rect 26882 10296 26938 10305
rect 26988 10266 27016 11222
rect 28000 11218 28028 13262
rect 28448 12844 28500 12850
rect 28448 12786 28500 12792
rect 28356 12708 28408 12714
rect 28356 12650 28408 12656
rect 28264 12640 28316 12646
rect 28184 12600 28264 12628
rect 27988 11212 28040 11218
rect 27988 11154 28040 11160
rect 27894 11112 27950 11121
rect 27894 11047 27896 11056
rect 27948 11047 27950 11056
rect 27896 11018 27948 11024
rect 27160 10736 27212 10742
rect 27160 10678 27212 10684
rect 26882 10231 26938 10240
rect 26976 10260 27028 10266
rect 26976 10202 27028 10208
rect 27172 9722 27200 10678
rect 27622 10364 27918 10384
rect 27678 10362 27702 10364
rect 27758 10362 27782 10364
rect 27838 10362 27862 10364
rect 27700 10310 27702 10362
rect 27764 10310 27776 10362
rect 27838 10310 27840 10362
rect 27678 10308 27702 10310
rect 27758 10308 27782 10310
rect 27838 10308 27862 10310
rect 27622 10288 27918 10308
rect 27528 10192 27580 10198
rect 27528 10134 27580 10140
rect 27160 9716 27212 9722
rect 27160 9658 27212 9664
rect 27540 9654 27568 10134
rect 28184 10062 28212 12600
rect 28264 12582 28316 12588
rect 28264 12436 28316 12442
rect 28264 12378 28316 12384
rect 28276 11626 28304 12378
rect 28368 12374 28396 12650
rect 28356 12368 28408 12374
rect 28354 12336 28356 12345
rect 28408 12336 28410 12345
rect 28354 12271 28410 12280
rect 28368 11830 28396 12271
rect 28460 12170 28488 12786
rect 28448 12164 28500 12170
rect 28448 12106 28500 12112
rect 28356 11824 28408 11830
rect 28356 11766 28408 11772
rect 28264 11620 28316 11626
rect 28264 11562 28316 11568
rect 28368 11354 28396 11766
rect 28356 11348 28408 11354
rect 28356 11290 28408 11296
rect 28356 11008 28408 11014
rect 28356 10950 28408 10956
rect 28368 10470 28396 10950
rect 28356 10464 28408 10470
rect 28356 10406 28408 10412
rect 28368 10062 28396 10406
rect 28172 10056 28224 10062
rect 28172 9998 28224 10004
rect 28356 10056 28408 10062
rect 28356 9998 28408 10004
rect 27988 9920 28040 9926
rect 27988 9862 28040 9868
rect 27528 9648 27580 9654
rect 27528 9590 27580 9596
rect 27622 9276 27918 9296
rect 27678 9274 27702 9276
rect 27758 9274 27782 9276
rect 27838 9274 27862 9276
rect 27700 9222 27702 9274
rect 27764 9222 27776 9274
rect 27838 9222 27840 9274
rect 27678 9220 27702 9222
rect 27758 9220 27782 9222
rect 27838 9220 27862 9222
rect 27158 9208 27214 9217
rect 27622 9200 27918 9220
rect 28000 9178 28028 9862
rect 28184 9625 28212 9998
rect 28170 9616 28226 9625
rect 28170 9551 28226 9560
rect 28184 9382 28212 9551
rect 28368 9450 28396 9998
rect 28552 9722 28580 13466
rect 28736 13394 28764 15520
rect 31220 13734 31248 15520
rect 32864 13932 32916 13938
rect 32864 13874 32916 13880
rect 31760 13864 31812 13870
rect 31760 13806 31812 13812
rect 30932 13728 30984 13734
rect 30932 13670 30984 13676
rect 31208 13728 31260 13734
rect 31208 13670 31260 13676
rect 31668 13728 31720 13734
rect 31668 13670 31720 13676
rect 28908 13456 28960 13462
rect 28908 13398 28960 13404
rect 28724 13388 28776 13394
rect 28724 13330 28776 13336
rect 28920 13190 28948 13398
rect 30104 13388 30156 13394
rect 30104 13330 30156 13336
rect 28908 13184 28960 13190
rect 28908 13126 28960 13132
rect 29000 13184 29052 13190
rect 29000 13126 29052 13132
rect 29828 13184 29880 13190
rect 29828 13126 29880 13132
rect 28920 12918 28948 13126
rect 28908 12912 28960 12918
rect 28908 12854 28960 12860
rect 29012 12238 29040 13126
rect 29368 12980 29420 12986
rect 29368 12922 29420 12928
rect 29460 12980 29512 12986
rect 29460 12922 29512 12928
rect 29092 12708 29144 12714
rect 29092 12650 29144 12656
rect 28816 12232 28868 12238
rect 29000 12232 29052 12238
rect 28816 12174 28868 12180
rect 28998 12200 29000 12209
rect 29052 12200 29054 12209
rect 28632 12164 28684 12170
rect 28632 12106 28684 12112
rect 28644 11286 28672 12106
rect 28828 11558 28856 12174
rect 28998 12135 29054 12144
rect 29012 12109 29040 12135
rect 29104 11778 29132 12650
rect 29380 12170 29408 12922
rect 29368 12164 29420 12170
rect 29368 12106 29420 12112
rect 29472 11898 29500 12922
rect 29736 12912 29788 12918
rect 29736 12854 29788 12860
rect 29644 12640 29696 12646
rect 29644 12582 29696 12588
rect 29460 11892 29512 11898
rect 29460 11834 29512 11840
rect 28920 11762 29132 11778
rect 28908 11756 29132 11762
rect 28960 11750 29132 11756
rect 28908 11698 28960 11704
rect 29184 11688 29236 11694
rect 29184 11630 29236 11636
rect 28908 11620 28960 11626
rect 28908 11562 28960 11568
rect 28816 11552 28868 11558
rect 28816 11494 28868 11500
rect 28632 11280 28684 11286
rect 28632 11222 28684 11228
rect 28644 10470 28672 11222
rect 28632 10464 28684 10470
rect 28632 10406 28684 10412
rect 28540 9716 28592 9722
rect 28540 9658 28592 9664
rect 28356 9444 28408 9450
rect 28356 9386 28408 9392
rect 28172 9376 28224 9382
rect 28172 9318 28224 9324
rect 27158 9143 27160 9152
rect 27212 9143 27214 9152
rect 27988 9172 28040 9178
rect 27160 9114 27212 9120
rect 27988 9114 28040 9120
rect 27434 9072 27490 9081
rect 27434 9007 27490 9016
rect 27252 8968 27304 8974
rect 27252 8910 27304 8916
rect 27264 8430 27292 8910
rect 27252 8424 27304 8430
rect 27252 8366 27304 8372
rect 27068 8356 27120 8362
rect 27068 8298 27120 8304
rect 26976 7880 27028 7886
rect 26882 7848 26938 7857
rect 26976 7822 27028 7828
rect 26882 7783 26938 7792
rect 26896 7313 26924 7783
rect 26882 7304 26938 7313
rect 26882 7239 26938 7248
rect 26884 7200 26936 7206
rect 26884 7142 26936 7148
rect 26792 6860 26844 6866
rect 26792 6802 26844 6808
rect 26804 5914 26832 6802
rect 26896 6361 26924 7142
rect 26988 6633 27016 7822
rect 27080 7721 27108 8298
rect 27342 8256 27398 8265
rect 27342 8191 27398 8200
rect 27066 7712 27122 7721
rect 27066 7647 27122 7656
rect 27160 7472 27212 7478
rect 27160 7414 27212 7420
rect 27172 7041 27200 7414
rect 27252 7268 27304 7274
rect 27252 7210 27304 7216
rect 27158 7032 27214 7041
rect 27264 7002 27292 7210
rect 27158 6967 27214 6976
rect 27252 6996 27304 7002
rect 27252 6938 27304 6944
rect 27068 6860 27120 6866
rect 27068 6802 27120 6808
rect 27080 6769 27108 6802
rect 27356 6769 27384 8191
rect 27066 6760 27122 6769
rect 27066 6695 27122 6704
rect 27342 6760 27398 6769
rect 27342 6695 27398 6704
rect 26974 6624 27030 6633
rect 26974 6559 27030 6568
rect 27080 6458 27108 6695
rect 27068 6452 27120 6458
rect 27068 6394 27120 6400
rect 26882 6352 26938 6361
rect 26882 6287 26938 6296
rect 26976 6112 27028 6118
rect 26976 6054 27028 6060
rect 26792 5908 26844 5914
rect 26792 5850 26844 5856
rect 26804 5273 26832 5850
rect 26988 5778 27016 6054
rect 27448 5914 27476 9007
rect 28000 8344 28028 9114
rect 28172 8492 28224 8498
rect 28172 8434 28224 8440
rect 28080 8356 28132 8362
rect 28000 8316 28080 8344
rect 28080 8298 28132 8304
rect 27622 8188 27918 8208
rect 27678 8186 27702 8188
rect 27758 8186 27782 8188
rect 27838 8186 27862 8188
rect 27700 8134 27702 8186
rect 27764 8134 27776 8186
rect 27838 8134 27840 8186
rect 27678 8132 27702 8134
rect 27758 8132 27782 8134
rect 27838 8132 27862 8134
rect 27622 8112 27918 8132
rect 28184 8090 28212 8434
rect 28264 8356 28316 8362
rect 28264 8298 28316 8304
rect 28172 8084 28224 8090
rect 28172 8026 28224 8032
rect 28080 7880 28132 7886
rect 28080 7822 28132 7828
rect 28092 7546 28120 7822
rect 28276 7750 28304 8298
rect 28356 8288 28408 8294
rect 28356 8230 28408 8236
rect 28446 8256 28502 8265
rect 28368 8129 28396 8230
rect 28446 8191 28502 8200
rect 28354 8120 28410 8129
rect 28354 8055 28410 8064
rect 28264 7744 28316 7750
rect 28264 7686 28316 7692
rect 28080 7540 28132 7546
rect 28080 7482 28132 7488
rect 27988 7268 28040 7274
rect 27988 7210 28040 7216
rect 27622 7100 27918 7120
rect 27678 7098 27702 7100
rect 27758 7098 27782 7100
rect 27838 7098 27862 7100
rect 27700 7046 27702 7098
rect 27764 7046 27776 7098
rect 27838 7046 27840 7098
rect 27678 7044 27702 7046
rect 27758 7044 27782 7046
rect 27838 7044 27862 7046
rect 27622 7024 27918 7044
rect 28000 6882 28028 7210
rect 27816 6854 28028 6882
rect 27816 6798 27844 6854
rect 27804 6792 27856 6798
rect 27804 6734 27856 6740
rect 27816 6390 27844 6734
rect 27896 6656 27948 6662
rect 27894 6624 27896 6633
rect 27948 6624 27950 6633
rect 27894 6559 27950 6568
rect 27804 6384 27856 6390
rect 27804 6326 27856 6332
rect 27622 6012 27918 6032
rect 27678 6010 27702 6012
rect 27758 6010 27782 6012
rect 27838 6010 27862 6012
rect 27700 5958 27702 6010
rect 27764 5958 27776 6010
rect 27838 5958 27840 6010
rect 27678 5956 27702 5958
rect 27758 5956 27782 5958
rect 27838 5956 27862 5958
rect 27622 5936 27918 5956
rect 28170 5944 28226 5953
rect 27436 5908 27488 5914
rect 27356 5868 27436 5896
rect 26976 5772 27028 5778
rect 26976 5714 27028 5720
rect 27356 5370 27384 5868
rect 28170 5879 28226 5888
rect 27436 5850 27488 5856
rect 27712 5772 27764 5778
rect 27712 5714 27764 5720
rect 27436 5704 27488 5710
rect 27434 5672 27436 5681
rect 27488 5672 27490 5681
rect 27434 5607 27490 5616
rect 27434 5400 27490 5409
rect 27344 5364 27396 5370
rect 27434 5335 27490 5344
rect 27344 5306 27396 5312
rect 26790 5264 26846 5273
rect 26790 5199 26846 5208
rect 27344 5092 27396 5098
rect 27448 5080 27476 5335
rect 27724 5234 27752 5714
rect 28184 5710 28212 5879
rect 28460 5778 28488 8191
rect 28448 5772 28500 5778
rect 28448 5714 28500 5720
rect 28172 5704 28224 5710
rect 28172 5646 28224 5652
rect 28184 5370 28212 5646
rect 28172 5364 28224 5370
rect 28172 5306 28224 5312
rect 27712 5228 27764 5234
rect 27712 5170 27764 5176
rect 27724 5080 27752 5170
rect 28460 5137 28488 5714
rect 27396 5052 27476 5080
rect 27540 5052 27752 5080
rect 28446 5128 28502 5137
rect 28446 5063 28448 5072
rect 27344 5034 27396 5040
rect 27356 4690 27384 5034
rect 27540 4758 27568 5052
rect 28500 5063 28502 5072
rect 28448 5034 28500 5040
rect 28552 5030 28580 9658
rect 28644 7313 28672 10406
rect 28828 10062 28856 11494
rect 28816 10056 28868 10062
rect 28816 9998 28868 10004
rect 28920 9586 28948 11562
rect 29092 11348 29144 11354
rect 29092 11290 29144 11296
rect 29000 11076 29052 11082
rect 29000 11018 29052 11024
rect 28908 9580 28960 9586
rect 28908 9522 28960 9528
rect 28724 9036 28776 9042
rect 28724 8978 28776 8984
rect 28736 8566 28764 8978
rect 29012 8922 29040 11018
rect 29104 10538 29132 11290
rect 29196 11218 29224 11630
rect 29184 11212 29236 11218
rect 29184 11154 29236 11160
rect 29092 10532 29144 10538
rect 29092 10474 29144 10480
rect 29196 10470 29224 11154
rect 29368 11008 29420 11014
rect 29368 10950 29420 10956
rect 29380 10606 29408 10950
rect 29368 10600 29420 10606
rect 29368 10542 29420 10548
rect 29184 10464 29236 10470
rect 29184 10406 29236 10412
rect 29196 10169 29224 10406
rect 29182 10160 29238 10169
rect 29182 10095 29238 10104
rect 29184 9920 29236 9926
rect 29184 9862 29236 9868
rect 29092 9444 29144 9450
rect 29092 9386 29144 9392
rect 29104 9217 29132 9386
rect 29196 9382 29224 9862
rect 29380 9654 29408 10542
rect 29368 9648 29420 9654
rect 29368 9590 29420 9596
rect 29276 9580 29328 9586
rect 29276 9522 29328 9528
rect 29184 9376 29236 9382
rect 29184 9318 29236 9324
rect 29090 9208 29146 9217
rect 29090 9143 29146 9152
rect 28828 8894 29040 8922
rect 28724 8560 28776 8566
rect 28724 8502 28776 8508
rect 28828 8498 28856 8894
rect 28908 8832 28960 8838
rect 28908 8774 28960 8780
rect 28920 8634 28948 8774
rect 28908 8628 28960 8634
rect 28908 8570 28960 8576
rect 28816 8492 28868 8498
rect 28816 8434 28868 8440
rect 28920 8430 28948 8570
rect 28908 8424 28960 8430
rect 28908 8366 28960 8372
rect 29104 8022 29132 9143
rect 29196 9042 29224 9318
rect 29184 9036 29236 9042
rect 29184 8978 29236 8984
rect 29184 8492 29236 8498
rect 29184 8434 29236 8440
rect 29092 8016 29144 8022
rect 29092 7958 29144 7964
rect 28724 7948 28776 7954
rect 28724 7890 28776 7896
rect 28736 7546 28764 7890
rect 28724 7540 28776 7546
rect 28724 7482 28776 7488
rect 29000 7404 29052 7410
rect 29000 7346 29052 7352
rect 28630 7304 28686 7313
rect 28630 7239 28686 7248
rect 29012 6798 29040 7346
rect 29104 6934 29132 7958
rect 29092 6928 29144 6934
rect 29092 6870 29144 6876
rect 29196 6866 29224 8434
rect 29288 7585 29316 9522
rect 29380 8974 29408 9590
rect 29368 8968 29420 8974
rect 29368 8910 29420 8916
rect 29552 8968 29604 8974
rect 29552 8910 29604 8916
rect 29564 8650 29592 8910
rect 29472 8634 29592 8650
rect 29472 8628 29604 8634
rect 29472 8622 29552 8628
rect 29368 8560 29420 8566
rect 29368 8502 29420 8508
rect 29380 8401 29408 8502
rect 29366 8392 29422 8401
rect 29366 8327 29422 8336
rect 29472 7954 29500 8622
rect 29552 8570 29604 8576
rect 29550 8528 29606 8537
rect 29550 8463 29606 8472
rect 29564 8362 29592 8463
rect 29552 8356 29604 8362
rect 29552 8298 29604 8304
rect 29460 7948 29512 7954
rect 29460 7890 29512 7896
rect 29274 7576 29330 7585
rect 29274 7511 29330 7520
rect 29184 6860 29236 6866
rect 29184 6802 29236 6808
rect 29368 6860 29420 6866
rect 29368 6802 29420 6808
rect 29000 6792 29052 6798
rect 29000 6734 29052 6740
rect 29012 6458 29040 6734
rect 28632 6452 28684 6458
rect 28632 6394 28684 6400
rect 29000 6452 29052 6458
rect 29000 6394 29052 6400
rect 28644 6089 28672 6394
rect 28998 6352 29054 6361
rect 28998 6287 29054 6296
rect 28908 6180 28960 6186
rect 28908 6122 28960 6128
rect 28630 6080 28686 6089
rect 28630 6015 28686 6024
rect 28632 5160 28684 5166
rect 28632 5102 28684 5108
rect 28540 5024 28592 5030
rect 28540 4966 28592 4972
rect 27622 4924 27918 4944
rect 27678 4922 27702 4924
rect 27758 4922 27782 4924
rect 27838 4922 27862 4924
rect 27700 4870 27702 4922
rect 27764 4870 27776 4922
rect 27838 4870 27840 4922
rect 27678 4868 27702 4870
rect 27758 4868 27782 4870
rect 27838 4868 27862 4870
rect 27622 4848 27918 4868
rect 28644 4826 28672 5102
rect 28632 4820 28684 4826
rect 28632 4762 28684 4768
rect 27528 4752 27580 4758
rect 27528 4694 27580 4700
rect 27344 4684 27396 4690
rect 27344 4626 27396 4632
rect 26792 4616 26844 4622
rect 26792 4558 26844 4564
rect 26804 4282 26832 4558
rect 26792 4276 26844 4282
rect 26792 4218 26844 4224
rect 26700 4208 26752 4214
rect 26700 4150 26752 4156
rect 27540 4146 27568 4694
rect 27528 4140 27580 4146
rect 27528 4082 27580 4088
rect 27344 4004 27396 4010
rect 27344 3946 27396 3952
rect 26606 3768 26662 3777
rect 26606 3703 26662 3712
rect 25780 3664 25832 3670
rect 25780 3606 25832 3612
rect 27356 3398 27384 3946
rect 27540 3738 27568 4082
rect 27622 3836 27918 3856
rect 27678 3834 27702 3836
rect 27758 3834 27782 3836
rect 27838 3834 27862 3836
rect 27700 3782 27702 3834
rect 27764 3782 27776 3834
rect 27838 3782 27840 3834
rect 27678 3780 27702 3782
rect 27758 3780 27782 3782
rect 27838 3780 27862 3782
rect 27622 3760 27918 3780
rect 28920 3754 28948 6122
rect 29012 5817 29040 6287
rect 29380 5846 29408 6802
rect 29184 5840 29236 5846
rect 28998 5808 29054 5817
rect 29184 5782 29236 5788
rect 29368 5840 29420 5846
rect 29368 5782 29420 5788
rect 28998 5743 29054 5752
rect 29000 5704 29052 5710
rect 29000 5646 29052 5652
rect 29012 5166 29040 5646
rect 29000 5160 29052 5166
rect 29000 5102 29052 5108
rect 29196 4486 29224 5782
rect 29656 4554 29684 12582
rect 29748 12220 29776 12854
rect 29840 12374 29868 13126
rect 30116 12889 30144 13330
rect 30380 13320 30432 13326
rect 30380 13262 30432 13268
rect 30102 12880 30158 12889
rect 30392 12850 30420 13262
rect 30654 12880 30710 12889
rect 30102 12815 30158 12824
rect 30196 12844 30248 12850
rect 30196 12786 30248 12792
rect 30380 12844 30432 12850
rect 30944 12850 30972 13670
rect 31208 13320 31260 13326
rect 31208 13262 31260 13268
rect 30654 12815 30656 12824
rect 30380 12786 30432 12792
rect 30708 12815 30710 12824
rect 30932 12844 30984 12850
rect 30656 12786 30708 12792
rect 30932 12786 30984 12792
rect 29920 12708 29972 12714
rect 29920 12650 29972 12656
rect 29932 12442 29960 12650
rect 29920 12436 29972 12442
rect 29920 12378 29972 12384
rect 29828 12368 29880 12374
rect 29828 12310 29880 12316
rect 30208 12306 30236 12786
rect 31220 12782 31248 13262
rect 31392 12912 31444 12918
rect 31392 12854 31444 12860
rect 31208 12776 31260 12782
rect 31208 12718 31260 12724
rect 30196 12300 30248 12306
rect 30196 12242 30248 12248
rect 30656 12300 30708 12306
rect 30656 12242 30708 12248
rect 29828 12232 29880 12238
rect 29748 12192 29828 12220
rect 29828 12174 29880 12180
rect 29920 12232 29972 12238
rect 29920 12174 29972 12180
rect 30564 12232 30616 12238
rect 30564 12174 30616 12180
rect 29840 11354 29868 12174
rect 29932 12073 29960 12174
rect 29918 12064 29974 12073
rect 29918 11999 29974 12008
rect 29932 11830 29960 11999
rect 30576 11937 30604 12174
rect 30562 11928 30618 11937
rect 30562 11863 30618 11872
rect 29920 11824 29972 11830
rect 29920 11766 29972 11772
rect 30380 11688 30432 11694
rect 30380 11630 30432 11636
rect 29828 11348 29880 11354
rect 29828 11290 29880 11296
rect 30392 11082 30420 11630
rect 30576 11558 30604 11863
rect 30668 11694 30696 12242
rect 30656 11688 30708 11694
rect 30656 11630 30708 11636
rect 30564 11552 30616 11558
rect 30564 11494 30616 11500
rect 30380 11076 30432 11082
rect 30380 11018 30432 11024
rect 30380 10464 30432 10470
rect 30208 10412 30380 10418
rect 30208 10406 30432 10412
rect 30208 10390 30420 10406
rect 29736 10056 29788 10062
rect 29736 9998 29788 10004
rect 29748 8838 29776 9998
rect 29736 8832 29788 8838
rect 29736 8774 29788 8780
rect 29748 6361 29776 8774
rect 30208 8265 30236 10390
rect 30288 9920 30340 9926
rect 30288 9862 30340 9868
rect 30300 9518 30328 9862
rect 30288 9512 30340 9518
rect 30288 9454 30340 9460
rect 30194 8256 30250 8265
rect 30194 8191 30250 8200
rect 30378 8256 30434 8265
rect 30378 8191 30434 8200
rect 30104 7744 30156 7750
rect 30104 7686 30156 7692
rect 30116 7342 30144 7686
rect 30104 7336 30156 7342
rect 30392 7313 30420 8191
rect 30104 7278 30156 7284
rect 30378 7304 30434 7313
rect 30378 7239 30434 7248
rect 30378 6760 30434 6769
rect 30378 6695 30434 6704
rect 30196 6384 30248 6390
rect 29734 6352 29790 6361
rect 30196 6326 30248 6332
rect 29734 6287 29790 6296
rect 29828 6316 29880 6322
rect 29828 6258 29880 6264
rect 29736 6112 29788 6118
rect 29736 6054 29788 6060
rect 29748 5545 29776 6054
rect 29840 5914 29868 6258
rect 29920 6248 29972 6254
rect 29920 6190 29972 6196
rect 29828 5908 29880 5914
rect 29828 5850 29880 5856
rect 29734 5536 29790 5545
rect 29734 5471 29790 5480
rect 29932 5234 29960 6190
rect 30104 5568 30156 5574
rect 30104 5510 30156 5516
rect 29920 5228 29972 5234
rect 29840 5188 29920 5216
rect 29840 4826 29868 5188
rect 29920 5170 29972 5176
rect 30116 5098 30144 5510
rect 29920 5092 29972 5098
rect 29920 5034 29972 5040
rect 30104 5092 30156 5098
rect 30104 5034 30156 5040
rect 29828 4820 29880 4826
rect 29828 4762 29880 4768
rect 29644 4548 29696 4554
rect 29644 4490 29696 4496
rect 29184 4480 29236 4486
rect 29184 4422 29236 4428
rect 29196 4282 29224 4422
rect 29932 4282 29960 5034
rect 30208 4826 30236 6326
rect 30392 5914 30420 6695
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30484 6497 30512 6598
rect 30470 6488 30526 6497
rect 30470 6423 30526 6432
rect 30380 5908 30432 5914
rect 30380 5850 30432 5856
rect 30392 5370 30420 5850
rect 30470 5808 30526 5817
rect 30470 5743 30526 5752
rect 30484 5710 30512 5743
rect 30472 5704 30524 5710
rect 30472 5646 30524 5652
rect 30380 5364 30432 5370
rect 30380 5306 30432 5312
rect 30288 5296 30340 5302
rect 30288 5238 30340 5244
rect 30196 4820 30248 4826
rect 30196 4762 30248 4768
rect 30300 4622 30328 5238
rect 30484 5030 30512 5646
rect 30576 5137 30604 11494
rect 30668 10810 30696 11630
rect 30932 11212 30984 11218
rect 30932 11154 30984 11160
rect 30656 10804 30708 10810
rect 30656 10746 30708 10752
rect 30944 10470 30972 11154
rect 30932 10464 30984 10470
rect 30932 10406 30984 10412
rect 30930 9208 30986 9217
rect 30930 9143 30932 9152
rect 30984 9143 30986 9152
rect 30932 9114 30984 9120
rect 30654 8528 30710 8537
rect 30654 8463 30710 8472
rect 30668 8090 30696 8463
rect 30932 8288 30984 8294
rect 30932 8230 30984 8236
rect 30656 8084 30708 8090
rect 30656 8026 30708 8032
rect 30656 7200 30708 7206
rect 30656 7142 30708 7148
rect 30668 6934 30696 7142
rect 30656 6928 30708 6934
rect 30656 6870 30708 6876
rect 30944 6730 30972 8230
rect 30932 6724 30984 6730
rect 30932 6666 30984 6672
rect 30748 6180 30800 6186
rect 30748 6122 30800 6128
rect 30760 5778 30788 6122
rect 30748 5772 30800 5778
rect 30748 5714 30800 5720
rect 30562 5128 30618 5137
rect 30562 5063 30618 5072
rect 30472 5024 30524 5030
rect 30378 4992 30434 5001
rect 30472 4966 30524 4972
rect 30378 4927 30434 4936
rect 30392 4758 30420 4927
rect 30380 4752 30432 4758
rect 30484 4729 30512 4966
rect 30760 4826 30788 5714
rect 30932 5364 30984 5370
rect 30932 5306 30984 5312
rect 30944 4865 30972 5306
rect 30930 4856 30986 4865
rect 30564 4820 30616 4826
rect 30564 4762 30616 4768
rect 30748 4820 30800 4826
rect 30930 4791 30986 4800
rect 30748 4762 30800 4768
rect 30380 4694 30432 4700
rect 30470 4720 30526 4729
rect 30288 4616 30340 4622
rect 30288 4558 30340 4564
rect 30392 4570 30420 4694
rect 30470 4655 30526 4664
rect 30300 4468 30328 4558
rect 30392 4542 30512 4570
rect 30300 4440 30420 4468
rect 29184 4276 29236 4282
rect 29184 4218 29236 4224
rect 29920 4276 29972 4282
rect 29920 4218 29972 4224
rect 30196 4004 30248 4010
rect 30196 3946 30248 3952
rect 29644 3936 29696 3942
rect 29644 3878 29696 3884
rect 28920 3738 29040 3754
rect 27528 3732 27580 3738
rect 28920 3732 29052 3738
rect 28920 3726 29000 3732
rect 27528 3674 27580 3680
rect 29000 3674 29052 3680
rect 29656 3641 29684 3878
rect 30208 3738 30236 3946
rect 30392 3738 30420 4440
rect 30484 4214 30512 4542
rect 30472 4208 30524 4214
rect 30472 4150 30524 4156
rect 30576 4146 30604 4762
rect 30564 4140 30616 4146
rect 30564 4082 30616 4088
rect 30760 4078 30788 4762
rect 31116 4480 31168 4486
rect 31116 4422 31168 4428
rect 31128 4282 31156 4422
rect 31116 4276 31168 4282
rect 31116 4218 31168 4224
rect 30748 4072 30800 4078
rect 30562 4040 30618 4049
rect 30748 4014 30800 4020
rect 30562 3975 30618 3984
rect 30576 3942 30604 3975
rect 30564 3936 30616 3942
rect 30564 3878 30616 3884
rect 30196 3732 30248 3738
rect 30196 3674 30248 3680
rect 30380 3732 30432 3738
rect 30380 3674 30432 3680
rect 30760 3670 30788 4014
rect 31220 3777 31248 12718
rect 31404 12442 31432 12854
rect 31680 12850 31708 13670
rect 31772 13530 31800 13806
rect 31760 13524 31812 13530
rect 31760 13466 31812 13472
rect 32128 13388 32180 13394
rect 32128 13330 32180 13336
rect 31668 12844 31720 12850
rect 31668 12786 31720 12792
rect 32140 12782 32168 13330
rect 32128 12776 32180 12782
rect 32128 12718 32180 12724
rect 31760 12708 31812 12714
rect 31680 12668 31760 12696
rect 31680 12442 31708 12668
rect 31760 12650 31812 12656
rect 32876 12442 32904 13874
rect 33416 13388 33468 13394
rect 33416 13330 33468 13336
rect 33428 12646 33456 13330
rect 33600 12844 33652 12850
rect 33600 12786 33652 12792
rect 33416 12640 33468 12646
rect 33416 12582 33468 12588
rect 31392 12436 31444 12442
rect 31392 12378 31444 12384
rect 31668 12436 31720 12442
rect 31668 12378 31720 12384
rect 32864 12436 32916 12442
rect 32864 12378 32916 12384
rect 31680 12345 31708 12378
rect 31666 12336 31722 12345
rect 31666 12271 31722 12280
rect 32680 12300 32732 12306
rect 32680 12242 32732 12248
rect 31298 12200 31354 12209
rect 31298 12135 31354 12144
rect 31312 8498 31340 12135
rect 31758 12064 31814 12073
rect 31758 11999 31814 12008
rect 31772 11898 31800 11999
rect 31760 11892 31812 11898
rect 31760 11834 31812 11840
rect 32692 11558 32720 12242
rect 33324 12096 33376 12102
rect 33324 12038 33376 12044
rect 33336 11626 33364 12038
rect 33324 11620 33376 11626
rect 33324 11562 33376 11568
rect 32404 11552 32456 11558
rect 32404 11494 32456 11500
rect 32680 11552 32732 11558
rect 32680 11494 32732 11500
rect 32310 11384 32366 11393
rect 32310 11319 32366 11328
rect 32324 10742 32352 11319
rect 32416 11082 32444 11494
rect 32404 11076 32456 11082
rect 32404 11018 32456 11024
rect 32692 10985 32720 11494
rect 33048 11144 33100 11150
rect 33048 11086 33100 11092
rect 33324 11144 33376 11150
rect 33324 11086 33376 11092
rect 32678 10976 32734 10985
rect 32678 10911 32734 10920
rect 32312 10736 32364 10742
rect 32126 10704 32182 10713
rect 32312 10678 32364 10684
rect 32954 10704 33010 10713
rect 32126 10639 32182 10648
rect 33060 10690 33088 11086
rect 33336 10810 33364 11086
rect 33324 10804 33376 10810
rect 33324 10746 33376 10752
rect 33060 10674 33180 10690
rect 33060 10668 33192 10674
rect 33060 10662 33140 10668
rect 32954 10639 33010 10648
rect 32140 10606 32168 10639
rect 32128 10600 32180 10606
rect 32128 10542 32180 10548
rect 31668 10532 31720 10538
rect 31668 10474 31720 10480
rect 31680 9897 31708 10474
rect 32968 10470 32996 10639
rect 33140 10610 33192 10616
rect 32956 10464 33008 10470
rect 32956 10406 33008 10412
rect 33324 10464 33376 10470
rect 33324 10406 33376 10412
rect 31760 10260 31812 10266
rect 31760 10202 31812 10208
rect 31666 9888 31722 9897
rect 31666 9823 31722 9832
rect 31300 8492 31352 8498
rect 31300 8434 31352 8440
rect 31772 7313 31800 10202
rect 32968 10198 32996 10406
rect 32956 10192 33008 10198
rect 32956 10134 33008 10140
rect 33048 10192 33100 10198
rect 33048 10134 33100 10140
rect 32126 9616 32182 9625
rect 33060 9586 33088 10134
rect 32126 9551 32182 9560
rect 33048 9580 33100 9586
rect 32140 9518 32168 9551
rect 33048 9522 33100 9528
rect 32128 9512 32180 9518
rect 32128 9454 32180 9460
rect 32312 9376 32364 9382
rect 32310 9344 32312 9353
rect 32772 9376 32824 9382
rect 32364 9344 32366 9353
rect 32772 9318 32824 9324
rect 32310 9279 32366 9288
rect 32784 9217 32812 9318
rect 32770 9208 32826 9217
rect 32770 9143 32826 9152
rect 31852 9104 31904 9110
rect 31852 9046 31904 9052
rect 31864 8362 31892 9046
rect 32956 9036 33008 9042
rect 32956 8978 33008 8984
rect 31852 8356 31904 8362
rect 31852 8298 31904 8304
rect 32588 8356 32640 8362
rect 32588 8298 32640 8304
rect 31758 7304 31814 7313
rect 31758 7239 31814 7248
rect 31864 5642 31892 8298
rect 32600 7818 32628 8298
rect 32588 7812 32640 7818
rect 32588 7754 32640 7760
rect 32312 7404 32364 7410
rect 32312 7346 32364 7352
rect 32324 7002 32352 7346
rect 32312 6996 32364 7002
rect 32312 6938 32364 6944
rect 32324 6254 32352 6938
rect 32312 6248 32364 6254
rect 32312 6190 32364 6196
rect 32128 6112 32180 6118
rect 32128 6054 32180 6060
rect 31852 5636 31904 5642
rect 31852 5578 31904 5584
rect 32140 5234 32168 6054
rect 32862 5944 32918 5953
rect 32862 5879 32918 5888
rect 32128 5228 32180 5234
rect 32128 5170 32180 5176
rect 32140 4826 32168 5170
rect 32128 4820 32180 4826
rect 32128 4762 32180 4768
rect 32876 4729 32904 5879
rect 32862 4720 32918 4729
rect 32862 4655 32918 4664
rect 32968 4554 32996 8978
rect 33060 8430 33088 9522
rect 33232 8968 33284 8974
rect 33232 8910 33284 8916
rect 33140 8832 33192 8838
rect 33140 8774 33192 8780
rect 33048 8424 33100 8430
rect 33048 8366 33100 8372
rect 33060 7954 33088 8366
rect 33048 7948 33100 7954
rect 33048 7890 33100 7896
rect 33060 7546 33088 7890
rect 33048 7540 33100 7546
rect 33048 7482 33100 7488
rect 33046 7440 33102 7449
rect 33046 7375 33102 7384
rect 33060 7274 33088 7375
rect 33048 7268 33100 7274
rect 33048 7210 33100 7216
rect 33060 6202 33088 7210
rect 33152 6866 33180 8774
rect 33244 8362 33272 8910
rect 33232 8356 33284 8362
rect 33232 8298 33284 8304
rect 33244 8022 33272 8298
rect 33232 8016 33284 8022
rect 33232 7958 33284 7964
rect 33244 7546 33272 7958
rect 33232 7540 33284 7546
rect 33232 7482 33284 7488
rect 33230 7304 33286 7313
rect 33230 7239 33286 7248
rect 33140 6860 33192 6866
rect 33140 6802 33192 6808
rect 33152 6458 33180 6802
rect 33140 6452 33192 6458
rect 33140 6394 33192 6400
rect 33244 6322 33272 7239
rect 33232 6316 33284 6322
rect 33232 6258 33284 6264
rect 33060 6174 33272 6202
rect 33046 5944 33102 5953
rect 33046 5879 33102 5888
rect 33140 5908 33192 5914
rect 33060 5846 33088 5879
rect 33140 5850 33192 5856
rect 33048 5840 33100 5846
rect 33048 5782 33100 5788
rect 33152 5386 33180 5850
rect 33244 5846 33272 6174
rect 33232 5840 33284 5846
rect 33232 5782 33284 5788
rect 33060 5370 33180 5386
rect 33048 5364 33180 5370
rect 33100 5358 33180 5364
rect 33048 5306 33100 5312
rect 33244 5250 33272 5782
rect 33152 5222 33272 5250
rect 33152 4826 33180 5222
rect 33230 5128 33286 5137
rect 33230 5063 33286 5072
rect 33140 4820 33192 4826
rect 33140 4762 33192 4768
rect 32956 4548 33008 4554
rect 32956 4490 33008 4496
rect 33152 4282 33180 4762
rect 33244 4758 33272 5063
rect 33232 4752 33284 4758
rect 33336 4729 33364 10406
rect 33428 5817 33456 12582
rect 33508 11144 33560 11150
rect 33508 11086 33560 11092
rect 33520 10713 33548 11086
rect 33506 10704 33562 10713
rect 33506 10639 33562 10648
rect 33612 10538 33640 12786
rect 33704 12209 33732 15520
rect 35806 15464 35862 15473
rect 35806 15399 35862 15408
rect 34518 15056 34574 15065
rect 34518 14991 34574 15000
rect 34532 13530 34560 14991
rect 34702 14648 34758 14657
rect 34702 14583 34758 14592
rect 34612 13864 34664 13870
rect 34610 13832 34612 13841
rect 34664 13832 34666 13841
rect 34610 13767 34666 13776
rect 34520 13524 34572 13530
rect 34520 13466 34572 13472
rect 34152 13388 34204 13394
rect 34152 13330 34204 13336
rect 34164 12628 34192 13330
rect 34716 13258 34744 14583
rect 34794 14240 34850 14249
rect 34794 14175 34850 14184
rect 34808 13938 34836 14175
rect 34796 13932 34848 13938
rect 34796 13874 34848 13880
rect 35164 13796 35216 13802
rect 35164 13738 35216 13744
rect 35072 13456 35124 13462
rect 34794 13424 34850 13433
rect 35072 13398 35124 13404
rect 34794 13359 34850 13368
rect 34704 13252 34756 13258
rect 34704 13194 34756 13200
rect 34289 13084 34585 13104
rect 34345 13082 34369 13084
rect 34425 13082 34449 13084
rect 34505 13082 34529 13084
rect 34367 13030 34369 13082
rect 34431 13030 34443 13082
rect 34505 13030 34507 13082
rect 34345 13028 34369 13030
rect 34425 13028 34449 13030
rect 34505 13028 34529 13030
rect 34289 13008 34585 13028
rect 34612 12980 34664 12986
rect 34612 12922 34664 12928
rect 34244 12640 34296 12646
rect 34164 12600 34244 12628
rect 34624 12617 34652 12922
rect 34808 12918 34836 13359
rect 34796 12912 34848 12918
rect 35084 12900 35112 13398
rect 34796 12854 34848 12860
rect 34992 12872 35112 12900
rect 34796 12640 34848 12646
rect 34244 12582 34296 12588
rect 34610 12608 34666 12617
rect 34060 12368 34112 12374
rect 34058 12336 34060 12345
rect 34112 12336 34114 12345
rect 33784 12300 33836 12306
rect 34058 12271 34114 12280
rect 33784 12242 33836 12248
rect 33690 12200 33746 12209
rect 33690 12135 33746 12144
rect 33692 12096 33744 12102
rect 33692 12038 33744 12044
rect 33704 11762 33732 12038
rect 33796 11898 33824 12242
rect 34256 12209 34284 12582
rect 34796 12582 34848 12588
rect 34610 12543 34666 12552
rect 34242 12200 34298 12209
rect 34242 12135 34298 12144
rect 34289 11996 34585 12016
rect 34345 11994 34369 11996
rect 34425 11994 34449 11996
rect 34505 11994 34529 11996
rect 34367 11942 34369 11994
rect 34431 11942 34443 11994
rect 34505 11942 34507 11994
rect 34345 11940 34369 11942
rect 34425 11940 34449 11942
rect 34505 11940 34529 11942
rect 34289 11920 34585 11940
rect 33784 11892 33836 11898
rect 33784 11834 33836 11840
rect 33692 11756 33744 11762
rect 33692 11698 33744 11704
rect 33704 11529 33732 11698
rect 34808 11665 34836 12582
rect 34992 12424 35020 12872
rect 35176 12832 35204 13738
rect 35532 13388 35584 13394
rect 35532 13330 35584 13336
rect 35544 12850 35572 13330
rect 35624 13184 35676 13190
rect 35624 13126 35676 13132
rect 34900 12396 35020 12424
rect 35084 12804 35204 12832
rect 35532 12844 35584 12850
rect 34794 11656 34850 11665
rect 33784 11620 33836 11626
rect 34794 11591 34850 11600
rect 33784 11562 33836 11568
rect 33690 11520 33746 11529
rect 33690 11455 33746 11464
rect 33600 10532 33652 10538
rect 33600 10474 33652 10480
rect 33796 9926 33824 11562
rect 34704 11552 34756 11558
rect 34704 11494 34756 11500
rect 34428 11280 34480 11286
rect 34480 11228 34652 11234
rect 34428 11222 34652 11228
rect 34440 11206 34652 11222
rect 34716 11218 34744 11494
rect 33876 11008 33928 11014
rect 33876 10950 33928 10956
rect 33888 10470 33916 10950
rect 34289 10908 34585 10928
rect 34345 10906 34369 10908
rect 34425 10906 34449 10908
rect 34505 10906 34529 10908
rect 34367 10854 34369 10906
rect 34431 10854 34443 10906
rect 34505 10854 34507 10906
rect 34345 10852 34369 10854
rect 34425 10852 34449 10854
rect 34505 10852 34529 10854
rect 34289 10832 34585 10852
rect 33876 10464 33928 10470
rect 34336 10464 34388 10470
rect 33876 10406 33928 10412
rect 34334 10432 34336 10441
rect 34388 10432 34390 10441
rect 34334 10367 34390 10376
rect 33784 9920 33836 9926
rect 33784 9862 33836 9868
rect 34289 9820 34585 9840
rect 34345 9818 34369 9820
rect 34425 9818 34449 9820
rect 34505 9818 34529 9820
rect 34367 9766 34369 9818
rect 34431 9766 34443 9818
rect 34505 9766 34507 9818
rect 34345 9764 34369 9766
rect 34425 9764 34449 9766
rect 34505 9764 34529 9766
rect 34289 9744 34585 9764
rect 34624 9654 34652 11206
rect 34704 11212 34756 11218
rect 34704 11154 34756 11160
rect 34716 10674 34744 11154
rect 34808 10810 34836 11591
rect 34796 10804 34848 10810
rect 34796 10746 34848 10752
rect 34900 10690 34928 12396
rect 34980 12300 35032 12306
rect 34980 12242 35032 12248
rect 34992 11558 35020 12242
rect 34980 11552 35032 11558
rect 34980 11494 35032 11500
rect 34704 10668 34756 10674
rect 34704 10610 34756 10616
rect 34808 10662 34928 10690
rect 33968 9648 34020 9654
rect 33968 9590 34020 9596
rect 34612 9648 34664 9654
rect 34612 9590 34664 9596
rect 33784 9580 33836 9586
rect 33784 9522 33836 9528
rect 33690 9480 33746 9489
rect 33508 9444 33560 9450
rect 33690 9415 33746 9424
rect 33508 9386 33560 9392
rect 33520 8838 33548 9386
rect 33704 9194 33732 9415
rect 33796 9382 33824 9522
rect 33876 9444 33928 9450
rect 33876 9386 33928 9392
rect 33784 9376 33836 9382
rect 33784 9318 33836 9324
rect 33704 9166 33824 9194
rect 33508 8832 33560 8838
rect 33508 8774 33560 8780
rect 33414 5808 33470 5817
rect 33414 5743 33470 5752
rect 33414 5672 33470 5681
rect 33414 5607 33470 5616
rect 33428 4826 33456 5607
rect 33520 5409 33548 8774
rect 33690 8120 33746 8129
rect 33690 8055 33746 8064
rect 33600 7744 33652 7750
rect 33600 7686 33652 7692
rect 33612 6934 33640 7686
rect 33704 7313 33732 8055
rect 33796 7698 33824 9166
rect 33888 9042 33916 9386
rect 33876 9036 33928 9042
rect 33876 8978 33928 8984
rect 33888 8634 33916 8978
rect 33980 8974 34008 9590
rect 34428 9376 34480 9382
rect 34428 9318 34480 9324
rect 34612 9376 34664 9382
rect 34612 9318 34664 9324
rect 34440 9042 34468 9318
rect 34624 9081 34652 9318
rect 34702 9208 34758 9217
rect 34702 9143 34758 9152
rect 34610 9072 34666 9081
rect 34428 9036 34480 9042
rect 34610 9007 34666 9016
rect 34428 8978 34480 8984
rect 33968 8968 34020 8974
rect 33968 8910 34020 8916
rect 33876 8628 33928 8634
rect 33876 8570 33928 8576
rect 33980 8430 34008 8910
rect 34060 8832 34112 8838
rect 34060 8774 34112 8780
rect 34072 8498 34100 8774
rect 34289 8732 34585 8752
rect 34345 8730 34369 8732
rect 34425 8730 34449 8732
rect 34505 8730 34529 8732
rect 34367 8678 34369 8730
rect 34431 8678 34443 8730
rect 34505 8678 34507 8730
rect 34345 8676 34369 8678
rect 34425 8676 34449 8678
rect 34505 8676 34529 8678
rect 34289 8656 34585 8676
rect 34152 8560 34204 8566
rect 34152 8502 34204 8508
rect 34060 8492 34112 8498
rect 34060 8434 34112 8440
rect 33968 8424 34020 8430
rect 33968 8366 34020 8372
rect 33966 8120 34022 8129
rect 33966 8055 34022 8064
rect 33980 7857 34008 8055
rect 33966 7848 34022 7857
rect 33966 7783 34022 7792
rect 33796 7670 34008 7698
rect 33784 7540 33836 7546
rect 33784 7482 33836 7488
rect 33690 7304 33746 7313
rect 33690 7239 33746 7248
rect 33692 7200 33744 7206
rect 33692 7142 33744 7148
rect 33600 6928 33652 6934
rect 33600 6870 33652 6876
rect 33704 6882 33732 7142
rect 33796 7002 33824 7482
rect 33980 7206 34008 7670
rect 33968 7200 34020 7206
rect 33968 7142 34020 7148
rect 33784 6996 33836 7002
rect 33784 6938 33836 6944
rect 33612 6390 33640 6870
rect 33704 6854 33824 6882
rect 33692 6792 33744 6798
rect 33692 6734 33744 6740
rect 33600 6384 33652 6390
rect 33600 6326 33652 6332
rect 33704 5846 33732 6734
rect 33692 5840 33744 5846
rect 33692 5782 33744 5788
rect 33506 5400 33562 5409
rect 33506 5335 33562 5344
rect 33692 5024 33744 5030
rect 33690 4992 33692 5001
rect 33744 4992 33746 5001
rect 33690 4927 33746 4936
rect 33416 4820 33468 4826
rect 33416 4762 33468 4768
rect 33232 4694 33284 4700
rect 33322 4720 33378 4729
rect 33140 4276 33192 4282
rect 33140 4218 33192 4224
rect 33244 4214 33272 4694
rect 33322 4655 33378 4664
rect 33428 4282 33456 4762
rect 33796 4593 33824 6854
rect 34060 6860 34112 6866
rect 34060 6802 34112 6808
rect 33876 6656 33928 6662
rect 33876 6598 33928 6604
rect 33888 5914 33916 6598
rect 34072 6458 34100 6802
rect 34164 6798 34192 8502
rect 34428 8424 34480 8430
rect 34480 8372 34652 8378
rect 34428 8366 34652 8372
rect 34440 8350 34652 8366
rect 34289 7644 34585 7664
rect 34345 7642 34369 7644
rect 34425 7642 34449 7644
rect 34505 7642 34529 7644
rect 34367 7590 34369 7642
rect 34431 7590 34443 7642
rect 34505 7590 34507 7642
rect 34345 7588 34369 7590
rect 34425 7588 34449 7590
rect 34505 7588 34529 7590
rect 34289 7568 34585 7588
rect 34336 7200 34388 7206
rect 34336 7142 34388 7148
rect 34348 6866 34376 7142
rect 34336 6860 34388 6866
rect 34336 6802 34388 6808
rect 34152 6792 34204 6798
rect 34152 6734 34204 6740
rect 34289 6556 34585 6576
rect 34345 6554 34369 6556
rect 34425 6554 34449 6556
rect 34505 6554 34529 6556
rect 34367 6502 34369 6554
rect 34431 6502 34443 6554
rect 34505 6502 34507 6554
rect 34345 6500 34369 6502
rect 34425 6500 34449 6502
rect 34505 6500 34529 6502
rect 34289 6480 34585 6500
rect 34060 6452 34112 6458
rect 34060 6394 34112 6400
rect 34624 6254 34652 8350
rect 34716 7206 34744 9143
rect 34808 7721 34836 10662
rect 34886 8256 34942 8265
rect 34886 8191 34942 8200
rect 34900 8090 34928 8191
rect 34992 8129 35020 11494
rect 34978 8120 35034 8129
rect 34888 8084 34940 8090
rect 35084 8090 35112 12804
rect 35532 12786 35584 12792
rect 35440 12776 35492 12782
rect 35440 12718 35492 12724
rect 35452 12646 35480 12718
rect 35440 12640 35492 12646
rect 35440 12582 35492 12588
rect 35636 12209 35664 13126
rect 35820 12986 35848 15399
rect 35898 13016 35954 13025
rect 35808 12980 35860 12986
rect 35898 12951 35954 12960
rect 35808 12922 35860 12928
rect 35622 12200 35678 12209
rect 35622 12135 35678 12144
rect 35624 12096 35676 12102
rect 35624 12038 35676 12044
rect 35256 11688 35308 11694
rect 35256 11630 35308 11636
rect 35164 11144 35216 11150
rect 35164 11086 35216 11092
rect 35176 10849 35204 11086
rect 35162 10840 35218 10849
rect 35162 10775 35218 10784
rect 35164 10056 35216 10062
rect 35164 9998 35216 10004
rect 35176 9722 35204 9998
rect 35164 9716 35216 9722
rect 35164 9658 35216 9664
rect 35268 9450 35296 11630
rect 35348 10532 35400 10538
rect 35348 10474 35400 10480
rect 35360 10198 35388 10474
rect 35440 10464 35492 10470
rect 35440 10406 35492 10412
rect 35452 10305 35480 10406
rect 35438 10296 35494 10305
rect 35438 10231 35494 10240
rect 35348 10192 35400 10198
rect 35348 10134 35400 10140
rect 35452 10010 35480 10231
rect 35532 10192 35584 10198
rect 35636 10169 35664 12038
rect 35808 11552 35860 11558
rect 35808 11494 35860 11500
rect 35716 11280 35768 11286
rect 35716 11222 35768 11228
rect 35728 10441 35756 11222
rect 35714 10432 35770 10441
rect 35714 10367 35770 10376
rect 35532 10134 35584 10140
rect 35622 10160 35678 10169
rect 35360 9982 35480 10010
rect 35360 9926 35388 9982
rect 35348 9920 35400 9926
rect 35348 9862 35400 9868
rect 35256 9444 35308 9450
rect 35256 9386 35308 9392
rect 34978 8055 35034 8064
rect 35072 8084 35124 8090
rect 34888 8026 34940 8032
rect 35072 8026 35124 8032
rect 34794 7712 34850 7721
rect 34794 7647 34850 7656
rect 34900 7342 34928 8026
rect 35256 7744 35308 7750
rect 35256 7686 35308 7692
rect 35360 7698 35388 9862
rect 35544 9518 35572 10134
rect 35622 10095 35678 10104
rect 35622 9752 35678 9761
rect 35622 9687 35678 9696
rect 35532 9512 35584 9518
rect 35532 9454 35584 9460
rect 35440 9444 35492 9450
rect 35440 9386 35492 9392
rect 35452 9178 35480 9386
rect 35440 9172 35492 9178
rect 35440 9114 35492 9120
rect 35544 8906 35572 9454
rect 35532 8900 35584 8906
rect 35532 8842 35584 8848
rect 35440 8356 35492 8362
rect 35440 8298 35492 8304
rect 35452 7818 35480 8298
rect 35440 7812 35492 7818
rect 35440 7754 35492 7760
rect 34980 7472 35032 7478
rect 35268 7449 35296 7686
rect 35360 7670 35480 7698
rect 34980 7414 35032 7420
rect 35254 7440 35310 7449
rect 34888 7336 34940 7342
rect 34888 7278 34940 7284
rect 34704 7200 34756 7206
rect 34704 7142 34756 7148
rect 34888 6928 34940 6934
rect 34886 6896 34888 6905
rect 34940 6896 34942 6905
rect 34886 6831 34942 6840
rect 34900 6322 34928 6831
rect 34888 6316 34940 6322
rect 34888 6258 34940 6264
rect 34060 6248 34112 6254
rect 34060 6190 34112 6196
rect 34612 6248 34664 6254
rect 34612 6190 34664 6196
rect 33876 5908 33928 5914
rect 33876 5850 33928 5856
rect 34072 5710 34100 6190
rect 34992 5953 35020 7414
rect 35254 7375 35310 7384
rect 35348 7336 35400 7342
rect 35348 7278 35400 7284
rect 35072 6792 35124 6798
rect 35072 6734 35124 6740
rect 35084 6361 35112 6734
rect 35256 6656 35308 6662
rect 35256 6598 35308 6604
rect 35070 6352 35126 6361
rect 35070 6287 35072 6296
rect 35124 6287 35126 6296
rect 35072 6258 35124 6264
rect 34978 5944 35034 5953
rect 34978 5879 35034 5888
rect 34152 5840 34204 5846
rect 34152 5782 34204 5788
rect 34060 5704 34112 5710
rect 34060 5646 34112 5652
rect 34072 5166 34100 5646
rect 34060 5160 34112 5166
rect 34060 5102 34112 5108
rect 34072 5030 34100 5102
rect 34164 5098 34192 5782
rect 35084 5522 35112 6258
rect 35268 6254 35296 6598
rect 35256 6248 35308 6254
rect 35256 6190 35308 6196
rect 35084 5494 35204 5522
rect 34289 5468 34585 5488
rect 34345 5466 34369 5468
rect 34425 5466 34449 5468
rect 34505 5466 34529 5468
rect 34367 5414 34369 5466
rect 34431 5414 34443 5466
rect 34505 5414 34507 5466
rect 34345 5412 34369 5414
rect 34425 5412 34449 5414
rect 34505 5412 34529 5414
rect 34289 5392 34585 5412
rect 34794 5264 34850 5273
rect 34794 5199 34850 5208
rect 34152 5092 34204 5098
rect 34152 5034 34204 5040
rect 34060 5024 34112 5030
rect 34060 4966 34112 4972
rect 34610 4720 34666 4729
rect 34610 4655 34666 4664
rect 33782 4584 33838 4593
rect 33782 4519 33838 4528
rect 34289 4380 34585 4400
rect 34345 4378 34369 4380
rect 34425 4378 34449 4380
rect 34505 4378 34529 4380
rect 34367 4326 34369 4378
rect 34431 4326 34443 4378
rect 34505 4326 34507 4378
rect 34345 4324 34369 4326
rect 34425 4324 34449 4326
rect 34505 4324 34529 4326
rect 34289 4304 34585 4324
rect 33416 4276 33468 4282
rect 33416 4218 33468 4224
rect 33232 4208 33284 4214
rect 33232 4150 33284 4156
rect 31206 3768 31262 3777
rect 31206 3703 31262 3712
rect 30748 3664 30800 3670
rect 29642 3632 29698 3641
rect 30748 3606 30800 3612
rect 29642 3567 29698 3576
rect 27344 3392 27396 3398
rect 27344 3334 27396 3340
rect 27356 2961 27384 3334
rect 34289 3292 34585 3312
rect 34345 3290 34369 3292
rect 34425 3290 34449 3292
rect 34505 3290 34529 3292
rect 34367 3238 34369 3290
rect 34431 3238 34443 3290
rect 34505 3238 34507 3290
rect 34345 3236 34369 3238
rect 34425 3236 34449 3238
rect 34505 3236 34529 3238
rect 34289 3216 34585 3236
rect 27342 2952 27398 2961
rect 27342 2887 27398 2896
rect 27622 2748 27918 2768
rect 27678 2746 27702 2748
rect 27758 2746 27782 2748
rect 27838 2746 27862 2748
rect 27700 2694 27702 2746
rect 27764 2694 27776 2746
rect 27838 2694 27840 2746
rect 27678 2692 27702 2694
rect 27758 2692 27782 2694
rect 27838 2692 27862 2694
rect 27622 2672 27918 2692
rect 34289 2204 34585 2224
rect 34345 2202 34369 2204
rect 34425 2202 34449 2204
rect 34505 2202 34529 2204
rect 34367 2150 34369 2202
rect 34431 2150 34443 2202
rect 34505 2150 34507 2202
rect 34345 2148 34369 2150
rect 34425 2148 34449 2150
rect 34505 2148 34529 2150
rect 34289 2128 34585 2148
rect 25134 1728 25190 1737
rect 25134 1663 25190 1672
rect 34624 921 34652 4655
rect 34610 912 34666 921
rect 34610 847 34666 856
rect 2686 232 2742 241
rect 2686 167 2742 176
rect 4986 0 5042 480
rect 14922 0 14978 480
rect 24950 0 25006 480
rect 34808 241 34836 5199
rect 34980 5024 35032 5030
rect 34980 4966 35032 4972
rect 34992 480 35020 4966
rect 35176 513 35204 5494
rect 35360 1329 35388 7278
rect 35452 5794 35480 7670
rect 35532 7268 35584 7274
rect 35532 7210 35584 7216
rect 35544 6866 35572 7210
rect 35532 6860 35584 6866
rect 35532 6802 35584 6808
rect 35544 6254 35572 6802
rect 35532 6248 35584 6254
rect 35532 6190 35584 6196
rect 35544 5914 35572 6190
rect 35532 5908 35584 5914
rect 35532 5850 35584 5856
rect 35452 5766 35572 5794
rect 35440 5160 35492 5166
rect 35440 5102 35492 5108
rect 35452 4185 35480 5102
rect 35438 4176 35494 4185
rect 35544 4162 35572 5766
rect 35636 5370 35664 9687
rect 35728 7449 35756 10367
rect 35820 9081 35848 11494
rect 35912 11354 35940 12951
rect 36188 12345 36216 15520
rect 36740 13530 36768 15807
rect 38658 15520 38714 16000
rect 36728 13524 36780 13530
rect 36728 13466 36780 13472
rect 36544 13388 36596 13394
rect 36544 13330 36596 13336
rect 36556 12986 36584 13330
rect 36544 12980 36596 12986
rect 36544 12922 36596 12928
rect 36556 12889 36584 12922
rect 36542 12880 36598 12889
rect 36542 12815 36598 12824
rect 36728 12640 36780 12646
rect 36728 12582 36780 12588
rect 36174 12336 36230 12345
rect 36174 12271 36230 12280
rect 36452 12300 36504 12306
rect 36452 12242 36504 12248
rect 36082 12064 36138 12073
rect 36082 11999 36138 12008
rect 35900 11348 35952 11354
rect 35900 11290 35952 11296
rect 35900 11008 35952 11014
rect 35900 10950 35952 10956
rect 35912 10674 35940 10950
rect 35900 10668 35952 10674
rect 35900 10610 35952 10616
rect 35806 9072 35862 9081
rect 35806 9007 35862 9016
rect 35900 9036 35952 9042
rect 35900 8978 35952 8984
rect 35912 8634 35940 8978
rect 35900 8628 35952 8634
rect 35900 8570 35952 8576
rect 35808 8492 35860 8498
rect 35860 8452 35940 8480
rect 35808 8434 35860 8440
rect 35806 7984 35862 7993
rect 35806 7919 35862 7928
rect 35714 7440 35770 7449
rect 35714 7375 35770 7384
rect 35714 6624 35770 6633
rect 35714 6559 35770 6568
rect 35624 5364 35676 5370
rect 35624 5306 35676 5312
rect 35622 4176 35678 4185
rect 35544 4134 35622 4162
rect 35438 4111 35494 4120
rect 35622 4111 35678 4120
rect 35728 4049 35756 6559
rect 35820 5817 35848 7919
rect 35912 7546 35940 8452
rect 36096 8022 36124 11999
rect 36268 11688 36320 11694
rect 36268 11630 36320 11636
rect 36176 11212 36228 11218
rect 36176 11154 36228 11160
rect 36188 10470 36216 11154
rect 36176 10464 36228 10470
rect 36176 10406 36228 10412
rect 35992 8016 36044 8022
rect 35992 7958 36044 7964
rect 36084 8016 36136 8022
rect 36084 7958 36136 7964
rect 36004 7721 36032 7958
rect 35990 7712 36046 7721
rect 35990 7647 36046 7656
rect 35900 7540 35952 7546
rect 35900 7482 35952 7488
rect 36004 7206 36032 7647
rect 36096 7478 36124 7958
rect 36084 7472 36136 7478
rect 36084 7414 36136 7420
rect 35992 7200 36044 7206
rect 35992 7142 36044 7148
rect 36084 6928 36136 6934
rect 36188 6905 36216 10406
rect 36280 7313 36308 11630
rect 36464 11558 36492 12242
rect 36740 11801 36768 12582
rect 37188 12096 37240 12102
rect 37188 12038 37240 12044
rect 36726 11792 36782 11801
rect 36726 11727 36782 11736
rect 36452 11552 36504 11558
rect 36728 11552 36780 11558
rect 36452 11494 36504 11500
rect 36542 11520 36598 11529
rect 36360 11076 36412 11082
rect 36360 11018 36412 11024
rect 36372 8537 36400 11018
rect 36358 8528 36414 8537
rect 36464 8514 36492 11494
rect 36728 11494 36780 11500
rect 36542 11455 36598 11464
rect 36556 10810 36584 11455
rect 36544 10804 36596 10810
rect 36544 10746 36596 10752
rect 36740 10577 36768 11494
rect 36818 11112 36874 11121
rect 36818 11047 36874 11056
rect 36726 10568 36782 10577
rect 36726 10503 36782 10512
rect 36636 8968 36688 8974
rect 36636 8910 36688 8916
rect 36464 8486 36584 8514
rect 36358 8463 36414 8472
rect 36452 8424 36504 8430
rect 36450 8392 36452 8401
rect 36504 8392 36506 8401
rect 36450 8327 36506 8336
rect 36556 8242 36584 8486
rect 36372 8214 36584 8242
rect 36266 7304 36322 7313
rect 36266 7239 36322 7248
rect 36372 6934 36400 8214
rect 36648 8090 36676 8910
rect 36832 8498 36860 11047
rect 36912 11008 36964 11014
rect 37200 10985 37228 12038
rect 38672 11121 38700 15520
rect 38658 11112 38714 11121
rect 38658 11047 38714 11056
rect 36912 10950 36964 10956
rect 37186 10976 37242 10985
rect 36924 10713 36952 10950
rect 37186 10911 37242 10920
rect 37554 10840 37610 10849
rect 37554 10775 37610 10784
rect 36910 10704 36966 10713
rect 36910 10639 36966 10648
rect 37096 10668 37148 10674
rect 36924 10470 36952 10639
rect 37096 10610 37148 10616
rect 36912 10464 36964 10470
rect 36912 10406 36964 10412
rect 36924 10266 36952 10406
rect 37108 10266 37136 10610
rect 36912 10260 36964 10266
rect 36912 10202 36964 10208
rect 37096 10260 37148 10266
rect 37096 10202 37148 10208
rect 37568 9586 37596 10775
rect 37556 9580 37608 9586
rect 37556 9522 37608 9528
rect 36912 9376 36964 9382
rect 36912 9318 36964 9324
rect 36820 8492 36872 8498
rect 36820 8434 36872 8440
rect 36924 8265 36952 9318
rect 36910 8256 36966 8265
rect 36910 8191 36966 8200
rect 36452 8084 36504 8090
rect 36452 8026 36504 8032
rect 36636 8084 36688 8090
rect 36636 8026 36688 8032
rect 36464 7274 36492 8026
rect 36544 7744 36596 7750
rect 36544 7686 36596 7692
rect 36556 7410 36584 7686
rect 36544 7404 36596 7410
rect 36544 7346 36596 7352
rect 36452 7268 36504 7274
rect 36452 7210 36504 7216
rect 36360 6928 36412 6934
rect 36084 6870 36136 6876
rect 36174 6896 36230 6905
rect 35992 6656 36044 6662
rect 35992 6598 36044 6604
rect 35898 6080 35954 6089
rect 35898 6015 35954 6024
rect 35806 5808 35862 5817
rect 35806 5743 35862 5752
rect 35912 5642 35940 6015
rect 36004 5681 36032 6598
rect 36096 6497 36124 6870
rect 36360 6870 36412 6876
rect 36174 6831 36230 6840
rect 36360 6792 36412 6798
rect 36360 6734 36412 6740
rect 36082 6488 36138 6497
rect 36082 6423 36138 6432
rect 36096 5914 36124 6423
rect 36084 5908 36136 5914
rect 36084 5850 36136 5856
rect 35990 5672 36046 5681
rect 35900 5636 35952 5642
rect 36372 5642 36400 6734
rect 36556 6662 36584 7346
rect 36648 7342 36676 8026
rect 36636 7336 36688 7342
rect 36636 7278 36688 7284
rect 37004 7268 37056 7274
rect 37004 7210 37056 7216
rect 36636 7200 36688 7206
rect 36636 7142 36688 7148
rect 36544 6656 36596 6662
rect 36544 6598 36596 6604
rect 36556 6458 36584 6598
rect 36544 6452 36596 6458
rect 36544 6394 36596 6400
rect 35990 5607 36046 5616
rect 36360 5636 36412 5642
rect 35900 5578 35952 5584
rect 36360 5578 36412 5584
rect 35912 5522 35940 5578
rect 35820 5494 35940 5522
rect 35714 4040 35770 4049
rect 35714 3975 35770 3984
rect 35820 2961 35848 5494
rect 36648 5409 36676 7142
rect 37016 7041 37044 7210
rect 37002 7032 37058 7041
rect 37002 6967 37058 6976
rect 36634 5400 36690 5409
rect 36634 5335 36690 5344
rect 35806 2952 35862 2961
rect 35806 2887 35862 2896
rect 35622 2136 35678 2145
rect 35622 2071 35678 2080
rect 35636 1465 35664 2071
rect 35622 1456 35678 1465
rect 35622 1391 35678 1400
rect 35346 1320 35402 1329
rect 35346 1255 35402 1264
rect 35162 504 35218 513
rect 34794 232 34850 241
rect 34794 167 34850 176
rect 34978 0 35034 480
rect 35162 439 35218 448
<< via2 >>
rect 3054 15816 3110 15872
rect 36726 15816 36782 15872
rect 3422 15408 3478 15464
rect 3330 15000 3386 15056
rect 1398 10104 1454 10160
rect 1582 11772 1584 11792
rect 1584 11772 1636 11792
rect 1636 11772 1638 11792
rect 1582 11736 1638 11772
rect 1858 11056 1914 11112
rect 1674 9560 1730 9616
rect 2778 13368 2834 13424
rect 2318 11192 2374 11248
rect 3422 11600 3478 11656
rect 2502 10260 2558 10296
rect 2502 10240 2504 10260
rect 2504 10240 2556 10260
rect 2556 10240 2558 10260
rect 2410 10004 2412 10024
rect 2412 10004 2464 10024
rect 2464 10004 2466 10024
rect 2410 9968 2466 10004
rect 1582 8200 1638 8256
rect 2042 6568 2098 6624
rect 2226 4120 2282 4176
rect 2410 4936 2466 4992
rect 2962 8200 3018 8256
rect 2594 7520 2650 7576
rect 3238 7112 3294 7168
rect 3146 5108 3148 5128
rect 3148 5108 3200 5128
rect 3200 5108 3202 5128
rect 3146 5072 3202 5108
rect 2502 4664 2558 4720
rect 1306 448 1362 504
rect 3146 1672 3202 1728
rect 4434 14592 4490 14648
rect 4066 14184 4122 14240
rect 4342 13776 4398 13832
rect 4158 12960 4214 13016
rect 4066 12552 4122 12608
rect 4250 12164 4306 12200
rect 4250 12144 4252 12164
rect 4252 12144 4304 12164
rect 4304 12144 4306 12164
rect 3698 11056 3754 11112
rect 3514 6976 3570 7032
rect 3514 5208 3570 5264
rect 3698 10376 3754 10432
rect 3974 10920 4030 10976
rect 4066 10512 4122 10568
rect 4066 9560 4122 9616
rect 4250 8880 4306 8936
rect 4158 8472 4214 8528
rect 3790 6860 3846 6896
rect 3790 6840 3792 6860
rect 3792 6840 3844 6860
rect 3844 6840 3846 6860
rect 3974 6976 4030 7032
rect 3698 5344 3754 5400
rect 4526 11872 4582 11928
rect 4802 11464 4858 11520
rect 4618 10240 4674 10296
rect 4526 9152 4582 9208
rect 4710 10104 4766 10160
rect 4618 8628 4674 8664
rect 4618 8608 4620 8628
rect 4620 8608 4672 8628
rect 4672 8608 4674 8628
rect 4894 11056 4950 11112
rect 4986 9968 5042 10024
rect 5170 12300 5226 12336
rect 5170 12280 5172 12300
rect 5172 12280 5224 12300
rect 5224 12280 5226 12300
rect 4894 7792 4950 7848
rect 7622 13082 7678 13084
rect 7702 13082 7758 13084
rect 7782 13082 7838 13084
rect 7862 13082 7918 13084
rect 7622 13030 7648 13082
rect 7648 13030 7678 13082
rect 7702 13030 7712 13082
rect 7712 13030 7758 13082
rect 7782 13030 7828 13082
rect 7828 13030 7838 13082
rect 7862 13030 7892 13082
rect 7892 13030 7918 13082
rect 7622 13028 7678 13030
rect 7702 13028 7758 13030
rect 7782 13028 7838 13030
rect 7862 13028 7918 13030
rect 6274 11756 6330 11792
rect 6274 11736 6276 11756
rect 6276 11736 6328 11756
rect 6328 11736 6330 11756
rect 5722 11328 5778 11384
rect 5906 11192 5962 11248
rect 5446 10412 5448 10432
rect 5448 10412 5500 10432
rect 5500 10412 5502 10432
rect 5446 10376 5502 10412
rect 5538 9596 5540 9616
rect 5540 9596 5592 9616
rect 5592 9596 5594 9616
rect 5538 9560 5594 9596
rect 6182 10240 6238 10296
rect 5814 9288 5870 9344
rect 6090 9052 6092 9072
rect 6092 9052 6144 9072
rect 6144 9052 6146 9072
rect 6090 9016 6146 9052
rect 5998 8880 6054 8936
rect 5722 8356 5778 8392
rect 5722 8336 5724 8356
rect 5724 8336 5776 8356
rect 5776 8336 5778 8356
rect 6182 7828 6184 7848
rect 6184 7828 6236 7848
rect 6236 7828 6238 7848
rect 4802 7384 4858 7440
rect 6182 7792 6238 7828
rect 5906 7248 5962 7304
rect 6366 8472 6422 8528
rect 5814 6296 5870 6352
rect 4066 4800 4122 4856
rect 3606 4528 3662 4584
rect 3238 1264 3294 1320
rect 4066 4120 4122 4176
rect 3974 3848 4030 3904
rect 4894 4972 4896 4992
rect 4896 4972 4948 4992
rect 4948 4972 4950 4992
rect 4894 4936 4950 4972
rect 5078 4936 5134 4992
rect 6274 6452 6330 6488
rect 6274 6432 6276 6452
rect 6276 6432 6328 6452
rect 6328 6432 6330 6452
rect 6090 5908 6146 5944
rect 6090 5888 6092 5908
rect 6092 5888 6144 5908
rect 6144 5888 6146 5908
rect 4526 4004 4582 4040
rect 4526 3984 4528 4004
rect 4528 3984 4580 4004
rect 4580 3984 4582 4004
rect 6642 6160 6698 6216
rect 4618 3712 4674 3768
rect 3974 3304 4030 3360
rect 7622 11994 7678 11996
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7622 11942 7648 11994
rect 7648 11942 7678 11994
rect 7702 11942 7712 11994
rect 7712 11942 7758 11994
rect 7782 11942 7828 11994
rect 7828 11942 7838 11994
rect 7862 11942 7892 11994
rect 7892 11942 7918 11994
rect 7622 11940 7678 11942
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 9586 12144 9642 12200
rect 9126 11636 9128 11656
rect 9128 11636 9180 11656
rect 9180 11636 9182 11656
rect 9126 11600 9182 11636
rect 8942 11500 8944 11520
rect 8944 11500 8996 11520
rect 8996 11500 8998 11520
rect 7622 10906 7678 10908
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7622 10854 7648 10906
rect 7648 10854 7678 10906
rect 7702 10854 7712 10906
rect 7712 10854 7758 10906
rect 7782 10854 7828 10906
rect 7828 10854 7838 10906
rect 7862 10854 7892 10906
rect 7892 10854 7918 10906
rect 7622 10852 7678 10854
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 8942 11464 8998 11500
rect 8114 10784 8170 10840
rect 8022 10648 8078 10704
rect 8114 10512 8170 10568
rect 7102 8608 7158 8664
rect 5262 3052 5318 3088
rect 5262 3032 5264 3052
rect 5264 3032 5316 3052
rect 5316 3032 5318 3052
rect 4342 2508 4398 2544
rect 4342 2488 4344 2508
rect 4344 2488 4396 2508
rect 4396 2488 4398 2508
rect 3882 2080 3938 2136
rect 3790 856 3846 912
rect 7470 9968 7526 10024
rect 7622 9818 7678 9820
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7622 9766 7648 9818
rect 7648 9766 7678 9818
rect 7702 9766 7712 9818
rect 7712 9766 7758 9818
rect 7782 9766 7828 9818
rect 7828 9766 7838 9818
rect 7862 9766 7892 9818
rect 7892 9766 7918 9818
rect 7622 9764 7678 9766
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 8298 10376 8354 10432
rect 7654 9288 7710 9344
rect 7102 6704 7158 6760
rect 7622 8730 7678 8732
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7622 8678 7648 8730
rect 7648 8678 7678 8730
rect 7702 8678 7712 8730
rect 7712 8678 7758 8730
rect 7782 8678 7828 8730
rect 7828 8678 7838 8730
rect 7862 8678 7892 8730
rect 7892 8678 7918 8730
rect 7622 8676 7678 8678
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 8022 8608 8078 8664
rect 7746 8064 7802 8120
rect 7654 7928 7710 7984
rect 7622 7642 7678 7644
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7622 7590 7648 7642
rect 7648 7590 7678 7642
rect 7702 7590 7712 7642
rect 7712 7590 7758 7642
rect 7782 7590 7828 7642
rect 7828 7590 7838 7642
rect 7862 7590 7892 7642
rect 7892 7590 7918 7642
rect 7622 7588 7678 7590
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 7562 6704 7618 6760
rect 8206 7520 8262 7576
rect 8114 6976 8170 7032
rect 9770 11076 9826 11112
rect 9770 11056 9772 11076
rect 9772 11056 9824 11076
rect 9824 11056 9826 11076
rect 10230 10648 10286 10704
rect 9862 9832 9918 9888
rect 10138 10240 10194 10296
rect 10598 9152 10654 9208
rect 10230 8744 10286 8800
rect 9954 8508 9956 8528
rect 9956 8508 10008 8528
rect 10008 8508 10010 8528
rect 9954 8472 10010 8508
rect 9770 8336 9826 8392
rect 10414 8064 10470 8120
rect 8942 7248 8998 7304
rect 8298 6976 8354 7032
rect 10414 7148 10416 7168
rect 10416 7148 10468 7168
rect 10468 7148 10470 7168
rect 7622 6554 7678 6556
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7622 6502 7648 6554
rect 7648 6502 7678 6554
rect 7702 6502 7712 6554
rect 7712 6502 7758 6554
rect 7782 6502 7828 6554
rect 7828 6502 7838 6554
rect 7862 6502 7892 6554
rect 7892 6502 7918 6554
rect 7622 6500 7678 6502
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 7622 5466 7678 5468
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7622 5414 7648 5466
rect 7648 5414 7678 5466
rect 7702 5414 7712 5466
rect 7712 5414 7758 5466
rect 7782 5414 7828 5466
rect 7828 5414 7838 5466
rect 7862 5414 7892 5466
rect 7892 5414 7918 5466
rect 7622 5412 7678 5414
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 7194 3984 7250 4040
rect 7102 3732 7158 3768
rect 8114 5344 8170 5400
rect 9954 6704 10010 6760
rect 9862 6316 9918 6352
rect 9862 6296 9864 6316
rect 9864 6296 9916 6316
rect 9916 6296 9918 6316
rect 9678 5888 9734 5944
rect 9954 5752 10010 5808
rect 10414 7112 10470 7148
rect 10506 6704 10562 6760
rect 8758 5208 8814 5264
rect 8942 5092 8998 5128
rect 8942 5072 8944 5092
rect 8944 5072 8996 5092
rect 8996 5072 8998 5092
rect 7470 4528 7526 4584
rect 7622 4378 7678 4380
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7622 4326 7648 4378
rect 7648 4326 7678 4378
rect 7702 4326 7712 4378
rect 7712 4326 7758 4378
rect 7782 4326 7828 4378
rect 7828 4326 7838 4378
rect 7862 4326 7892 4378
rect 7892 4326 7918 4378
rect 7622 4324 7678 4326
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 8942 4120 8998 4176
rect 9218 4004 9274 4040
rect 9586 5092 9642 5128
rect 9586 5072 9588 5092
rect 9588 5072 9640 5092
rect 9640 5072 9642 5092
rect 9494 4800 9550 4856
rect 10322 5752 10378 5808
rect 10138 4564 10140 4584
rect 10140 4564 10192 4584
rect 10192 4564 10194 4584
rect 10138 4528 10194 4564
rect 9218 3984 9220 4004
rect 9220 3984 9272 4004
rect 9272 3984 9274 4004
rect 8666 3884 8668 3904
rect 8668 3884 8720 3904
rect 8720 3884 8722 3904
rect 8666 3848 8722 3884
rect 7102 3712 7104 3732
rect 7104 3712 7156 3732
rect 7156 3712 7158 3732
rect 9678 3304 9734 3360
rect 7622 3290 7678 3292
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7622 3238 7648 3290
rect 7648 3238 7678 3290
rect 7702 3238 7712 3290
rect 7712 3238 7758 3290
rect 7782 3238 7828 3290
rect 7828 3238 7838 3290
rect 7862 3238 7892 3290
rect 7892 3238 7918 3290
rect 7622 3236 7678 3238
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 12254 10920 12310 10976
rect 11150 9444 11206 9480
rect 11150 9424 11152 9444
rect 11152 9424 11204 9444
rect 11204 9424 11206 9444
rect 12070 10512 12126 10568
rect 11978 9968 12034 10024
rect 11426 9580 11482 9616
rect 11426 9560 11428 9580
rect 11428 9560 11480 9580
rect 11480 9560 11482 9580
rect 11426 9052 11428 9072
rect 11428 9052 11480 9072
rect 11480 9052 11482 9072
rect 11426 9016 11482 9052
rect 10966 8880 11022 8936
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 12806 11056 12862 11112
rect 12254 9288 12310 9344
rect 12530 8880 12586 8936
rect 12714 8880 12770 8936
rect 11794 8200 11850 8256
rect 11334 7812 11390 7848
rect 11334 7792 11336 7812
rect 11336 7792 11388 7812
rect 11388 7792 11390 7812
rect 10966 7656 11022 7712
rect 13542 11600 13598 11656
rect 13450 9560 13506 9616
rect 12990 9152 13046 9208
rect 12898 8608 12954 8664
rect 12530 8472 12586 8528
rect 11794 7248 11850 7304
rect 10966 6840 11022 6896
rect 11426 6296 11482 6352
rect 12438 6840 12494 6896
rect 12254 6704 12310 6760
rect 12162 6452 12218 6488
rect 12162 6432 12164 6452
rect 12164 6432 12216 6452
rect 12216 6432 12218 6452
rect 11426 5480 11482 5536
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 13818 9596 13820 9616
rect 13820 9596 13872 9616
rect 13872 9596 13874 9616
rect 13818 9560 13874 9596
rect 14186 10104 14242 10160
rect 14002 9560 14058 9616
rect 14002 9152 14058 9208
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 13818 8780 13820 8800
rect 13820 8780 13872 8800
rect 13872 8780 13874 8800
rect 13818 8744 13874 8780
rect 14278 8744 14334 8800
rect 15198 11736 15254 11792
rect 15382 11464 15438 11520
rect 15382 11192 15438 11248
rect 15198 9696 15254 9752
rect 14278 8472 14334 8528
rect 14462 8492 14518 8528
rect 14462 8472 14464 8492
rect 14464 8472 14516 8492
rect 14516 8472 14518 8492
rect 15382 8472 15438 8528
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 14646 7248 14702 7304
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 14646 6432 14702 6488
rect 14002 6332 14004 6352
rect 14004 6332 14056 6352
rect 14056 6332 14058 6352
rect 14002 6296 14058 6332
rect 14738 6296 14794 6352
rect 14002 6160 14058 6216
rect 14738 6024 14794 6080
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 15658 8356 15714 8392
rect 15658 8336 15660 8356
rect 15660 8336 15712 8356
rect 15712 8336 15714 8356
rect 15658 7656 15714 7712
rect 15474 7520 15530 7576
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 12530 4800 12586 4856
rect 16026 11600 16082 11656
rect 16210 12008 16266 12064
rect 16946 11600 17002 11656
rect 17958 12008 18014 12064
rect 16670 8880 16726 8936
rect 17130 8472 17186 8528
rect 17314 8236 17316 8256
rect 17316 8236 17368 8256
rect 17368 8236 17370 8256
rect 17314 8200 17370 8236
rect 16302 7828 16304 7848
rect 16304 7828 16356 7848
rect 16356 7828 16358 7848
rect 16302 7792 16358 7828
rect 16578 7404 16634 7440
rect 17038 7656 17094 7712
rect 16578 7384 16580 7404
rect 16580 7384 16632 7404
rect 16632 7384 16634 7404
rect 16670 7268 16726 7304
rect 16670 7248 16672 7268
rect 16672 7248 16724 7268
rect 16724 7248 16726 7268
rect 16210 6976 16266 7032
rect 16670 6432 16726 6488
rect 17038 6704 17094 6760
rect 16854 6024 16910 6080
rect 16486 5480 16542 5536
rect 16394 4820 16450 4856
rect 16394 4800 16396 4820
rect 16396 4800 16448 4820
rect 16448 4800 16450 4820
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 10322 2896 10378 2952
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 6918 2624 6974 2680
rect 14922 2488 14978 2544
rect 7622 2202 7678 2204
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7622 2150 7648 2202
rect 7648 2150 7678 2202
rect 7702 2150 7712 2202
rect 7712 2150 7758 2202
rect 7782 2150 7828 2202
rect 7828 2150 7838 2202
rect 7862 2150 7892 2202
rect 7892 2150 7918 2202
rect 7622 2148 7678 2150
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 17314 5752 17370 5808
rect 17406 5616 17462 5672
rect 18234 6296 18290 6352
rect 18142 6160 18198 6216
rect 17774 5364 17830 5400
rect 17774 5344 17776 5364
rect 17776 5344 17828 5364
rect 17828 5344 17830 5364
rect 18234 5616 18290 5672
rect 18142 4800 18198 4856
rect 18602 11736 18658 11792
rect 18694 11620 18750 11656
rect 18694 11600 18696 11620
rect 18696 11600 18748 11620
rect 18748 11600 18750 11620
rect 19982 11192 20038 11248
rect 18602 10920 18658 10976
rect 19062 10376 19118 10432
rect 18786 9968 18842 10024
rect 18602 9152 18658 9208
rect 19430 10240 19486 10296
rect 19062 8880 19118 8936
rect 18694 8336 18750 8392
rect 18602 6976 18658 7032
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 21454 11328 21510 11384
rect 27622 13626 27678 13628
rect 27702 13626 27758 13628
rect 27782 13626 27838 13628
rect 27862 13626 27918 13628
rect 27622 13574 27648 13626
rect 27648 13574 27678 13626
rect 27702 13574 27712 13626
rect 27712 13574 27758 13626
rect 27782 13574 27828 13626
rect 27828 13574 27838 13626
rect 27862 13574 27892 13626
rect 27892 13574 27918 13626
rect 27622 13572 27678 13574
rect 27702 13572 27758 13574
rect 27782 13572 27838 13574
rect 27862 13572 27918 13574
rect 24030 13232 24086 13288
rect 24030 12960 24086 13016
rect 22926 12144 22982 12200
rect 22926 11636 22928 11656
rect 22928 11636 22980 11656
rect 22980 11636 22982 11656
rect 22926 11600 22982 11636
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 20810 10512 20866 10568
rect 22190 10784 22246 10840
rect 20626 10376 20682 10432
rect 22190 10512 22246 10568
rect 22466 10512 22522 10568
rect 22282 10376 22338 10432
rect 20166 9832 20222 9888
rect 20074 9580 20130 9616
rect 20074 9560 20076 9580
rect 20076 9560 20128 9580
rect 20128 9560 20130 9580
rect 19798 8744 19854 8800
rect 19338 7692 19340 7712
rect 19340 7692 19392 7712
rect 19392 7692 19394 7712
rect 19338 7656 19394 7692
rect 19430 7520 19486 7576
rect 19614 7420 19616 7440
rect 19616 7420 19668 7440
rect 19668 7420 19670 7440
rect 19614 7384 19670 7420
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 21270 9016 21326 9072
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 21454 8356 21510 8392
rect 21454 8336 21456 8356
rect 21456 8336 21508 8356
rect 21508 8336 21510 8356
rect 20902 8236 20904 8256
rect 20904 8236 20956 8256
rect 20956 8236 20958 8256
rect 20902 8200 20958 8236
rect 21730 8472 21786 8528
rect 22374 9016 22430 9072
rect 22006 8472 22062 8528
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 21638 7520 21694 7576
rect 18878 6840 18934 6896
rect 18510 5228 18566 5264
rect 18510 5208 18512 5228
rect 18512 5208 18564 5228
rect 18564 5208 18566 5228
rect 18602 5092 18658 5128
rect 18602 5072 18604 5092
rect 18604 5072 18656 5092
rect 18656 5072 18658 5092
rect 18786 5072 18842 5128
rect 18602 4664 18658 4720
rect 18786 4256 18842 4312
rect 18326 3984 18382 4040
rect 17682 3576 17738 3632
rect 19522 5364 19578 5400
rect 19522 5344 19524 5364
rect 19524 5344 19576 5364
rect 19576 5344 19578 5364
rect 20166 6840 20222 6896
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 20810 6024 20866 6080
rect 22374 6860 22430 6896
rect 22374 6840 22376 6860
rect 22376 6840 22428 6860
rect 22428 6840 22430 6860
rect 21546 5752 21602 5808
rect 21822 5772 21878 5808
rect 21822 5752 21824 5772
rect 21824 5752 21876 5772
rect 21876 5752 21878 5772
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 19798 4664 19854 4720
rect 20442 3576 20498 3632
rect 19338 3304 19394 3360
rect 20534 3068 20536 3088
rect 20536 3068 20588 3088
rect 20588 3068 20590 3088
rect 20534 3032 20590 3068
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 21086 4020 21088 4040
rect 21088 4020 21140 4040
rect 21140 4020 21142 4040
rect 21086 3984 21142 4020
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 18878 2896 18934 2952
rect 22926 9152 22982 9208
rect 23294 12316 23296 12336
rect 23296 12316 23348 12336
rect 23348 12316 23350 12336
rect 23294 12280 23350 12316
rect 23202 8880 23258 8936
rect 24398 12044 24400 12064
rect 24400 12044 24452 12064
rect 24452 12044 24454 12064
rect 24398 12008 24454 12044
rect 24950 11872 25006 11928
rect 24674 11464 24730 11520
rect 23478 10004 23480 10024
rect 23480 10004 23532 10024
rect 23532 10004 23534 10024
rect 23478 9968 23534 10004
rect 23386 8200 23442 8256
rect 24030 9424 24086 9480
rect 23846 9152 23902 9208
rect 23938 8064 23994 8120
rect 23662 5072 23718 5128
rect 24306 9696 24362 9752
rect 25134 11348 25190 11384
rect 25134 11328 25136 11348
rect 25136 11328 25188 11348
rect 25188 11328 25190 11348
rect 24950 10648 25006 10704
rect 24306 9444 24362 9480
rect 24306 9424 24308 9444
rect 24308 9424 24360 9444
rect 24360 9424 24362 9444
rect 25502 12300 25558 12336
rect 25502 12280 25504 12300
rect 25504 12280 25556 12300
rect 25556 12280 25558 12300
rect 25686 11056 25742 11112
rect 27066 13232 27122 13288
rect 26238 12960 26294 13016
rect 26054 11192 26110 11248
rect 24214 8336 24270 8392
rect 24214 7384 24270 7440
rect 24122 6568 24178 6624
rect 24950 9016 25006 9072
rect 24490 6976 24546 7032
rect 24306 5616 24362 5672
rect 24582 6180 24638 6216
rect 24582 6160 24584 6180
rect 24584 6160 24636 6180
rect 24636 6160 24638 6180
rect 24674 5616 24730 5672
rect 24306 4004 24362 4040
rect 24306 3984 24308 4004
rect 24308 3984 24360 4004
rect 24360 3984 24362 4004
rect 24582 3732 24638 3768
rect 24582 3712 24584 3732
rect 24584 3712 24636 3732
rect 24636 3712 24638 3732
rect 23018 3340 23020 3360
rect 23020 3340 23072 3360
rect 23072 3340 23074 3360
rect 23018 3304 23074 3340
rect 25226 7792 25282 7848
rect 25318 7384 25374 7440
rect 27622 12538 27678 12540
rect 27702 12538 27758 12540
rect 27782 12538 27838 12540
rect 27862 12538 27918 12540
rect 27622 12486 27648 12538
rect 27648 12486 27678 12538
rect 27702 12486 27712 12538
rect 27712 12486 27758 12538
rect 27782 12486 27828 12538
rect 27828 12486 27838 12538
rect 27862 12486 27892 12538
rect 27892 12486 27918 12538
rect 27622 12484 27678 12486
rect 27702 12484 27758 12486
rect 27782 12484 27838 12486
rect 27862 12484 27918 12486
rect 27434 12180 27436 12200
rect 27436 12180 27488 12200
rect 27488 12180 27490 12200
rect 26606 11736 26662 11792
rect 27434 12144 27490 12180
rect 27802 12044 27804 12064
rect 27804 12044 27856 12064
rect 27856 12044 27858 12064
rect 27802 12008 27858 12044
rect 27622 11450 27678 11452
rect 27702 11450 27758 11452
rect 27782 11450 27838 11452
rect 27862 11450 27918 11452
rect 27622 11398 27648 11450
rect 27648 11398 27678 11450
rect 27702 11398 27712 11450
rect 27712 11398 27758 11450
rect 27782 11398 27828 11450
rect 27828 11398 27838 11450
rect 27862 11398 27892 11450
rect 27892 11398 27918 11450
rect 27622 11396 27678 11398
rect 27702 11396 27758 11398
rect 27782 11396 27838 11398
rect 27862 11396 27918 11398
rect 26790 10920 26846 10976
rect 26698 8472 26754 8528
rect 25226 7112 25282 7168
rect 25410 6452 25466 6488
rect 25410 6432 25412 6452
rect 25412 6432 25464 6452
rect 25464 6432 25466 6452
rect 25410 5888 25466 5944
rect 25778 6432 25834 6488
rect 25594 5480 25650 5536
rect 25318 4936 25374 4992
rect 26606 6160 26662 6216
rect 25134 4140 25190 4176
rect 25134 4120 25136 4140
rect 25136 4120 25188 4140
rect 25188 4120 25190 4140
rect 25318 4156 25320 4176
rect 25320 4156 25372 4176
rect 25372 4156 25374 4176
rect 25318 4120 25374 4156
rect 24950 3304 25006 3360
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 17222 1400 17278 1456
rect 26882 10648 26938 10704
rect 26882 10240 26938 10296
rect 27894 11076 27950 11112
rect 27894 11056 27896 11076
rect 27896 11056 27948 11076
rect 27948 11056 27950 11076
rect 27622 10362 27678 10364
rect 27702 10362 27758 10364
rect 27782 10362 27838 10364
rect 27862 10362 27918 10364
rect 27622 10310 27648 10362
rect 27648 10310 27678 10362
rect 27702 10310 27712 10362
rect 27712 10310 27758 10362
rect 27782 10310 27828 10362
rect 27828 10310 27838 10362
rect 27862 10310 27892 10362
rect 27892 10310 27918 10362
rect 27622 10308 27678 10310
rect 27702 10308 27758 10310
rect 27782 10308 27838 10310
rect 27862 10308 27918 10310
rect 28354 12316 28356 12336
rect 28356 12316 28408 12336
rect 28408 12316 28410 12336
rect 28354 12280 28410 12316
rect 27622 9274 27678 9276
rect 27702 9274 27758 9276
rect 27782 9274 27838 9276
rect 27862 9274 27918 9276
rect 27622 9222 27648 9274
rect 27648 9222 27678 9274
rect 27702 9222 27712 9274
rect 27712 9222 27758 9274
rect 27782 9222 27828 9274
rect 27828 9222 27838 9274
rect 27862 9222 27892 9274
rect 27892 9222 27918 9274
rect 27622 9220 27678 9222
rect 27702 9220 27758 9222
rect 27782 9220 27838 9222
rect 27862 9220 27918 9222
rect 27158 9172 27214 9208
rect 28170 9560 28226 9616
rect 28998 12180 29000 12200
rect 29000 12180 29052 12200
rect 29052 12180 29054 12200
rect 28998 12144 29054 12180
rect 27158 9152 27160 9172
rect 27160 9152 27212 9172
rect 27212 9152 27214 9172
rect 27434 9016 27490 9072
rect 26882 7792 26938 7848
rect 26882 7248 26938 7304
rect 27342 8200 27398 8256
rect 27066 7656 27122 7712
rect 27158 6976 27214 7032
rect 27066 6704 27122 6760
rect 27342 6704 27398 6760
rect 26974 6568 27030 6624
rect 26882 6296 26938 6352
rect 27622 8186 27678 8188
rect 27702 8186 27758 8188
rect 27782 8186 27838 8188
rect 27862 8186 27918 8188
rect 27622 8134 27648 8186
rect 27648 8134 27678 8186
rect 27702 8134 27712 8186
rect 27712 8134 27758 8186
rect 27782 8134 27828 8186
rect 27828 8134 27838 8186
rect 27862 8134 27892 8186
rect 27892 8134 27918 8186
rect 27622 8132 27678 8134
rect 27702 8132 27758 8134
rect 27782 8132 27838 8134
rect 27862 8132 27918 8134
rect 28446 8200 28502 8256
rect 28354 8064 28410 8120
rect 27622 7098 27678 7100
rect 27702 7098 27758 7100
rect 27782 7098 27838 7100
rect 27862 7098 27918 7100
rect 27622 7046 27648 7098
rect 27648 7046 27678 7098
rect 27702 7046 27712 7098
rect 27712 7046 27758 7098
rect 27782 7046 27828 7098
rect 27828 7046 27838 7098
rect 27862 7046 27892 7098
rect 27892 7046 27918 7098
rect 27622 7044 27678 7046
rect 27702 7044 27758 7046
rect 27782 7044 27838 7046
rect 27862 7044 27918 7046
rect 27894 6604 27896 6624
rect 27896 6604 27948 6624
rect 27948 6604 27950 6624
rect 27894 6568 27950 6604
rect 27622 6010 27678 6012
rect 27702 6010 27758 6012
rect 27782 6010 27838 6012
rect 27862 6010 27918 6012
rect 27622 5958 27648 6010
rect 27648 5958 27678 6010
rect 27702 5958 27712 6010
rect 27712 5958 27758 6010
rect 27782 5958 27828 6010
rect 27828 5958 27838 6010
rect 27862 5958 27892 6010
rect 27892 5958 27918 6010
rect 27622 5956 27678 5958
rect 27702 5956 27758 5958
rect 27782 5956 27838 5958
rect 27862 5956 27918 5958
rect 28170 5888 28226 5944
rect 27434 5652 27436 5672
rect 27436 5652 27488 5672
rect 27488 5652 27490 5672
rect 27434 5616 27490 5652
rect 27434 5344 27490 5400
rect 26790 5208 26846 5264
rect 28446 5092 28502 5128
rect 28446 5072 28448 5092
rect 28448 5072 28500 5092
rect 28500 5072 28502 5092
rect 29182 10104 29238 10160
rect 29090 9152 29146 9208
rect 28630 7248 28686 7304
rect 29366 8336 29422 8392
rect 29550 8472 29606 8528
rect 29274 7520 29330 7576
rect 28998 6296 29054 6352
rect 28630 6024 28686 6080
rect 27622 4922 27678 4924
rect 27702 4922 27758 4924
rect 27782 4922 27838 4924
rect 27862 4922 27918 4924
rect 27622 4870 27648 4922
rect 27648 4870 27678 4922
rect 27702 4870 27712 4922
rect 27712 4870 27758 4922
rect 27782 4870 27828 4922
rect 27828 4870 27838 4922
rect 27862 4870 27892 4922
rect 27892 4870 27918 4922
rect 27622 4868 27678 4870
rect 27702 4868 27758 4870
rect 27782 4868 27838 4870
rect 27862 4868 27918 4870
rect 26606 3712 26662 3768
rect 27622 3834 27678 3836
rect 27702 3834 27758 3836
rect 27782 3834 27838 3836
rect 27862 3834 27918 3836
rect 27622 3782 27648 3834
rect 27648 3782 27678 3834
rect 27702 3782 27712 3834
rect 27712 3782 27758 3834
rect 27782 3782 27828 3834
rect 27828 3782 27838 3834
rect 27862 3782 27892 3834
rect 27892 3782 27918 3834
rect 27622 3780 27678 3782
rect 27702 3780 27758 3782
rect 27782 3780 27838 3782
rect 27862 3780 27918 3782
rect 28998 5752 29054 5808
rect 30102 12824 30158 12880
rect 30654 12844 30710 12880
rect 30654 12824 30656 12844
rect 30656 12824 30708 12844
rect 30708 12824 30710 12844
rect 29918 12008 29974 12064
rect 30562 11872 30618 11928
rect 30194 8200 30250 8256
rect 30378 8200 30434 8256
rect 30378 7248 30434 7304
rect 30378 6704 30434 6760
rect 29734 6296 29790 6352
rect 29734 5480 29790 5536
rect 30470 6432 30526 6488
rect 30470 5752 30526 5808
rect 30930 9172 30986 9208
rect 30930 9152 30932 9172
rect 30932 9152 30984 9172
rect 30984 9152 30986 9172
rect 30654 8472 30710 8528
rect 30562 5072 30618 5128
rect 30378 4936 30434 4992
rect 30930 4800 30986 4856
rect 30470 4664 30526 4720
rect 30562 3984 30618 4040
rect 31666 12280 31722 12336
rect 31298 12144 31354 12200
rect 31758 12008 31814 12064
rect 32310 11328 32366 11384
rect 32678 10920 32734 10976
rect 32126 10648 32182 10704
rect 32954 10648 33010 10704
rect 31666 9832 31722 9888
rect 32126 9560 32182 9616
rect 32310 9324 32312 9344
rect 32312 9324 32364 9344
rect 32364 9324 32366 9344
rect 32310 9288 32366 9324
rect 32770 9152 32826 9208
rect 31758 7248 31814 7304
rect 32862 5888 32918 5944
rect 32862 4664 32918 4720
rect 33046 7384 33102 7440
rect 33230 7248 33286 7304
rect 33046 5888 33102 5944
rect 33230 5072 33286 5128
rect 33506 10648 33562 10704
rect 35806 15408 35862 15464
rect 34518 15000 34574 15056
rect 34702 14592 34758 14648
rect 34610 13812 34612 13832
rect 34612 13812 34664 13832
rect 34664 13812 34666 13832
rect 34610 13776 34666 13812
rect 34794 14184 34850 14240
rect 34794 13368 34850 13424
rect 34289 13082 34345 13084
rect 34369 13082 34425 13084
rect 34449 13082 34505 13084
rect 34529 13082 34585 13084
rect 34289 13030 34315 13082
rect 34315 13030 34345 13082
rect 34369 13030 34379 13082
rect 34379 13030 34425 13082
rect 34449 13030 34495 13082
rect 34495 13030 34505 13082
rect 34529 13030 34559 13082
rect 34559 13030 34585 13082
rect 34289 13028 34345 13030
rect 34369 13028 34425 13030
rect 34449 13028 34505 13030
rect 34529 13028 34585 13030
rect 34058 12316 34060 12336
rect 34060 12316 34112 12336
rect 34112 12316 34114 12336
rect 34058 12280 34114 12316
rect 33690 12144 33746 12200
rect 34610 12552 34666 12608
rect 34242 12144 34298 12200
rect 34289 11994 34345 11996
rect 34369 11994 34425 11996
rect 34449 11994 34505 11996
rect 34529 11994 34585 11996
rect 34289 11942 34315 11994
rect 34315 11942 34345 11994
rect 34369 11942 34379 11994
rect 34379 11942 34425 11994
rect 34449 11942 34495 11994
rect 34495 11942 34505 11994
rect 34529 11942 34559 11994
rect 34559 11942 34585 11994
rect 34289 11940 34345 11942
rect 34369 11940 34425 11942
rect 34449 11940 34505 11942
rect 34529 11940 34585 11942
rect 34794 11600 34850 11656
rect 33690 11464 33746 11520
rect 34289 10906 34345 10908
rect 34369 10906 34425 10908
rect 34449 10906 34505 10908
rect 34529 10906 34585 10908
rect 34289 10854 34315 10906
rect 34315 10854 34345 10906
rect 34369 10854 34379 10906
rect 34379 10854 34425 10906
rect 34449 10854 34495 10906
rect 34495 10854 34505 10906
rect 34529 10854 34559 10906
rect 34559 10854 34585 10906
rect 34289 10852 34345 10854
rect 34369 10852 34425 10854
rect 34449 10852 34505 10854
rect 34529 10852 34585 10854
rect 34334 10412 34336 10432
rect 34336 10412 34388 10432
rect 34388 10412 34390 10432
rect 34334 10376 34390 10412
rect 34289 9818 34345 9820
rect 34369 9818 34425 9820
rect 34449 9818 34505 9820
rect 34529 9818 34585 9820
rect 34289 9766 34315 9818
rect 34315 9766 34345 9818
rect 34369 9766 34379 9818
rect 34379 9766 34425 9818
rect 34449 9766 34495 9818
rect 34495 9766 34505 9818
rect 34529 9766 34559 9818
rect 34559 9766 34585 9818
rect 34289 9764 34345 9766
rect 34369 9764 34425 9766
rect 34449 9764 34505 9766
rect 34529 9764 34585 9766
rect 33690 9424 33746 9480
rect 33414 5752 33470 5808
rect 33414 5616 33470 5672
rect 33690 8064 33746 8120
rect 34702 9152 34758 9208
rect 34610 9016 34666 9072
rect 34289 8730 34345 8732
rect 34369 8730 34425 8732
rect 34449 8730 34505 8732
rect 34529 8730 34585 8732
rect 34289 8678 34315 8730
rect 34315 8678 34345 8730
rect 34369 8678 34379 8730
rect 34379 8678 34425 8730
rect 34449 8678 34495 8730
rect 34495 8678 34505 8730
rect 34529 8678 34559 8730
rect 34559 8678 34585 8730
rect 34289 8676 34345 8678
rect 34369 8676 34425 8678
rect 34449 8676 34505 8678
rect 34529 8676 34585 8678
rect 33966 8064 34022 8120
rect 33966 7792 34022 7848
rect 33690 7248 33746 7304
rect 33506 5344 33562 5400
rect 33690 4972 33692 4992
rect 33692 4972 33744 4992
rect 33744 4972 33746 4992
rect 33690 4936 33746 4972
rect 33322 4664 33378 4720
rect 34289 7642 34345 7644
rect 34369 7642 34425 7644
rect 34449 7642 34505 7644
rect 34529 7642 34585 7644
rect 34289 7590 34315 7642
rect 34315 7590 34345 7642
rect 34369 7590 34379 7642
rect 34379 7590 34425 7642
rect 34449 7590 34495 7642
rect 34495 7590 34505 7642
rect 34529 7590 34559 7642
rect 34559 7590 34585 7642
rect 34289 7588 34345 7590
rect 34369 7588 34425 7590
rect 34449 7588 34505 7590
rect 34529 7588 34585 7590
rect 34289 6554 34345 6556
rect 34369 6554 34425 6556
rect 34449 6554 34505 6556
rect 34529 6554 34585 6556
rect 34289 6502 34315 6554
rect 34315 6502 34345 6554
rect 34369 6502 34379 6554
rect 34379 6502 34425 6554
rect 34449 6502 34495 6554
rect 34495 6502 34505 6554
rect 34529 6502 34559 6554
rect 34559 6502 34585 6554
rect 34289 6500 34345 6502
rect 34369 6500 34425 6502
rect 34449 6500 34505 6502
rect 34529 6500 34585 6502
rect 34886 8200 34942 8256
rect 34978 8064 35034 8120
rect 35898 12960 35954 13016
rect 35622 12144 35678 12200
rect 35162 10784 35218 10840
rect 35438 10240 35494 10296
rect 35714 10376 35770 10432
rect 34794 7656 34850 7712
rect 35622 10104 35678 10160
rect 35622 9696 35678 9752
rect 34886 6876 34888 6896
rect 34888 6876 34940 6896
rect 34940 6876 34942 6896
rect 34886 6840 34942 6876
rect 35254 7384 35310 7440
rect 35070 6316 35126 6352
rect 35070 6296 35072 6316
rect 35072 6296 35124 6316
rect 35124 6296 35126 6316
rect 34978 5888 35034 5944
rect 34289 5466 34345 5468
rect 34369 5466 34425 5468
rect 34449 5466 34505 5468
rect 34529 5466 34585 5468
rect 34289 5414 34315 5466
rect 34315 5414 34345 5466
rect 34369 5414 34379 5466
rect 34379 5414 34425 5466
rect 34449 5414 34495 5466
rect 34495 5414 34505 5466
rect 34529 5414 34559 5466
rect 34559 5414 34585 5466
rect 34289 5412 34345 5414
rect 34369 5412 34425 5414
rect 34449 5412 34505 5414
rect 34529 5412 34585 5414
rect 34794 5208 34850 5264
rect 34610 4664 34666 4720
rect 33782 4528 33838 4584
rect 34289 4378 34345 4380
rect 34369 4378 34425 4380
rect 34449 4378 34505 4380
rect 34529 4378 34585 4380
rect 34289 4326 34315 4378
rect 34315 4326 34345 4378
rect 34369 4326 34379 4378
rect 34379 4326 34425 4378
rect 34449 4326 34495 4378
rect 34495 4326 34505 4378
rect 34529 4326 34559 4378
rect 34559 4326 34585 4378
rect 34289 4324 34345 4326
rect 34369 4324 34425 4326
rect 34449 4324 34505 4326
rect 34529 4324 34585 4326
rect 31206 3712 31262 3768
rect 29642 3576 29698 3632
rect 34289 3290 34345 3292
rect 34369 3290 34425 3292
rect 34449 3290 34505 3292
rect 34529 3290 34585 3292
rect 34289 3238 34315 3290
rect 34315 3238 34345 3290
rect 34369 3238 34379 3290
rect 34379 3238 34425 3290
rect 34449 3238 34495 3290
rect 34495 3238 34505 3290
rect 34529 3238 34559 3290
rect 34559 3238 34585 3290
rect 34289 3236 34345 3238
rect 34369 3236 34425 3238
rect 34449 3236 34505 3238
rect 34529 3236 34585 3238
rect 27342 2896 27398 2952
rect 27622 2746 27678 2748
rect 27702 2746 27758 2748
rect 27782 2746 27838 2748
rect 27862 2746 27918 2748
rect 27622 2694 27648 2746
rect 27648 2694 27678 2746
rect 27702 2694 27712 2746
rect 27712 2694 27758 2746
rect 27782 2694 27828 2746
rect 27828 2694 27838 2746
rect 27862 2694 27892 2746
rect 27892 2694 27918 2746
rect 27622 2692 27678 2694
rect 27702 2692 27758 2694
rect 27782 2692 27838 2694
rect 27862 2692 27918 2694
rect 34289 2202 34345 2204
rect 34369 2202 34425 2204
rect 34449 2202 34505 2204
rect 34529 2202 34585 2204
rect 34289 2150 34315 2202
rect 34315 2150 34345 2202
rect 34369 2150 34379 2202
rect 34379 2150 34425 2202
rect 34449 2150 34495 2202
rect 34495 2150 34505 2202
rect 34529 2150 34559 2202
rect 34559 2150 34585 2202
rect 34289 2148 34345 2150
rect 34369 2148 34425 2150
rect 34449 2148 34505 2150
rect 34529 2148 34585 2150
rect 25134 1672 25190 1728
rect 34610 856 34666 912
rect 2686 176 2742 232
rect 35438 4120 35494 4176
rect 36542 12824 36598 12880
rect 36174 12280 36230 12336
rect 36082 12008 36138 12064
rect 35806 9016 35862 9072
rect 35806 7928 35862 7984
rect 35714 7384 35770 7440
rect 35714 6568 35770 6624
rect 35622 4120 35678 4176
rect 35990 7656 36046 7712
rect 36726 11736 36782 11792
rect 36358 8472 36414 8528
rect 36542 11464 36598 11520
rect 36818 11056 36874 11112
rect 36726 10512 36782 10568
rect 36450 8372 36452 8392
rect 36452 8372 36504 8392
rect 36504 8372 36506 8392
rect 36450 8336 36506 8372
rect 36266 7248 36322 7304
rect 38658 11056 38714 11112
rect 37186 10920 37242 10976
rect 37554 10784 37610 10840
rect 36910 10648 36966 10704
rect 36910 8200 36966 8256
rect 35898 6024 35954 6080
rect 35806 5752 35862 5808
rect 36174 6840 36230 6896
rect 36082 6432 36138 6488
rect 35990 5616 36046 5672
rect 35714 3984 35770 4040
rect 37002 6976 37058 7032
rect 36634 5344 36690 5400
rect 35806 2896 35862 2952
rect 35622 2080 35678 2136
rect 35622 1400 35678 1456
rect 35346 1264 35402 1320
rect 34794 176 34850 232
rect 35162 448 35218 504
<< metal3 >>
rect 0 15874 480 15904
rect 3049 15874 3115 15877
rect 0 15872 3115 15874
rect 0 15816 3054 15872
rect 3110 15816 3115 15872
rect 0 15814 3115 15816
rect 0 15784 480 15814
rect 3049 15811 3115 15814
rect 36721 15874 36787 15877
rect 39520 15874 40000 15904
rect 36721 15872 40000 15874
rect 36721 15816 36726 15872
rect 36782 15816 40000 15872
rect 36721 15814 40000 15816
rect 36721 15811 36787 15814
rect 39520 15784 40000 15814
rect 0 15466 480 15496
rect 3417 15466 3483 15469
rect 0 15464 3483 15466
rect 0 15408 3422 15464
rect 3478 15408 3483 15464
rect 0 15406 3483 15408
rect 0 15376 480 15406
rect 3417 15403 3483 15406
rect 35801 15466 35867 15469
rect 39520 15466 40000 15496
rect 35801 15464 40000 15466
rect 35801 15408 35806 15464
rect 35862 15408 40000 15464
rect 35801 15406 40000 15408
rect 35801 15403 35867 15406
rect 39520 15376 40000 15406
rect 0 15058 480 15088
rect 3325 15058 3391 15061
rect 0 15056 3391 15058
rect 0 15000 3330 15056
rect 3386 15000 3391 15056
rect 0 14998 3391 15000
rect 0 14968 480 14998
rect 3325 14995 3391 14998
rect 34513 15058 34579 15061
rect 39520 15058 40000 15088
rect 34513 15056 40000 15058
rect 34513 15000 34518 15056
rect 34574 15000 40000 15056
rect 34513 14998 40000 15000
rect 34513 14995 34579 14998
rect 39520 14968 40000 14998
rect 0 14650 480 14680
rect 4429 14650 4495 14653
rect 0 14648 4495 14650
rect 0 14592 4434 14648
rect 4490 14592 4495 14648
rect 0 14590 4495 14592
rect 0 14560 480 14590
rect 4429 14587 4495 14590
rect 34697 14650 34763 14653
rect 39520 14650 40000 14680
rect 34697 14648 40000 14650
rect 34697 14592 34702 14648
rect 34758 14592 40000 14648
rect 34697 14590 40000 14592
rect 34697 14587 34763 14590
rect 39520 14560 40000 14590
rect 0 14242 480 14272
rect 4061 14242 4127 14245
rect 0 14240 4127 14242
rect 0 14184 4066 14240
rect 4122 14184 4127 14240
rect 0 14182 4127 14184
rect 0 14152 480 14182
rect 4061 14179 4127 14182
rect 34789 14242 34855 14245
rect 39520 14242 40000 14272
rect 34789 14240 40000 14242
rect 34789 14184 34794 14240
rect 34850 14184 40000 14240
rect 34789 14182 40000 14184
rect 34789 14179 34855 14182
rect 39520 14152 40000 14182
rect 0 13834 480 13864
rect 4337 13834 4403 13837
rect 0 13832 4403 13834
rect 0 13776 4342 13832
rect 4398 13776 4403 13832
rect 0 13774 4403 13776
rect 0 13744 480 13774
rect 4337 13771 4403 13774
rect 34605 13834 34671 13837
rect 39520 13834 40000 13864
rect 34605 13832 40000 13834
rect 34605 13776 34610 13832
rect 34666 13776 40000 13832
rect 34605 13774 40000 13776
rect 34605 13771 34671 13774
rect 39520 13744 40000 13774
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 27610 13632 27930 13633
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 13567 27930 13568
rect 0 13426 480 13456
rect 2773 13426 2839 13429
rect 0 13424 2839 13426
rect 0 13368 2778 13424
rect 2834 13368 2839 13424
rect 0 13366 2839 13368
rect 0 13336 480 13366
rect 2773 13363 2839 13366
rect 34789 13426 34855 13429
rect 39520 13426 40000 13456
rect 34789 13424 40000 13426
rect 34789 13368 34794 13424
rect 34850 13368 40000 13424
rect 34789 13366 40000 13368
rect 34789 13363 34855 13366
rect 39520 13336 40000 13366
rect 24025 13290 24091 13293
rect 27061 13290 27127 13293
rect 24025 13288 27127 13290
rect 24025 13232 24030 13288
rect 24086 13232 27066 13288
rect 27122 13232 27127 13288
rect 24025 13230 27127 13232
rect 24025 13227 24091 13230
rect 27061 13227 27127 13230
rect 7610 13088 7930 13089
rect 0 13018 480 13048
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7930 13088
rect 7610 13023 7930 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 34277 13088 34597 13089
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 13023 34597 13024
rect 4153 13018 4219 13021
rect 0 13016 4219 13018
rect 0 12960 4158 13016
rect 4214 12960 4219 13016
rect 0 12958 4219 12960
rect 0 12928 480 12958
rect 4153 12955 4219 12958
rect 24025 13018 24091 13021
rect 26233 13018 26299 13021
rect 24025 13016 26299 13018
rect 24025 12960 24030 13016
rect 24086 12960 26238 13016
rect 26294 12960 26299 13016
rect 24025 12958 26299 12960
rect 24025 12955 24091 12958
rect 26233 12955 26299 12958
rect 35893 13018 35959 13021
rect 39520 13018 40000 13048
rect 35893 13016 40000 13018
rect 35893 12960 35898 13016
rect 35954 12960 40000 13016
rect 35893 12958 40000 12960
rect 35893 12955 35959 12958
rect 39520 12928 40000 12958
rect 30097 12882 30163 12885
rect 30649 12882 30715 12885
rect 36537 12882 36603 12885
rect 30097 12880 36603 12882
rect 30097 12824 30102 12880
rect 30158 12824 30654 12880
rect 30710 12824 36542 12880
rect 36598 12824 36603 12880
rect 30097 12822 36603 12824
rect 30097 12819 30163 12822
rect 30649 12819 30715 12822
rect 36537 12819 36603 12822
rect 0 12610 480 12640
rect 4061 12610 4127 12613
rect 0 12608 4127 12610
rect 0 12552 4066 12608
rect 4122 12552 4127 12608
rect 0 12550 4127 12552
rect 0 12520 480 12550
rect 4061 12547 4127 12550
rect 34605 12610 34671 12613
rect 39520 12610 40000 12640
rect 34605 12608 40000 12610
rect 34605 12552 34610 12608
rect 34666 12552 40000 12608
rect 34605 12550 40000 12552
rect 34605 12547 34671 12550
rect 14277 12544 14597 12545
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 27610 12544 27930 12545
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 39520 12520 40000 12550
rect 27610 12479 27930 12480
rect 5165 12338 5231 12341
rect 23289 12338 23355 12341
rect 5165 12336 23355 12338
rect 5165 12280 5170 12336
rect 5226 12280 23294 12336
rect 23350 12280 23355 12336
rect 5165 12278 23355 12280
rect 5165 12275 5231 12278
rect 23289 12275 23355 12278
rect 25497 12338 25563 12341
rect 28349 12338 28415 12341
rect 31661 12338 31727 12341
rect 25497 12336 28274 12338
rect 25497 12280 25502 12336
rect 25558 12280 28274 12336
rect 25497 12278 28274 12280
rect 25497 12275 25563 12278
rect 0 12202 480 12232
rect 4245 12202 4311 12205
rect 0 12200 4311 12202
rect 0 12144 4250 12200
rect 4306 12144 4311 12200
rect 0 12142 4311 12144
rect 0 12112 480 12142
rect 4245 12139 4311 12142
rect 9581 12202 9647 12205
rect 22921 12202 22987 12205
rect 9581 12200 22987 12202
rect 9581 12144 9586 12200
rect 9642 12144 22926 12200
rect 22982 12144 22987 12200
rect 9581 12142 22987 12144
rect 9581 12139 9647 12142
rect 22921 12139 22987 12142
rect 27429 12202 27495 12205
rect 28214 12202 28274 12278
rect 28349 12336 31727 12338
rect 28349 12280 28354 12336
rect 28410 12280 31666 12336
rect 31722 12280 31727 12336
rect 28349 12278 31727 12280
rect 28349 12275 28415 12278
rect 31661 12275 31727 12278
rect 34053 12338 34119 12341
rect 36169 12338 36235 12341
rect 34053 12336 36235 12338
rect 34053 12280 34058 12336
rect 34114 12280 36174 12336
rect 36230 12280 36235 12336
rect 34053 12278 36235 12280
rect 34053 12275 34119 12278
rect 36169 12275 36235 12278
rect 28993 12202 29059 12205
rect 27429 12200 28090 12202
rect 27429 12144 27434 12200
rect 27490 12144 28090 12200
rect 27429 12142 28090 12144
rect 28214 12200 29059 12202
rect 28214 12144 28998 12200
rect 29054 12144 29059 12200
rect 28214 12142 29059 12144
rect 27429 12139 27495 12142
rect 16205 12066 16271 12069
rect 17953 12066 18019 12069
rect 16205 12064 18019 12066
rect 16205 12008 16210 12064
rect 16266 12008 17958 12064
rect 18014 12008 18019 12064
rect 16205 12006 18019 12008
rect 16205 12003 16271 12006
rect 17953 12003 18019 12006
rect 24393 12066 24459 12069
rect 27797 12066 27863 12069
rect 24393 12064 27863 12066
rect 24393 12008 24398 12064
rect 24454 12008 27802 12064
rect 27858 12008 27863 12064
rect 24393 12006 27863 12008
rect 28030 12066 28090 12142
rect 28993 12139 29059 12142
rect 31293 12202 31359 12205
rect 33685 12202 33751 12205
rect 31293 12200 33751 12202
rect 31293 12144 31298 12200
rect 31354 12144 33690 12200
rect 33746 12144 33751 12200
rect 31293 12142 33751 12144
rect 31293 12139 31359 12142
rect 33685 12139 33751 12142
rect 33910 12140 33916 12204
rect 33980 12202 33986 12204
rect 34237 12202 34303 12205
rect 35617 12202 35683 12205
rect 39520 12202 40000 12232
rect 33980 12200 35450 12202
rect 33980 12144 34242 12200
rect 34298 12144 35450 12200
rect 33980 12142 35450 12144
rect 33980 12140 33986 12142
rect 34237 12139 34303 12142
rect 29913 12066 29979 12069
rect 31753 12066 31819 12069
rect 28030 12064 31819 12066
rect 28030 12008 29918 12064
rect 29974 12008 31758 12064
rect 31814 12008 31819 12064
rect 28030 12006 31819 12008
rect 35390 12066 35450 12142
rect 35617 12200 40000 12202
rect 35617 12144 35622 12200
rect 35678 12144 40000 12200
rect 35617 12142 40000 12144
rect 35617 12139 35683 12142
rect 39520 12112 40000 12142
rect 36077 12066 36143 12069
rect 35390 12064 36143 12066
rect 35390 12008 36082 12064
rect 36138 12008 36143 12064
rect 35390 12006 36143 12008
rect 24393 12003 24459 12006
rect 27797 12003 27863 12006
rect 29913 12003 29979 12006
rect 31753 12003 31819 12006
rect 36077 12003 36143 12006
rect 7610 12000 7930 12001
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7930 12000
rect 7610 11935 7930 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 34277 12000 34597 12001
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 11935 34597 11936
rect 4521 11930 4587 11933
rect 4654 11930 4660 11932
rect 4521 11928 4660 11930
rect 4521 11872 4526 11928
rect 4582 11872 4660 11928
rect 4521 11870 4660 11872
rect 4521 11867 4587 11870
rect 4654 11868 4660 11870
rect 4724 11868 4730 11932
rect 24945 11930 25011 11933
rect 30557 11930 30623 11933
rect 24945 11928 30623 11930
rect 24945 11872 24950 11928
rect 25006 11872 30562 11928
rect 30618 11872 30623 11928
rect 24945 11870 30623 11872
rect 24945 11867 25011 11870
rect 30557 11867 30623 11870
rect 0 11794 480 11824
rect 1577 11794 1643 11797
rect 0 11792 1643 11794
rect 0 11736 1582 11792
rect 1638 11736 1643 11792
rect 0 11734 1643 11736
rect 0 11704 480 11734
rect 1577 11731 1643 11734
rect 6269 11794 6335 11797
rect 15193 11794 15259 11797
rect 6269 11792 15259 11794
rect 6269 11736 6274 11792
rect 6330 11736 15198 11792
rect 15254 11736 15259 11792
rect 6269 11734 15259 11736
rect 6269 11731 6335 11734
rect 15193 11731 15259 11734
rect 18597 11794 18663 11797
rect 26601 11794 26667 11797
rect 18597 11792 26667 11794
rect 18597 11736 18602 11792
rect 18658 11736 26606 11792
rect 26662 11736 26667 11792
rect 18597 11734 26667 11736
rect 18597 11731 18663 11734
rect 26601 11731 26667 11734
rect 36721 11794 36787 11797
rect 39520 11794 40000 11824
rect 36721 11792 40000 11794
rect 36721 11736 36726 11792
rect 36782 11736 40000 11792
rect 36721 11734 40000 11736
rect 36721 11731 36787 11734
rect 39520 11704 40000 11734
rect 3417 11658 3483 11661
rect 9121 11658 9187 11661
rect 3417 11656 9187 11658
rect 3417 11600 3422 11656
rect 3478 11600 9126 11656
rect 9182 11600 9187 11656
rect 3417 11598 9187 11600
rect 3417 11595 3483 11598
rect 9121 11595 9187 11598
rect 13537 11658 13603 11661
rect 16021 11658 16087 11661
rect 13537 11656 16087 11658
rect 13537 11600 13542 11656
rect 13598 11600 16026 11656
rect 16082 11600 16087 11656
rect 13537 11598 16087 11600
rect 13537 11595 13603 11598
rect 16021 11595 16087 11598
rect 16941 11658 17007 11661
rect 18689 11658 18755 11661
rect 16941 11656 18755 11658
rect 16941 11600 16946 11656
rect 17002 11600 18694 11656
rect 18750 11600 18755 11656
rect 16941 11598 18755 11600
rect 16941 11595 17007 11598
rect 18689 11595 18755 11598
rect 22921 11658 22987 11661
rect 34789 11658 34855 11661
rect 22921 11656 34855 11658
rect 22921 11600 22926 11656
rect 22982 11600 34794 11656
rect 34850 11600 34855 11656
rect 22921 11598 34855 11600
rect 22921 11595 22987 11598
rect 34789 11595 34855 11598
rect 4797 11522 4863 11525
rect 8937 11522 9003 11525
rect 4797 11520 9003 11522
rect 4797 11464 4802 11520
rect 4858 11464 8942 11520
rect 8998 11464 9003 11520
rect 4797 11462 9003 11464
rect 4797 11459 4863 11462
rect 8937 11459 9003 11462
rect 15377 11522 15443 11525
rect 24669 11522 24735 11525
rect 15377 11520 24735 11522
rect 15377 11464 15382 11520
rect 15438 11464 24674 11520
rect 24730 11464 24735 11520
rect 15377 11462 24735 11464
rect 15377 11459 15443 11462
rect 24669 11459 24735 11462
rect 33685 11522 33751 11525
rect 36537 11522 36603 11525
rect 33685 11520 36603 11522
rect 33685 11464 33690 11520
rect 33746 11464 36542 11520
rect 36598 11464 36603 11520
rect 33685 11462 36603 11464
rect 33685 11459 33751 11462
rect 36537 11459 36603 11462
rect 14277 11456 14597 11457
rect 0 11386 480 11416
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 27610 11456 27930 11457
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 11391 27930 11392
rect 5717 11386 5783 11389
rect 0 11384 5783 11386
rect 0 11328 5722 11384
rect 5778 11328 5783 11384
rect 0 11326 5783 11328
rect 0 11296 480 11326
rect 5717 11323 5783 11326
rect 21449 11386 21515 11389
rect 25129 11386 25195 11389
rect 21449 11384 25195 11386
rect 21449 11328 21454 11384
rect 21510 11328 25134 11384
rect 25190 11328 25195 11384
rect 21449 11326 25195 11328
rect 21449 11323 21515 11326
rect 25129 11323 25195 11326
rect 32305 11386 32371 11389
rect 39520 11386 40000 11416
rect 32305 11384 40000 11386
rect 32305 11328 32310 11384
rect 32366 11328 40000 11384
rect 32305 11326 40000 11328
rect 32305 11323 32371 11326
rect 39520 11296 40000 11326
rect 2313 11250 2379 11253
rect 5901 11250 5967 11253
rect 15377 11250 15443 11253
rect 2313 11248 5967 11250
rect 2313 11192 2318 11248
rect 2374 11192 5906 11248
rect 5962 11192 5967 11248
rect 2313 11190 5967 11192
rect 2313 11187 2379 11190
rect 5901 11187 5967 11190
rect 6134 11248 15443 11250
rect 6134 11192 15382 11248
rect 15438 11192 15443 11248
rect 6134 11190 15443 11192
rect 1853 11114 1919 11117
rect 3693 11114 3759 11117
rect 1853 11112 3759 11114
rect 1853 11056 1858 11112
rect 1914 11056 3698 11112
rect 3754 11056 3759 11112
rect 1853 11054 3759 11056
rect 1853 11051 1919 11054
rect 3693 11051 3759 11054
rect 4889 11114 4955 11117
rect 6134 11114 6194 11190
rect 15377 11187 15443 11190
rect 19977 11250 20043 11253
rect 26049 11250 26115 11253
rect 19977 11248 26115 11250
rect 19977 11192 19982 11248
rect 20038 11192 26054 11248
rect 26110 11192 26115 11248
rect 19977 11190 26115 11192
rect 19977 11187 20043 11190
rect 26049 11187 26115 11190
rect 4889 11112 6194 11114
rect 4889 11056 4894 11112
rect 4950 11056 6194 11112
rect 4889 11054 6194 11056
rect 9765 11114 9831 11117
rect 12801 11114 12867 11117
rect 9765 11112 12867 11114
rect 9765 11056 9770 11112
rect 9826 11056 12806 11112
rect 12862 11056 12867 11112
rect 9765 11054 12867 11056
rect 4889 11051 4955 11054
rect 9765 11051 9831 11054
rect 12801 11051 12867 11054
rect 25681 11114 25747 11117
rect 27889 11114 27955 11117
rect 25681 11112 27955 11114
rect 25681 11056 25686 11112
rect 25742 11056 27894 11112
rect 27950 11056 27955 11112
rect 25681 11054 27955 11056
rect 25681 11051 25747 11054
rect 27889 11051 27955 11054
rect 36813 11114 36879 11117
rect 38653 11114 38719 11117
rect 36813 11112 38719 11114
rect 36813 11056 36818 11112
rect 36874 11056 38658 11112
rect 38714 11056 38719 11112
rect 36813 11054 38719 11056
rect 36813 11051 36879 11054
rect 38653 11051 38719 11054
rect 0 10978 480 11008
rect 3969 10978 4035 10981
rect 0 10976 4035 10978
rect 0 10920 3974 10976
rect 4030 10920 4035 10976
rect 0 10918 4035 10920
rect 0 10888 480 10918
rect 3969 10915 4035 10918
rect 12249 10978 12315 10981
rect 18597 10978 18663 10981
rect 12249 10976 18663 10978
rect 12249 10920 12254 10976
rect 12310 10920 18602 10976
rect 18658 10920 18663 10976
rect 12249 10918 18663 10920
rect 12249 10915 12315 10918
rect 18597 10915 18663 10918
rect 26785 10978 26851 10981
rect 32673 10978 32739 10981
rect 26785 10976 32739 10978
rect 26785 10920 26790 10976
rect 26846 10920 32678 10976
rect 32734 10920 32739 10976
rect 26785 10918 32739 10920
rect 26785 10915 26851 10918
rect 32673 10915 32739 10918
rect 37181 10978 37247 10981
rect 39520 10978 40000 11008
rect 37181 10976 40000 10978
rect 37181 10920 37186 10976
rect 37242 10920 40000 10976
rect 37181 10918 40000 10920
rect 37181 10915 37247 10918
rect 7610 10912 7930 10913
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7930 10912
rect 7610 10847 7930 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 34277 10912 34597 10913
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 39520 10888 40000 10918
rect 34277 10847 34597 10848
rect 8109 10842 8175 10845
rect 22185 10842 22251 10845
rect 35157 10842 35223 10845
rect 37549 10842 37615 10845
rect 8109 10840 17234 10842
rect 8109 10784 8114 10840
rect 8170 10784 17234 10840
rect 8109 10782 17234 10784
rect 8109 10779 8175 10782
rect 8017 10706 8083 10709
rect 10225 10706 10291 10709
rect 17174 10706 17234 10782
rect 22185 10840 32874 10842
rect 22185 10784 22190 10840
rect 22246 10784 32874 10840
rect 22185 10782 32874 10784
rect 22185 10779 22251 10782
rect 24945 10706 25011 10709
rect 8017 10704 17050 10706
rect 8017 10648 8022 10704
rect 8078 10648 10230 10704
rect 10286 10648 17050 10704
rect 8017 10646 17050 10648
rect 17174 10704 25011 10706
rect 17174 10648 24950 10704
rect 25006 10648 25011 10704
rect 17174 10646 25011 10648
rect 8017 10643 8083 10646
rect 10225 10643 10291 10646
rect 0 10570 480 10600
rect 4061 10570 4127 10573
rect 8109 10570 8175 10573
rect 0 10568 4127 10570
rect 0 10512 4066 10568
rect 4122 10512 4127 10568
rect 0 10510 4127 10512
rect 0 10480 480 10510
rect 4061 10507 4127 10510
rect 4294 10568 8175 10570
rect 4294 10512 8114 10568
rect 8170 10512 8175 10568
rect 4294 10510 8175 10512
rect 3693 10434 3759 10437
rect 4294 10434 4354 10510
rect 8109 10507 8175 10510
rect 12065 10570 12131 10573
rect 16990 10570 17050 10646
rect 24945 10643 25011 10646
rect 26877 10706 26943 10709
rect 32121 10706 32187 10709
rect 26877 10704 32187 10706
rect 26877 10648 26882 10704
rect 26938 10648 32126 10704
rect 32182 10648 32187 10704
rect 26877 10646 32187 10648
rect 26877 10643 26943 10646
rect 32121 10643 32187 10646
rect 20805 10570 20871 10573
rect 22185 10570 22251 10573
rect 12065 10568 16866 10570
rect 12065 10512 12070 10568
rect 12126 10512 16866 10568
rect 12065 10510 16866 10512
rect 16990 10568 22251 10570
rect 16990 10512 20810 10568
rect 20866 10512 22190 10568
rect 22246 10512 22251 10568
rect 16990 10510 22251 10512
rect 12065 10507 12131 10510
rect 3693 10432 4354 10434
rect 3693 10376 3698 10432
rect 3754 10376 4354 10432
rect 3693 10374 4354 10376
rect 5441 10434 5507 10437
rect 8293 10434 8359 10437
rect 5441 10432 8359 10434
rect 5441 10376 5446 10432
rect 5502 10376 8298 10432
rect 8354 10376 8359 10432
rect 5441 10374 8359 10376
rect 16806 10434 16866 10510
rect 20805 10507 20871 10510
rect 22185 10507 22251 10510
rect 22461 10570 22527 10573
rect 22461 10568 32690 10570
rect 22461 10512 22466 10568
rect 22522 10512 32690 10568
rect 22461 10510 32690 10512
rect 22461 10507 22527 10510
rect 19057 10434 19123 10437
rect 16806 10432 19123 10434
rect 16806 10376 19062 10432
rect 19118 10376 19123 10432
rect 16806 10374 19123 10376
rect 3693 10371 3759 10374
rect 5441 10371 5507 10374
rect 8293 10371 8359 10374
rect 19057 10371 19123 10374
rect 20621 10434 20687 10437
rect 22277 10434 22343 10437
rect 20621 10432 22343 10434
rect 20621 10376 20626 10432
rect 20682 10376 22282 10432
rect 22338 10376 22343 10432
rect 20621 10374 22343 10376
rect 20621 10371 20687 10374
rect 22277 10371 22343 10374
rect 14277 10368 14597 10369
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 27610 10368 27930 10369
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 10303 27930 10304
rect 2497 10298 2563 10301
rect 4613 10298 4679 10301
rect 2497 10296 4679 10298
rect 2497 10240 2502 10296
rect 2558 10240 4618 10296
rect 4674 10240 4679 10296
rect 2497 10238 4679 10240
rect 2497 10235 2563 10238
rect 4613 10235 4679 10238
rect 6177 10298 6243 10301
rect 10133 10298 10199 10301
rect 6177 10296 10199 10298
rect 6177 10240 6182 10296
rect 6238 10240 10138 10296
rect 10194 10240 10199 10296
rect 6177 10238 10199 10240
rect 6177 10235 6243 10238
rect 10133 10235 10199 10238
rect 19425 10298 19491 10301
rect 26877 10298 26943 10301
rect 19425 10296 26943 10298
rect 19425 10240 19430 10296
rect 19486 10240 26882 10296
rect 26938 10240 26943 10296
rect 19425 10238 26943 10240
rect 32630 10298 32690 10510
rect 32814 10434 32874 10782
rect 35157 10840 37615 10842
rect 35157 10784 35162 10840
rect 35218 10784 37554 10840
rect 37610 10784 37615 10840
rect 35157 10782 37615 10784
rect 35157 10779 35223 10782
rect 37549 10779 37615 10782
rect 32949 10706 33015 10709
rect 33501 10706 33567 10709
rect 36905 10706 36971 10709
rect 32949 10704 36971 10706
rect 32949 10648 32954 10704
rect 33010 10648 33506 10704
rect 33562 10648 36910 10704
rect 36966 10648 36971 10704
rect 32949 10646 36971 10648
rect 32949 10643 33015 10646
rect 33501 10643 33567 10646
rect 36905 10643 36971 10646
rect 36721 10570 36787 10573
rect 39520 10570 40000 10600
rect 36721 10568 40000 10570
rect 36721 10512 36726 10568
rect 36782 10512 40000 10568
rect 36721 10510 40000 10512
rect 36721 10507 36787 10510
rect 39520 10480 40000 10510
rect 34329 10434 34395 10437
rect 35709 10434 35775 10437
rect 32814 10432 35775 10434
rect 32814 10376 34334 10432
rect 34390 10376 35714 10432
rect 35770 10376 35775 10432
rect 32814 10374 35775 10376
rect 34329 10371 34395 10374
rect 35709 10371 35775 10374
rect 35433 10298 35499 10301
rect 32630 10296 35499 10298
rect 32630 10240 35438 10296
rect 35494 10240 35499 10296
rect 32630 10238 35499 10240
rect 19425 10235 19491 10238
rect 26877 10235 26943 10238
rect 35433 10235 35499 10238
rect 0 10162 480 10192
rect 1393 10162 1459 10165
rect 0 10160 1459 10162
rect 0 10104 1398 10160
rect 1454 10104 1459 10160
rect 0 10102 1459 10104
rect 0 10072 480 10102
rect 1393 10099 1459 10102
rect 4705 10162 4771 10165
rect 14181 10162 14247 10165
rect 29177 10162 29243 10165
rect 4705 10160 29243 10162
rect 4705 10104 4710 10160
rect 4766 10104 14186 10160
rect 14242 10104 29182 10160
rect 29238 10104 29243 10160
rect 4705 10102 29243 10104
rect 4705 10099 4771 10102
rect 14181 10099 14247 10102
rect 29177 10099 29243 10102
rect 35617 10162 35683 10165
rect 39520 10162 40000 10192
rect 35617 10160 40000 10162
rect 35617 10104 35622 10160
rect 35678 10104 40000 10160
rect 35617 10102 40000 10104
rect 35617 10099 35683 10102
rect 39520 10072 40000 10102
rect 2405 10026 2471 10029
rect 4981 10026 5047 10029
rect 2405 10024 5047 10026
rect 2405 9968 2410 10024
rect 2466 9968 4986 10024
rect 5042 9968 5047 10024
rect 2405 9966 5047 9968
rect 2405 9963 2471 9966
rect 4981 9963 5047 9966
rect 7465 10026 7531 10029
rect 11973 10026 12039 10029
rect 7465 10024 12039 10026
rect 7465 9968 7470 10024
rect 7526 9968 11978 10024
rect 12034 9968 12039 10024
rect 7465 9966 12039 9968
rect 7465 9963 7531 9966
rect 11973 9963 12039 9966
rect 18781 10026 18847 10029
rect 23473 10026 23539 10029
rect 18781 10024 23539 10026
rect 18781 9968 18786 10024
rect 18842 9968 23478 10024
rect 23534 9968 23539 10024
rect 18781 9966 23539 9968
rect 18781 9963 18847 9966
rect 23473 9963 23539 9966
rect 9857 9890 9923 9893
rect 20161 9890 20227 9893
rect 31661 9890 31727 9893
rect 9857 9888 20227 9890
rect 9857 9832 9862 9888
rect 9918 9832 20166 9888
rect 20222 9832 20227 9888
rect 9857 9830 20227 9832
rect 9857 9827 9923 9830
rect 20161 9827 20227 9830
rect 24534 9888 31727 9890
rect 24534 9832 31666 9888
rect 31722 9832 31727 9888
rect 24534 9830 31727 9832
rect 7610 9824 7930 9825
rect 0 9754 480 9784
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7930 9824
rect 7610 9759 7930 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 15193 9754 15259 9757
rect 24301 9754 24367 9757
rect 0 9694 1594 9754
rect 0 9664 480 9694
rect 1534 9618 1594 9694
rect 15193 9752 20730 9754
rect 15193 9696 15198 9752
rect 15254 9696 20730 9752
rect 15193 9694 20730 9696
rect 15193 9691 15259 9694
rect 1669 9618 1735 9621
rect 1534 9616 1735 9618
rect 1534 9560 1674 9616
rect 1730 9560 1735 9616
rect 1534 9558 1735 9560
rect 1669 9555 1735 9558
rect 4061 9618 4127 9621
rect 5533 9618 5599 9621
rect 4061 9616 5599 9618
rect 4061 9560 4066 9616
rect 4122 9560 5538 9616
rect 5594 9560 5599 9616
rect 4061 9558 5599 9560
rect 4061 9555 4127 9558
rect 5533 9555 5599 9558
rect 11421 9618 11487 9621
rect 13445 9618 13511 9621
rect 13813 9618 13879 9621
rect 11421 9616 13879 9618
rect 11421 9560 11426 9616
rect 11482 9560 13450 9616
rect 13506 9560 13818 9616
rect 13874 9560 13879 9616
rect 11421 9558 13879 9560
rect 11421 9555 11487 9558
rect 13445 9555 13511 9558
rect 13813 9555 13879 9558
rect 13997 9618 14063 9621
rect 20069 9618 20135 9621
rect 13997 9616 20135 9618
rect 13997 9560 14002 9616
rect 14058 9560 20074 9616
rect 20130 9560 20135 9616
rect 13997 9558 20135 9560
rect 20670 9618 20730 9694
rect 21406 9752 24367 9754
rect 21406 9696 24306 9752
rect 24362 9696 24367 9752
rect 21406 9694 24367 9696
rect 21406 9618 21466 9694
rect 24301 9691 24367 9694
rect 24534 9618 24594 9830
rect 31661 9827 31727 9830
rect 34277 9824 34597 9825
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 9759 34597 9760
rect 35617 9754 35683 9757
rect 39520 9754 40000 9784
rect 35617 9752 40000 9754
rect 35617 9696 35622 9752
rect 35678 9696 40000 9752
rect 35617 9694 40000 9696
rect 35617 9691 35683 9694
rect 39520 9664 40000 9694
rect 20670 9558 21466 9618
rect 24166 9558 24594 9618
rect 28165 9618 28231 9621
rect 32121 9618 32187 9621
rect 28165 9616 32187 9618
rect 28165 9560 28170 9616
rect 28226 9560 32126 9616
rect 32182 9560 32187 9616
rect 28165 9558 32187 9560
rect 13997 9555 14063 9558
rect 20069 9555 20135 9558
rect 11145 9482 11211 9485
rect 24025 9482 24091 9485
rect 24166 9482 24226 9558
rect 28165 9555 28231 9558
rect 32121 9555 32187 9558
rect 11145 9480 24226 9482
rect 11145 9424 11150 9480
rect 11206 9424 24030 9480
rect 24086 9424 24226 9480
rect 11145 9422 24226 9424
rect 24301 9482 24367 9485
rect 33685 9482 33751 9485
rect 24301 9480 33751 9482
rect 24301 9424 24306 9480
rect 24362 9424 33690 9480
rect 33746 9424 33751 9480
rect 24301 9422 33751 9424
rect 11145 9419 11211 9422
rect 24025 9419 24091 9422
rect 24301 9419 24367 9422
rect 33685 9419 33751 9422
rect 0 9346 480 9376
rect 5809 9346 5875 9349
rect 0 9344 5875 9346
rect 0 9288 5814 9344
rect 5870 9288 5875 9344
rect 0 9286 5875 9288
rect 0 9256 480 9286
rect 5809 9283 5875 9286
rect 7649 9346 7715 9349
rect 12249 9346 12315 9349
rect 7649 9344 12315 9346
rect 7649 9288 7654 9344
rect 7710 9288 12254 9344
rect 12310 9288 12315 9344
rect 7649 9286 12315 9288
rect 7649 9283 7715 9286
rect 12249 9283 12315 9286
rect 32305 9346 32371 9349
rect 39520 9346 40000 9376
rect 32305 9344 40000 9346
rect 32305 9288 32310 9344
rect 32366 9288 40000 9344
rect 32305 9286 40000 9288
rect 32305 9283 32371 9286
rect 14277 9280 14597 9281
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 27610 9280 27930 9281
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 39520 9256 40000 9286
rect 27610 9215 27930 9216
rect 4521 9210 4587 9213
rect 10593 9210 10659 9213
rect 12985 9210 13051 9213
rect 13997 9210 14063 9213
rect 4521 9208 10659 9210
rect 4521 9152 4526 9208
rect 4582 9152 10598 9208
rect 10654 9152 10659 9208
rect 4521 9150 10659 9152
rect 4521 9147 4587 9150
rect 10593 9147 10659 9150
rect 10734 9208 14063 9210
rect 10734 9152 12990 9208
rect 13046 9152 14002 9208
rect 14058 9152 14063 9208
rect 10734 9150 14063 9152
rect 6085 9074 6151 9077
rect 10734 9074 10794 9150
rect 12985 9147 13051 9150
rect 13997 9147 14063 9150
rect 18597 9210 18663 9213
rect 22921 9210 22987 9213
rect 18597 9208 22987 9210
rect 18597 9152 18602 9208
rect 18658 9152 22926 9208
rect 22982 9152 22987 9208
rect 18597 9150 22987 9152
rect 18597 9147 18663 9150
rect 22921 9147 22987 9150
rect 23841 9210 23907 9213
rect 27153 9210 27219 9213
rect 23841 9208 27219 9210
rect 23841 9152 23846 9208
rect 23902 9152 27158 9208
rect 27214 9152 27219 9208
rect 23841 9150 27219 9152
rect 23841 9147 23907 9150
rect 27153 9147 27219 9150
rect 29085 9210 29151 9213
rect 30925 9210 30991 9213
rect 29085 9208 30991 9210
rect 29085 9152 29090 9208
rect 29146 9152 30930 9208
rect 30986 9152 30991 9208
rect 29085 9150 30991 9152
rect 29085 9147 29151 9150
rect 30925 9147 30991 9150
rect 32765 9210 32831 9213
rect 34697 9210 34763 9213
rect 32765 9208 34763 9210
rect 32765 9152 32770 9208
rect 32826 9152 34702 9208
rect 34758 9152 34763 9208
rect 32765 9150 34763 9152
rect 32765 9147 32831 9150
rect 34697 9147 34763 9150
rect 6085 9072 10794 9074
rect 6085 9016 6090 9072
rect 6146 9016 10794 9072
rect 6085 9014 10794 9016
rect 11421 9074 11487 9077
rect 21265 9074 21331 9077
rect 11421 9072 21331 9074
rect 11421 9016 11426 9072
rect 11482 9016 21270 9072
rect 21326 9016 21331 9072
rect 11421 9014 21331 9016
rect 6085 9011 6151 9014
rect 11421 9011 11487 9014
rect 21265 9011 21331 9014
rect 22369 9074 22435 9077
rect 24945 9074 25011 9077
rect 27429 9074 27495 9077
rect 34605 9074 34671 9077
rect 22369 9072 34671 9074
rect 22369 9016 22374 9072
rect 22430 9016 24950 9072
rect 25006 9016 27434 9072
rect 27490 9016 34610 9072
rect 34666 9016 34671 9072
rect 22369 9014 34671 9016
rect 22369 9011 22435 9014
rect 24945 9011 25011 9014
rect 27429 9011 27495 9014
rect 34605 9011 34671 9014
rect 35801 9074 35867 9077
rect 35801 9072 37658 9074
rect 35801 9016 35806 9072
rect 35862 9016 37658 9072
rect 35801 9014 37658 9016
rect 35801 9011 35867 9014
rect 0 8938 480 8968
rect 4245 8938 4311 8941
rect 0 8936 4311 8938
rect 0 8880 4250 8936
rect 4306 8880 4311 8936
rect 0 8878 4311 8880
rect 0 8848 480 8878
rect 4245 8875 4311 8878
rect 5993 8938 6059 8941
rect 10961 8938 11027 8941
rect 12525 8938 12591 8941
rect 5993 8936 12591 8938
rect 5993 8880 5998 8936
rect 6054 8880 10966 8936
rect 11022 8880 12530 8936
rect 12586 8880 12591 8936
rect 5993 8878 12591 8880
rect 5993 8875 6059 8878
rect 10961 8875 11027 8878
rect 12525 8875 12591 8878
rect 12709 8938 12775 8941
rect 16665 8938 16731 8941
rect 12709 8936 16731 8938
rect 12709 8880 12714 8936
rect 12770 8880 16670 8936
rect 16726 8880 16731 8936
rect 12709 8878 16731 8880
rect 12709 8875 12775 8878
rect 16665 8875 16731 8878
rect 19057 8938 19123 8941
rect 23197 8938 23263 8941
rect 19057 8936 23263 8938
rect 19057 8880 19062 8936
rect 19118 8880 23202 8936
rect 23258 8880 23263 8936
rect 19057 8878 23263 8880
rect 37598 8938 37658 9014
rect 39520 8938 40000 8968
rect 37598 8878 40000 8938
rect 19057 8875 19123 8878
rect 23197 8875 23263 8878
rect 39520 8848 40000 8878
rect 10225 8802 10291 8805
rect 13813 8802 13879 8805
rect 10225 8800 13879 8802
rect 10225 8744 10230 8800
rect 10286 8744 13818 8800
rect 13874 8744 13879 8800
rect 10225 8742 13879 8744
rect 10225 8739 10291 8742
rect 13813 8739 13879 8742
rect 14273 8802 14339 8805
rect 19793 8802 19859 8805
rect 14273 8800 19859 8802
rect 14273 8744 14278 8800
rect 14334 8744 19798 8800
rect 19854 8744 19859 8800
rect 14273 8742 19859 8744
rect 14273 8739 14339 8742
rect 19793 8739 19859 8742
rect 7610 8736 7930 8737
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7930 8736
rect 7610 8671 7930 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 34277 8736 34597 8737
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 8671 34597 8672
rect 4613 8666 4679 8669
rect 7097 8666 7163 8669
rect 4613 8664 7163 8666
rect 4613 8608 4618 8664
rect 4674 8608 7102 8664
rect 7158 8608 7163 8664
rect 4613 8606 7163 8608
rect 4613 8603 4679 8606
rect 7097 8603 7163 8606
rect 8017 8666 8083 8669
rect 12893 8666 12959 8669
rect 8017 8664 17418 8666
rect 8017 8608 8022 8664
rect 8078 8608 12898 8664
rect 12954 8608 17418 8664
rect 8017 8606 17418 8608
rect 8017 8603 8083 8606
rect 12893 8603 12959 8606
rect 0 8530 480 8560
rect 4153 8530 4219 8533
rect 0 8528 4219 8530
rect 0 8472 4158 8528
rect 4214 8472 4219 8528
rect 0 8470 4219 8472
rect 0 8440 480 8470
rect 4153 8467 4219 8470
rect 6361 8530 6427 8533
rect 9949 8530 10015 8533
rect 6361 8528 10015 8530
rect 6361 8472 6366 8528
rect 6422 8472 9954 8528
rect 10010 8472 10015 8528
rect 6361 8470 10015 8472
rect 6361 8467 6427 8470
rect 9949 8467 10015 8470
rect 12525 8530 12591 8533
rect 14273 8530 14339 8533
rect 12525 8528 14339 8530
rect 12525 8472 12530 8528
rect 12586 8472 14278 8528
rect 14334 8472 14339 8528
rect 12525 8470 14339 8472
rect 12525 8467 12591 8470
rect 14273 8467 14339 8470
rect 14457 8530 14523 8533
rect 15377 8530 15443 8533
rect 17125 8530 17191 8533
rect 14457 8528 17191 8530
rect 14457 8472 14462 8528
rect 14518 8472 15382 8528
rect 15438 8472 17130 8528
rect 17186 8472 17191 8528
rect 14457 8470 17191 8472
rect 17358 8530 17418 8606
rect 21725 8530 21791 8533
rect 17358 8528 21791 8530
rect 17358 8472 21730 8528
rect 21786 8472 21791 8528
rect 17358 8470 21791 8472
rect 14457 8467 14523 8470
rect 15377 8467 15443 8470
rect 17125 8467 17191 8470
rect 21725 8467 21791 8470
rect 22001 8530 22067 8533
rect 26693 8530 26759 8533
rect 29545 8530 29611 8533
rect 30649 8530 30715 8533
rect 22001 8528 26618 8530
rect 22001 8472 22006 8528
rect 22062 8472 26618 8528
rect 22001 8470 26618 8472
rect 22001 8467 22067 8470
rect 5717 8394 5783 8397
rect 9765 8394 9831 8397
rect 5717 8392 9831 8394
rect 5717 8336 5722 8392
rect 5778 8336 9770 8392
rect 9826 8336 9831 8392
rect 5717 8334 9831 8336
rect 5717 8331 5783 8334
rect 9765 8331 9831 8334
rect 15653 8394 15719 8397
rect 18689 8394 18755 8397
rect 15653 8392 18755 8394
rect 15653 8336 15658 8392
rect 15714 8336 18694 8392
rect 18750 8336 18755 8392
rect 15653 8334 18755 8336
rect 15653 8331 15719 8334
rect 18689 8331 18755 8334
rect 21449 8394 21515 8397
rect 24209 8394 24275 8397
rect 21449 8392 24275 8394
rect 21449 8336 21454 8392
rect 21510 8336 24214 8392
rect 24270 8336 24275 8392
rect 21449 8334 24275 8336
rect 26558 8394 26618 8470
rect 26693 8528 30715 8530
rect 26693 8472 26698 8528
rect 26754 8472 29550 8528
rect 29606 8472 30654 8528
rect 30710 8472 30715 8528
rect 26693 8470 30715 8472
rect 26693 8467 26759 8470
rect 29545 8467 29611 8470
rect 30649 8467 30715 8470
rect 36353 8530 36419 8533
rect 39520 8530 40000 8560
rect 36353 8528 40000 8530
rect 36353 8472 36358 8528
rect 36414 8472 40000 8528
rect 36353 8470 40000 8472
rect 36353 8467 36419 8470
rect 39520 8440 40000 8470
rect 29361 8394 29427 8397
rect 36445 8394 36511 8397
rect 26558 8334 28090 8394
rect 21449 8331 21515 8334
rect 24209 8331 24275 8334
rect 0 8258 480 8288
rect 1577 8258 1643 8261
rect 0 8256 1643 8258
rect 0 8200 1582 8256
rect 1638 8200 1643 8256
rect 0 8198 1643 8200
rect 0 8168 480 8198
rect 1577 8195 1643 8198
rect 2957 8258 3023 8261
rect 11789 8258 11855 8261
rect 2957 8256 11855 8258
rect 2957 8200 2962 8256
rect 3018 8200 11794 8256
rect 11850 8200 11855 8256
rect 2957 8198 11855 8200
rect 2957 8195 3023 8198
rect 11789 8195 11855 8198
rect 17309 8258 17375 8261
rect 20897 8258 20963 8261
rect 17309 8256 20963 8258
rect 17309 8200 17314 8256
rect 17370 8200 20902 8256
rect 20958 8200 20963 8256
rect 17309 8198 20963 8200
rect 17309 8195 17375 8198
rect 20897 8195 20963 8198
rect 23381 8258 23447 8261
rect 27337 8258 27403 8261
rect 23381 8256 27403 8258
rect 23381 8200 23386 8256
rect 23442 8200 27342 8256
rect 27398 8200 27403 8256
rect 23381 8198 27403 8200
rect 23381 8195 23447 8198
rect 27337 8195 27403 8198
rect 14277 8192 14597 8193
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 27610 8192 27930 8193
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 8127 27930 8128
rect 7741 8122 7807 8125
rect 10409 8122 10475 8125
rect 23933 8122 23999 8125
rect 7741 8120 10475 8122
rect 7741 8064 7746 8120
rect 7802 8064 10414 8120
rect 10470 8064 10475 8120
rect 7741 8062 10475 8064
rect 7741 8059 7807 8062
rect 10409 8059 10475 8062
rect 17174 8120 23999 8122
rect 17174 8064 23938 8120
rect 23994 8064 23999 8120
rect 17174 8062 23999 8064
rect 7649 7986 7715 7989
rect 17174 7986 17234 8062
rect 23933 8059 23999 8062
rect 7649 7984 17234 7986
rect 7649 7928 7654 7984
rect 7710 7928 17234 7984
rect 7649 7926 17234 7928
rect 28030 7986 28090 8334
rect 29361 8392 36511 8394
rect 29361 8336 29366 8392
rect 29422 8336 36450 8392
rect 36506 8336 36511 8392
rect 29361 8334 36511 8336
rect 29361 8331 29427 8334
rect 36445 8331 36511 8334
rect 28441 8258 28507 8261
rect 30189 8258 30255 8261
rect 28441 8256 30255 8258
rect 28441 8200 28446 8256
rect 28502 8200 30194 8256
rect 30250 8200 30255 8256
rect 28441 8198 30255 8200
rect 28441 8195 28507 8198
rect 30189 8195 30255 8198
rect 30373 8258 30439 8261
rect 34881 8258 34947 8261
rect 30373 8256 34947 8258
rect 30373 8200 30378 8256
rect 30434 8200 34886 8256
rect 34942 8200 34947 8256
rect 30373 8198 34947 8200
rect 30373 8195 30439 8198
rect 34881 8195 34947 8198
rect 36905 8258 36971 8261
rect 39520 8258 40000 8288
rect 36905 8256 40000 8258
rect 36905 8200 36910 8256
rect 36966 8200 40000 8256
rect 36905 8198 40000 8200
rect 36905 8195 36971 8198
rect 39520 8168 40000 8198
rect 28349 8122 28415 8125
rect 33685 8122 33751 8125
rect 28349 8120 33751 8122
rect 28349 8064 28354 8120
rect 28410 8064 33690 8120
rect 33746 8064 33751 8120
rect 28349 8062 33751 8064
rect 28349 8059 28415 8062
rect 33685 8059 33751 8062
rect 33961 8122 34027 8125
rect 34973 8122 35039 8125
rect 33961 8120 35039 8122
rect 33961 8064 33966 8120
rect 34022 8064 34978 8120
rect 35034 8064 35039 8120
rect 33961 8062 35039 8064
rect 33961 8059 34027 8062
rect 34973 8059 35039 8062
rect 35801 7986 35867 7989
rect 28030 7984 35867 7986
rect 28030 7928 35806 7984
rect 35862 7928 35867 7984
rect 28030 7926 35867 7928
rect 7649 7923 7715 7926
rect 35801 7923 35867 7926
rect 0 7850 480 7880
rect 4889 7850 4955 7853
rect 0 7848 4955 7850
rect 0 7792 4894 7848
rect 4950 7792 4955 7848
rect 0 7790 4955 7792
rect 0 7760 480 7790
rect 4889 7787 4955 7790
rect 6177 7850 6243 7853
rect 11329 7850 11395 7853
rect 6177 7848 11395 7850
rect 6177 7792 6182 7848
rect 6238 7792 11334 7848
rect 11390 7792 11395 7848
rect 6177 7790 11395 7792
rect 6177 7787 6243 7790
rect 11329 7787 11395 7790
rect 16297 7850 16363 7853
rect 25221 7850 25287 7853
rect 16297 7848 25287 7850
rect 16297 7792 16302 7848
rect 16358 7792 25226 7848
rect 25282 7792 25287 7848
rect 16297 7790 25287 7792
rect 16297 7787 16363 7790
rect 25221 7787 25287 7790
rect 26877 7850 26943 7853
rect 33961 7850 34027 7853
rect 39520 7850 40000 7880
rect 26877 7848 34027 7850
rect 26877 7792 26882 7848
rect 26938 7792 33966 7848
rect 34022 7792 34027 7848
rect 26877 7790 34027 7792
rect 26877 7787 26943 7790
rect 33961 7787 34027 7790
rect 34102 7790 40000 7850
rect 10961 7714 11027 7717
rect 15653 7714 15719 7717
rect 17033 7714 17099 7717
rect 19333 7714 19399 7717
rect 10961 7712 16866 7714
rect 10961 7656 10966 7712
rect 11022 7656 15658 7712
rect 15714 7656 16866 7712
rect 10961 7654 16866 7656
rect 10961 7651 11027 7654
rect 15653 7651 15719 7654
rect 7610 7648 7930 7649
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7930 7648
rect 7610 7583 7930 7584
rect 2589 7578 2655 7581
rect 8201 7578 8267 7581
rect 15469 7578 15535 7581
rect 2589 7576 7482 7578
rect 2589 7520 2594 7576
rect 2650 7520 7482 7576
rect 2589 7518 7482 7520
rect 2589 7515 2655 7518
rect 0 7442 480 7472
rect 4797 7442 4863 7445
rect 0 7440 4863 7442
rect 0 7384 4802 7440
rect 4858 7384 4863 7440
rect 0 7382 4863 7384
rect 7422 7442 7482 7518
rect 8201 7576 15535 7578
rect 8201 7520 8206 7576
rect 8262 7520 15474 7576
rect 15530 7520 15535 7576
rect 8201 7518 15535 7520
rect 16806 7578 16866 7654
rect 17033 7712 19399 7714
rect 17033 7656 17038 7712
rect 17094 7656 19338 7712
rect 19394 7656 19399 7712
rect 17033 7654 19399 7656
rect 17033 7651 17099 7654
rect 19333 7651 19399 7654
rect 27061 7714 27127 7717
rect 34102 7714 34162 7790
rect 39520 7760 40000 7790
rect 27061 7712 34162 7714
rect 27061 7656 27066 7712
rect 27122 7656 34162 7712
rect 27061 7654 34162 7656
rect 34789 7714 34855 7717
rect 35985 7714 36051 7717
rect 34789 7712 36051 7714
rect 34789 7656 34794 7712
rect 34850 7656 35990 7712
rect 36046 7656 36051 7712
rect 34789 7654 36051 7656
rect 27061 7651 27127 7654
rect 34789 7651 34855 7654
rect 35985 7651 36051 7654
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 34277 7648 34597 7649
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 7583 34597 7584
rect 19425 7578 19491 7581
rect 16806 7576 19491 7578
rect 16806 7520 19430 7576
rect 19486 7520 19491 7576
rect 16806 7518 19491 7520
rect 8201 7515 8267 7518
rect 15469 7515 15535 7518
rect 19425 7515 19491 7518
rect 21633 7578 21699 7581
rect 29269 7578 29335 7581
rect 21633 7576 30666 7578
rect 21633 7520 21638 7576
rect 21694 7520 29274 7576
rect 29330 7520 30666 7576
rect 21633 7518 30666 7520
rect 21633 7515 21699 7518
rect 29269 7515 29335 7518
rect 16573 7442 16639 7445
rect 7422 7440 16639 7442
rect 7422 7384 16578 7440
rect 16634 7384 16639 7440
rect 7422 7382 16639 7384
rect 0 7352 480 7382
rect 4797 7379 4863 7382
rect 16573 7379 16639 7382
rect 19609 7442 19675 7445
rect 24209 7442 24275 7445
rect 25313 7442 25379 7445
rect 19609 7440 25379 7442
rect 19609 7384 19614 7440
rect 19670 7384 24214 7440
rect 24270 7384 25318 7440
rect 25374 7384 25379 7440
rect 19609 7382 25379 7384
rect 19609 7379 19675 7382
rect 24209 7379 24275 7382
rect 25313 7379 25379 7382
rect 5901 7306 5967 7309
rect 8937 7306 9003 7309
rect 5901 7304 9003 7306
rect 5901 7248 5906 7304
rect 5962 7248 8942 7304
rect 8998 7248 9003 7304
rect 5901 7246 9003 7248
rect 5901 7243 5967 7246
rect 8937 7243 9003 7246
rect 11789 7306 11855 7309
rect 14641 7306 14707 7309
rect 11789 7304 14707 7306
rect 11789 7248 11794 7304
rect 11850 7248 14646 7304
rect 14702 7248 14707 7304
rect 11789 7246 14707 7248
rect 11789 7243 11855 7246
rect 14641 7243 14707 7246
rect 16665 7306 16731 7309
rect 26877 7306 26943 7309
rect 28625 7306 28691 7309
rect 30373 7306 30439 7309
rect 16665 7304 26943 7306
rect 16665 7248 16670 7304
rect 16726 7248 26882 7304
rect 26938 7248 26943 7304
rect 16665 7246 26943 7248
rect 16665 7243 16731 7246
rect 26877 7243 26943 7246
rect 27478 7304 30439 7306
rect 27478 7248 28630 7304
rect 28686 7248 30378 7304
rect 30434 7248 30439 7304
rect 27478 7246 30439 7248
rect 30606 7306 30666 7518
rect 33041 7442 33107 7445
rect 35249 7442 35315 7445
rect 33041 7440 35315 7442
rect 33041 7384 33046 7440
rect 33102 7384 35254 7440
rect 35310 7384 35315 7440
rect 33041 7382 35315 7384
rect 33041 7379 33107 7382
rect 35249 7379 35315 7382
rect 35709 7442 35775 7445
rect 39520 7442 40000 7472
rect 35709 7440 40000 7442
rect 35709 7384 35714 7440
rect 35770 7384 40000 7440
rect 35709 7382 40000 7384
rect 35709 7379 35775 7382
rect 39520 7352 40000 7382
rect 31753 7306 31819 7309
rect 33225 7306 33291 7309
rect 30606 7304 33291 7306
rect 30606 7248 31758 7304
rect 31814 7248 33230 7304
rect 33286 7248 33291 7304
rect 30606 7246 33291 7248
rect 3233 7170 3299 7173
rect 10409 7170 10475 7173
rect 3233 7168 10475 7170
rect 3233 7112 3238 7168
rect 3294 7112 10414 7168
rect 10470 7112 10475 7168
rect 3233 7110 10475 7112
rect 3233 7107 3299 7110
rect 10409 7107 10475 7110
rect 25221 7170 25287 7173
rect 27478 7170 27538 7246
rect 28625 7243 28691 7246
rect 30373 7243 30439 7246
rect 31753 7243 31819 7246
rect 33225 7243 33291 7246
rect 33685 7306 33751 7309
rect 36261 7306 36327 7309
rect 33685 7304 36327 7306
rect 33685 7248 33690 7304
rect 33746 7248 36266 7304
rect 36322 7248 36327 7304
rect 33685 7246 36327 7248
rect 33685 7243 33751 7246
rect 36261 7243 36327 7246
rect 25221 7168 27538 7170
rect 25221 7112 25226 7168
rect 25282 7112 27538 7168
rect 25221 7110 27538 7112
rect 25221 7107 25287 7110
rect 14277 7104 14597 7105
rect 0 7034 480 7064
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 7039 14597 7040
rect 27610 7104 27930 7105
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 7039 27930 7040
rect 3509 7034 3575 7037
rect 0 7032 3575 7034
rect 0 6976 3514 7032
rect 3570 6976 3575 7032
rect 0 6974 3575 6976
rect 0 6944 480 6974
rect 3509 6971 3575 6974
rect 3969 7034 4035 7037
rect 8109 7034 8175 7037
rect 3969 7032 8175 7034
rect 3969 6976 3974 7032
rect 4030 6976 8114 7032
rect 8170 6976 8175 7032
rect 3969 6974 8175 6976
rect 3969 6971 4035 6974
rect 8109 6971 8175 6974
rect 8293 7034 8359 7037
rect 16205 7034 16271 7037
rect 18597 7034 18663 7037
rect 8293 7032 11162 7034
rect 8293 6976 8298 7032
rect 8354 6976 11162 7032
rect 8293 6974 11162 6976
rect 8293 6971 8359 6974
rect 3785 6898 3851 6901
rect 10961 6898 11027 6901
rect 3785 6896 11027 6898
rect 3785 6840 3790 6896
rect 3846 6840 10966 6896
rect 11022 6840 11027 6896
rect 3785 6838 11027 6840
rect 11102 6898 11162 6974
rect 16205 7032 18663 7034
rect 16205 6976 16210 7032
rect 16266 6976 18602 7032
rect 18658 6976 18663 7032
rect 16205 6974 18663 6976
rect 16205 6971 16271 6974
rect 18597 6971 18663 6974
rect 24485 7034 24551 7037
rect 27153 7034 27219 7037
rect 24485 7032 27219 7034
rect 24485 6976 24490 7032
rect 24546 6976 27158 7032
rect 27214 6976 27219 7032
rect 24485 6974 27219 6976
rect 24485 6971 24551 6974
rect 27153 6971 27219 6974
rect 36997 7034 37063 7037
rect 39520 7034 40000 7064
rect 36997 7032 40000 7034
rect 36997 6976 37002 7032
rect 37058 6976 40000 7032
rect 36997 6974 40000 6976
rect 36997 6971 37063 6974
rect 39520 6944 40000 6974
rect 12433 6898 12499 6901
rect 18873 6898 18939 6901
rect 11102 6896 18939 6898
rect 11102 6840 12438 6896
rect 12494 6840 18878 6896
rect 18934 6840 18939 6896
rect 11102 6838 18939 6840
rect 3785 6835 3851 6838
rect 10961 6835 11027 6838
rect 12433 6835 12499 6838
rect 18873 6835 18939 6838
rect 20161 6898 20227 6901
rect 22369 6898 22435 6901
rect 20161 6896 22435 6898
rect 20161 6840 20166 6896
rect 20222 6840 22374 6896
rect 22430 6840 22435 6896
rect 20161 6838 22435 6840
rect 20161 6835 20227 6838
rect 22369 6835 22435 6838
rect 34881 6898 34947 6901
rect 36169 6898 36235 6901
rect 34881 6896 36235 6898
rect 34881 6840 34886 6896
rect 34942 6840 36174 6896
rect 36230 6840 36235 6896
rect 34881 6838 36235 6840
rect 34881 6835 34947 6838
rect 36169 6835 36235 6838
rect 7097 6762 7163 6765
rect 7557 6762 7623 6765
rect 9949 6762 10015 6765
rect 10501 6762 10567 6765
rect 12249 6762 12315 6765
rect 17033 6762 17099 6765
rect 27061 6762 27127 6765
rect 7097 6760 8218 6762
rect 7097 6704 7102 6760
rect 7158 6704 7562 6760
rect 7618 6704 8218 6760
rect 7097 6702 8218 6704
rect 7097 6699 7163 6702
rect 7557 6699 7623 6702
rect 0 6626 480 6656
rect 2037 6626 2103 6629
rect 0 6624 2103 6626
rect 0 6568 2042 6624
rect 2098 6568 2103 6624
rect 0 6566 2103 6568
rect 8158 6626 8218 6702
rect 9949 6760 17099 6762
rect 9949 6704 9954 6760
rect 10010 6704 10506 6760
rect 10562 6704 12254 6760
rect 12310 6704 17038 6760
rect 17094 6704 17099 6760
rect 9949 6702 17099 6704
rect 9949 6699 10015 6702
rect 10501 6699 10567 6702
rect 12249 6699 12315 6702
rect 17033 6699 17099 6702
rect 17174 6760 27127 6762
rect 17174 6704 27066 6760
rect 27122 6704 27127 6760
rect 17174 6702 27127 6704
rect 17174 6626 17234 6702
rect 27061 6699 27127 6702
rect 27337 6762 27403 6765
rect 30373 6762 30439 6765
rect 27337 6760 30439 6762
rect 27337 6704 27342 6760
rect 27398 6704 30378 6760
rect 30434 6704 30439 6760
rect 27337 6702 30439 6704
rect 27337 6699 27403 6702
rect 30373 6699 30439 6702
rect 8158 6566 17234 6626
rect 24117 6626 24183 6629
rect 26969 6626 27035 6629
rect 27889 6626 27955 6629
rect 24117 6624 27955 6626
rect 24117 6568 24122 6624
rect 24178 6568 26974 6624
rect 27030 6568 27894 6624
rect 27950 6568 27955 6624
rect 24117 6566 27955 6568
rect 0 6536 480 6566
rect 2037 6563 2103 6566
rect 24117 6563 24183 6566
rect 26969 6563 27035 6566
rect 27889 6563 27955 6566
rect 35709 6626 35775 6629
rect 39520 6626 40000 6656
rect 35709 6624 40000 6626
rect 35709 6568 35714 6624
rect 35770 6568 40000 6624
rect 35709 6566 40000 6568
rect 35709 6563 35775 6566
rect 7610 6560 7930 6561
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7930 6560
rect 7610 6495 7930 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 34277 6560 34597 6561
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 39520 6536 40000 6566
rect 34277 6495 34597 6496
rect 6269 6492 6335 6493
rect 6269 6490 6316 6492
rect 6224 6488 6316 6490
rect 6224 6432 6274 6488
rect 6224 6430 6316 6432
rect 6269 6428 6316 6430
rect 6380 6428 6386 6492
rect 12157 6490 12223 6493
rect 14641 6490 14707 6493
rect 16665 6490 16731 6493
rect 25405 6492 25471 6493
rect 25405 6490 25452 6492
rect 12157 6488 14474 6490
rect 12157 6432 12162 6488
rect 12218 6432 14474 6488
rect 12157 6430 14474 6432
rect 6269 6427 6335 6428
rect 12157 6427 12223 6430
rect 5809 6354 5875 6357
rect 9857 6354 9923 6357
rect 5809 6352 9923 6354
rect 5809 6296 5814 6352
rect 5870 6296 9862 6352
rect 9918 6296 9923 6352
rect 5809 6294 9923 6296
rect 5809 6291 5875 6294
rect 9857 6291 9923 6294
rect 11421 6354 11487 6357
rect 13997 6354 14063 6357
rect 11421 6352 14063 6354
rect 11421 6296 11426 6352
rect 11482 6296 14002 6352
rect 14058 6296 14063 6352
rect 11421 6294 14063 6296
rect 14414 6354 14474 6430
rect 14641 6488 16731 6490
rect 14641 6432 14646 6488
rect 14702 6432 16670 6488
rect 16726 6432 16731 6488
rect 14641 6430 16731 6432
rect 25360 6488 25452 6490
rect 25360 6432 25410 6488
rect 25360 6430 25452 6432
rect 14641 6427 14707 6430
rect 16665 6427 16731 6430
rect 25405 6428 25452 6430
rect 25516 6428 25522 6492
rect 25773 6490 25839 6493
rect 30465 6490 30531 6493
rect 25773 6488 30531 6490
rect 25773 6432 25778 6488
rect 25834 6432 30470 6488
rect 30526 6432 30531 6488
rect 25773 6430 30531 6432
rect 25405 6427 25471 6428
rect 25773 6427 25839 6430
rect 30465 6427 30531 6430
rect 35934 6428 35940 6492
rect 36004 6490 36010 6492
rect 36077 6490 36143 6493
rect 36004 6488 36143 6490
rect 36004 6432 36082 6488
rect 36138 6432 36143 6488
rect 36004 6430 36143 6432
rect 36004 6428 36010 6430
rect 36077 6427 36143 6430
rect 14733 6354 14799 6357
rect 14414 6352 14799 6354
rect 14414 6296 14738 6352
rect 14794 6296 14799 6352
rect 14414 6294 14799 6296
rect 11421 6291 11487 6294
rect 13997 6291 14063 6294
rect 14733 6291 14799 6294
rect 18229 6354 18295 6357
rect 26877 6354 26943 6357
rect 28993 6354 29059 6357
rect 29729 6354 29795 6357
rect 35065 6354 35131 6357
rect 18229 6352 27170 6354
rect 18229 6296 18234 6352
rect 18290 6296 26882 6352
rect 26938 6296 27170 6352
rect 18229 6294 27170 6296
rect 18229 6291 18295 6294
rect 26877 6291 26943 6294
rect 0 6218 480 6248
rect 6637 6218 6703 6221
rect 0 6216 6703 6218
rect 0 6160 6642 6216
rect 6698 6160 6703 6216
rect 0 6158 6703 6160
rect 0 6128 480 6158
rect 6637 6155 6703 6158
rect 13997 6218 14063 6221
rect 18137 6218 18203 6221
rect 13997 6216 18203 6218
rect 13997 6160 14002 6216
rect 14058 6160 18142 6216
rect 18198 6160 18203 6216
rect 13997 6158 18203 6160
rect 13997 6155 14063 6158
rect 18137 6155 18203 6158
rect 24577 6218 24643 6221
rect 26601 6218 26667 6221
rect 24577 6216 26667 6218
rect 24577 6160 24582 6216
rect 24638 6160 26606 6216
rect 26662 6160 26667 6216
rect 24577 6158 26667 6160
rect 27110 6218 27170 6294
rect 28993 6352 35131 6354
rect 28993 6296 28998 6352
rect 29054 6296 29734 6352
rect 29790 6296 35070 6352
rect 35126 6296 35131 6352
rect 28993 6294 35131 6296
rect 28993 6291 29059 6294
rect 29729 6291 29795 6294
rect 35065 6291 35131 6294
rect 39520 6218 40000 6248
rect 27110 6158 40000 6218
rect 24577 6155 24643 6158
rect 26601 6155 26667 6158
rect 39520 6128 40000 6158
rect 14733 6082 14799 6085
rect 16849 6082 16915 6085
rect 20805 6082 20871 6085
rect 14733 6080 20871 6082
rect 14733 6024 14738 6080
rect 14794 6024 16854 6080
rect 16910 6024 20810 6080
rect 20866 6024 20871 6080
rect 14733 6022 20871 6024
rect 14733 6019 14799 6022
rect 16849 6019 16915 6022
rect 20805 6019 20871 6022
rect 28625 6082 28691 6085
rect 35893 6082 35959 6085
rect 28625 6080 35959 6082
rect 28625 6024 28630 6080
rect 28686 6024 35898 6080
rect 35954 6024 35959 6080
rect 28625 6022 35959 6024
rect 28625 6019 28691 6022
rect 35893 6019 35959 6022
rect 14277 6016 14597 6017
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 27610 6016 27930 6017
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 5951 27930 5952
rect 6085 5946 6151 5949
rect 9673 5946 9739 5949
rect 25405 5946 25471 5949
rect 6085 5944 9739 5946
rect 6085 5888 6090 5944
rect 6146 5888 9678 5944
rect 9734 5888 9739 5944
rect 6085 5886 9739 5888
rect 6085 5883 6151 5886
rect 9673 5883 9739 5886
rect 17174 5944 25471 5946
rect 17174 5888 25410 5944
rect 25466 5888 25471 5944
rect 17174 5886 25471 5888
rect 0 5810 480 5840
rect 9949 5810 10015 5813
rect 0 5808 10015 5810
rect 0 5752 9954 5808
rect 10010 5752 10015 5808
rect 0 5750 10015 5752
rect 0 5720 480 5750
rect 9949 5747 10015 5750
rect 10317 5810 10383 5813
rect 17174 5810 17234 5886
rect 25405 5883 25471 5886
rect 28165 5946 28231 5949
rect 32857 5946 32923 5949
rect 28165 5944 32923 5946
rect 28165 5888 28170 5944
rect 28226 5888 32862 5944
rect 32918 5888 32923 5944
rect 28165 5886 32923 5888
rect 28165 5883 28231 5886
rect 32857 5883 32923 5886
rect 33041 5946 33107 5949
rect 34973 5946 35039 5949
rect 33041 5944 35039 5946
rect 33041 5888 33046 5944
rect 33102 5888 34978 5944
rect 35034 5888 35039 5944
rect 33041 5886 35039 5888
rect 33041 5883 33107 5886
rect 34973 5883 35039 5886
rect 10317 5808 17234 5810
rect 10317 5752 10322 5808
rect 10378 5752 17234 5808
rect 10317 5750 17234 5752
rect 17309 5810 17375 5813
rect 21541 5810 21607 5813
rect 17309 5808 21607 5810
rect 17309 5752 17314 5808
rect 17370 5752 21546 5808
rect 21602 5752 21607 5808
rect 17309 5750 21607 5752
rect 10317 5747 10383 5750
rect 17309 5747 17375 5750
rect 21541 5747 21607 5750
rect 21817 5810 21883 5813
rect 28993 5810 29059 5813
rect 21817 5808 29059 5810
rect 21817 5752 21822 5808
rect 21878 5752 28998 5808
rect 29054 5752 29059 5808
rect 21817 5750 29059 5752
rect 21817 5747 21883 5750
rect 28993 5747 29059 5750
rect 30465 5810 30531 5813
rect 33409 5810 33475 5813
rect 30465 5808 33475 5810
rect 30465 5752 30470 5808
rect 30526 5752 33414 5808
rect 33470 5752 33475 5808
rect 30465 5750 33475 5752
rect 30465 5747 30531 5750
rect 33409 5747 33475 5750
rect 35801 5810 35867 5813
rect 39520 5810 40000 5840
rect 35801 5808 40000 5810
rect 35801 5752 35806 5808
rect 35862 5752 40000 5808
rect 35801 5750 40000 5752
rect 35801 5747 35867 5750
rect 39520 5720 40000 5750
rect 17401 5676 17467 5677
rect 17350 5612 17356 5676
rect 17420 5674 17467 5676
rect 18229 5674 18295 5677
rect 17420 5672 18295 5674
rect 17462 5616 18234 5672
rect 18290 5616 18295 5672
rect 17420 5614 18295 5616
rect 17420 5612 17467 5614
rect 17401 5611 17467 5612
rect 18229 5611 18295 5614
rect 24301 5674 24367 5677
rect 24669 5674 24735 5677
rect 27429 5674 27495 5677
rect 24301 5672 27495 5674
rect 24301 5616 24306 5672
rect 24362 5616 24674 5672
rect 24730 5616 27434 5672
rect 27490 5616 27495 5672
rect 24301 5614 27495 5616
rect 24301 5611 24367 5614
rect 24669 5611 24735 5614
rect 27429 5611 27495 5614
rect 33409 5674 33475 5677
rect 35985 5674 36051 5677
rect 33409 5672 36051 5674
rect 33409 5616 33414 5672
rect 33470 5616 35990 5672
rect 36046 5616 36051 5672
rect 33409 5614 36051 5616
rect 33409 5611 33475 5614
rect 35985 5611 36051 5614
rect 11421 5538 11487 5541
rect 16481 5538 16547 5541
rect 11421 5536 16547 5538
rect 11421 5480 11426 5536
rect 11482 5480 16486 5536
rect 16542 5480 16547 5536
rect 11421 5478 16547 5480
rect 11421 5475 11487 5478
rect 16481 5475 16547 5478
rect 25589 5538 25655 5541
rect 29729 5538 29795 5541
rect 25589 5536 29795 5538
rect 25589 5480 25594 5536
rect 25650 5480 29734 5536
rect 29790 5480 29795 5536
rect 25589 5478 29795 5480
rect 25589 5475 25655 5478
rect 29729 5475 29795 5478
rect 7610 5472 7930 5473
rect 0 5402 480 5432
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7930 5472
rect 7610 5407 7930 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 34277 5472 34597 5473
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 5407 34597 5408
rect 3693 5402 3759 5405
rect 0 5400 3759 5402
rect 0 5344 3698 5400
rect 3754 5344 3759 5400
rect 0 5342 3759 5344
rect 0 5312 480 5342
rect 3693 5339 3759 5342
rect 8109 5402 8175 5405
rect 17769 5402 17835 5405
rect 19517 5402 19583 5405
rect 8109 5400 17835 5402
rect 8109 5344 8114 5400
rect 8170 5344 17774 5400
rect 17830 5344 17835 5400
rect 8109 5342 17835 5344
rect 8109 5339 8175 5342
rect 17769 5339 17835 5342
rect 18278 5400 19583 5402
rect 18278 5344 19522 5400
rect 19578 5344 19583 5400
rect 18278 5342 19583 5344
rect 3509 5266 3575 5269
rect 8753 5266 8819 5269
rect 18278 5266 18338 5342
rect 19517 5339 19583 5342
rect 27429 5402 27495 5405
rect 33501 5402 33567 5405
rect 27429 5400 33567 5402
rect 27429 5344 27434 5400
rect 27490 5344 33506 5400
rect 33562 5344 33567 5400
rect 27429 5342 33567 5344
rect 27429 5339 27495 5342
rect 3509 5264 8819 5266
rect 3509 5208 3514 5264
rect 3570 5208 8758 5264
rect 8814 5208 8819 5264
rect 3509 5206 8819 5208
rect 3509 5203 3575 5206
rect 8753 5203 8819 5206
rect 9078 5206 18338 5266
rect 18505 5266 18571 5269
rect 26785 5266 26851 5269
rect 18505 5264 26851 5266
rect 18505 5208 18510 5264
rect 18566 5208 26790 5264
rect 26846 5208 26851 5264
rect 18505 5206 26851 5208
rect 33366 5266 33426 5342
rect 33501 5339 33567 5342
rect 36629 5402 36695 5405
rect 39520 5402 40000 5432
rect 36629 5400 40000 5402
rect 36629 5344 36634 5400
rect 36690 5344 40000 5400
rect 36629 5342 40000 5344
rect 36629 5339 36695 5342
rect 39520 5312 40000 5342
rect 34789 5266 34855 5269
rect 33366 5264 34855 5266
rect 33366 5208 34794 5264
rect 34850 5208 34855 5264
rect 33366 5206 34855 5208
rect 3141 5130 3207 5133
rect 8937 5130 9003 5133
rect 3141 5128 9003 5130
rect 3141 5072 3146 5128
rect 3202 5072 8942 5128
rect 8998 5072 9003 5128
rect 3141 5070 9003 5072
rect 3141 5067 3207 5070
rect 8937 5067 9003 5070
rect 0 4994 480 5024
rect 2405 4994 2471 4997
rect 4889 4994 4955 4997
rect 0 4934 1410 4994
rect 0 4904 480 4934
rect 1350 4858 1410 4934
rect 2405 4992 4955 4994
rect 2405 4936 2410 4992
rect 2466 4936 4894 4992
rect 4950 4936 4955 4992
rect 2405 4934 4955 4936
rect 2405 4931 2471 4934
rect 4889 4931 4955 4934
rect 5073 4994 5139 4997
rect 9078 4994 9138 5206
rect 18505 5203 18571 5206
rect 26785 5203 26851 5206
rect 34789 5203 34855 5206
rect 9581 5130 9647 5133
rect 18597 5132 18663 5133
rect 18597 5130 18644 5132
rect 9581 5128 17234 5130
rect 9581 5072 9586 5128
rect 9642 5072 17234 5128
rect 9581 5070 17234 5072
rect 18552 5128 18644 5130
rect 18552 5072 18602 5128
rect 18552 5070 18644 5072
rect 9581 5067 9647 5070
rect 5073 4992 9138 4994
rect 5073 4936 5078 4992
rect 5134 4936 9138 4992
rect 5073 4934 9138 4936
rect 17174 4994 17234 5070
rect 18597 5068 18644 5070
rect 18708 5068 18714 5132
rect 18781 5130 18847 5133
rect 23657 5130 23723 5133
rect 28441 5130 28507 5133
rect 18781 5128 28507 5130
rect 18781 5072 18786 5128
rect 18842 5072 23662 5128
rect 23718 5072 28446 5128
rect 28502 5072 28507 5128
rect 18781 5070 28507 5072
rect 18597 5067 18663 5068
rect 18781 5067 18847 5070
rect 23657 5067 23723 5070
rect 28441 5067 28507 5070
rect 30557 5130 30623 5133
rect 33225 5130 33291 5133
rect 30557 5128 33291 5130
rect 30557 5072 30562 5128
rect 30618 5072 33230 5128
rect 33286 5072 33291 5128
rect 30557 5070 33291 5072
rect 30557 5067 30623 5070
rect 33225 5067 33291 5070
rect 25313 4994 25379 4997
rect 17174 4992 25379 4994
rect 17174 4936 25318 4992
rect 25374 4936 25379 4992
rect 17174 4934 25379 4936
rect 5073 4931 5139 4934
rect 25313 4931 25379 4934
rect 30373 4994 30439 4997
rect 33685 4994 33751 4997
rect 39520 4994 40000 5024
rect 30373 4992 33751 4994
rect 30373 4936 30378 4992
rect 30434 4936 33690 4992
rect 33746 4936 33751 4992
rect 30373 4934 33751 4936
rect 30373 4931 30439 4934
rect 33685 4931 33751 4934
rect 35574 4934 40000 4994
rect 14277 4928 14597 4929
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 27610 4928 27930 4929
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 4863 27930 4864
rect 4061 4858 4127 4861
rect 1350 4856 4127 4858
rect 1350 4800 4066 4856
rect 4122 4800 4127 4856
rect 1350 4798 4127 4800
rect 4061 4795 4127 4798
rect 9489 4858 9555 4861
rect 12525 4858 12591 4861
rect 9489 4856 12591 4858
rect 9489 4800 9494 4856
rect 9550 4800 12530 4856
rect 12586 4800 12591 4856
rect 9489 4798 12591 4800
rect 9489 4795 9555 4798
rect 12525 4795 12591 4798
rect 16389 4858 16455 4861
rect 18137 4858 18203 4861
rect 16389 4856 18203 4858
rect 16389 4800 16394 4856
rect 16450 4800 18142 4856
rect 18198 4800 18203 4856
rect 16389 4798 18203 4800
rect 16389 4795 16455 4798
rect 18137 4795 18203 4798
rect 30925 4858 30991 4861
rect 35574 4858 35634 4934
rect 39520 4904 40000 4934
rect 30925 4856 35634 4858
rect 30925 4800 30930 4856
rect 30986 4800 35634 4856
rect 30925 4798 35634 4800
rect 30925 4795 30991 4798
rect 2497 4722 2563 4725
rect 18597 4722 18663 4725
rect 2497 4720 18663 4722
rect 2497 4664 2502 4720
rect 2558 4664 18602 4720
rect 18658 4664 18663 4720
rect 2497 4662 18663 4664
rect 2497 4659 2563 4662
rect 18597 4659 18663 4662
rect 19793 4722 19859 4725
rect 30465 4722 30531 4725
rect 19793 4720 30531 4722
rect 19793 4664 19798 4720
rect 19854 4664 30470 4720
rect 30526 4664 30531 4720
rect 19793 4662 30531 4664
rect 19793 4659 19859 4662
rect 30465 4659 30531 4662
rect 32857 4722 32923 4725
rect 33317 4722 33383 4725
rect 34605 4722 34671 4725
rect 32857 4720 34671 4722
rect 32857 4664 32862 4720
rect 32918 4664 33322 4720
rect 33378 4664 34610 4720
rect 34666 4664 34671 4720
rect 32857 4662 34671 4664
rect 32857 4659 32923 4662
rect 33317 4659 33383 4662
rect 34605 4659 34671 4662
rect 0 4586 480 4616
rect 3601 4586 3667 4589
rect 0 4584 3667 4586
rect 0 4528 3606 4584
rect 3662 4528 3667 4584
rect 0 4526 3667 4528
rect 0 4496 480 4526
rect 3601 4523 3667 4526
rect 7465 4586 7531 4589
rect 10133 4586 10199 4589
rect 7465 4584 10199 4586
rect 7465 4528 7470 4584
rect 7526 4528 10138 4584
rect 10194 4528 10199 4584
rect 7465 4526 10199 4528
rect 7465 4523 7531 4526
rect 10133 4523 10199 4526
rect 33777 4586 33843 4589
rect 39520 4586 40000 4616
rect 33777 4584 40000 4586
rect 33777 4528 33782 4584
rect 33838 4528 40000 4584
rect 33777 4526 40000 4528
rect 33777 4523 33843 4526
rect 39520 4496 40000 4526
rect 7610 4384 7930 4385
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7930 4384
rect 7610 4319 7930 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 34277 4384 34597 4385
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 4319 34597 4320
rect 18781 4314 18847 4317
rect 8158 4312 18847 4314
rect 8158 4256 18786 4312
rect 18842 4256 18847 4312
rect 8158 4254 18847 4256
rect 0 4178 480 4208
rect 2221 4178 2287 4181
rect 0 4176 2287 4178
rect 0 4120 2226 4176
rect 2282 4120 2287 4176
rect 0 4118 2287 4120
rect 0 4088 480 4118
rect 2221 4115 2287 4118
rect 4061 4178 4127 4181
rect 8158 4178 8218 4254
rect 18781 4251 18847 4254
rect 4061 4176 8218 4178
rect 4061 4120 4066 4176
rect 4122 4120 8218 4176
rect 4061 4118 8218 4120
rect 8937 4178 9003 4181
rect 25129 4178 25195 4181
rect 8937 4176 25195 4178
rect 8937 4120 8942 4176
rect 8998 4120 25134 4176
rect 25190 4120 25195 4176
rect 8937 4118 25195 4120
rect 4061 4115 4127 4118
rect 8937 4115 9003 4118
rect 25129 4115 25195 4118
rect 25313 4178 25379 4181
rect 35433 4178 35499 4181
rect 25313 4176 35499 4178
rect 25313 4120 25318 4176
rect 25374 4120 35438 4176
rect 35494 4120 35499 4176
rect 25313 4118 35499 4120
rect 25313 4115 25379 4118
rect 35433 4115 35499 4118
rect 35617 4178 35683 4181
rect 39520 4178 40000 4208
rect 35617 4176 40000 4178
rect 35617 4120 35622 4176
rect 35678 4120 40000 4176
rect 35617 4118 40000 4120
rect 35617 4115 35683 4118
rect 39520 4088 40000 4118
rect 4521 4042 4587 4045
rect 7189 4042 7255 4045
rect 4521 4040 7255 4042
rect 4521 3984 4526 4040
rect 4582 3984 7194 4040
rect 7250 3984 7255 4040
rect 4521 3982 7255 3984
rect 4521 3979 4587 3982
rect 7189 3979 7255 3982
rect 9213 4042 9279 4045
rect 18321 4042 18387 4045
rect 9213 4040 18387 4042
rect 9213 3984 9218 4040
rect 9274 3984 18326 4040
rect 18382 3984 18387 4040
rect 9213 3982 18387 3984
rect 9213 3979 9279 3982
rect 18321 3979 18387 3982
rect 21081 4042 21147 4045
rect 24301 4042 24367 4045
rect 21081 4040 24367 4042
rect 21081 3984 21086 4040
rect 21142 3984 24306 4040
rect 24362 3984 24367 4040
rect 21081 3982 24367 3984
rect 21081 3979 21147 3982
rect 24301 3979 24367 3982
rect 30557 4042 30623 4045
rect 35709 4042 35775 4045
rect 30557 4040 35775 4042
rect 30557 3984 30562 4040
rect 30618 3984 35714 4040
rect 35770 3984 35775 4040
rect 30557 3982 35775 3984
rect 30557 3979 30623 3982
rect 35709 3979 35775 3982
rect 3969 3906 4035 3909
rect 8661 3906 8727 3909
rect 3969 3904 8727 3906
rect 3969 3848 3974 3904
rect 4030 3848 8666 3904
rect 8722 3848 8727 3904
rect 3969 3846 8727 3848
rect 3969 3843 4035 3846
rect 8661 3843 8727 3846
rect 14277 3840 14597 3841
rect 0 3770 480 3800
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 27610 3840 27930 3841
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 3775 27930 3776
rect 4613 3770 4679 3773
rect 7097 3770 7163 3773
rect 0 3710 4538 3770
rect 0 3680 480 3710
rect 4478 3634 4538 3710
rect 4613 3768 7163 3770
rect 4613 3712 4618 3768
rect 4674 3712 7102 3768
rect 7158 3712 7163 3768
rect 4613 3710 7163 3712
rect 4613 3707 4679 3710
rect 7097 3707 7163 3710
rect 24577 3770 24643 3773
rect 26601 3770 26667 3773
rect 24577 3768 26667 3770
rect 24577 3712 24582 3768
rect 24638 3712 26606 3768
rect 26662 3712 26667 3768
rect 24577 3710 26667 3712
rect 24577 3707 24643 3710
rect 26601 3707 26667 3710
rect 30414 3708 30420 3772
rect 30484 3770 30490 3772
rect 31201 3770 31267 3773
rect 39520 3770 40000 3800
rect 30484 3768 40000 3770
rect 30484 3712 31206 3768
rect 31262 3712 40000 3768
rect 30484 3710 40000 3712
rect 30484 3708 30490 3710
rect 31201 3707 31267 3710
rect 39520 3680 40000 3710
rect 17677 3634 17743 3637
rect 4478 3632 17743 3634
rect 4478 3576 17682 3632
rect 17738 3576 17743 3632
rect 4478 3574 17743 3576
rect 17677 3571 17743 3574
rect 20437 3634 20503 3637
rect 29637 3634 29703 3637
rect 20437 3632 29703 3634
rect 20437 3576 20442 3632
rect 20498 3576 29642 3632
rect 29698 3576 29703 3632
rect 20437 3574 29703 3576
rect 20437 3571 20503 3574
rect 29637 3571 29703 3574
rect 0 3362 480 3392
rect 3969 3362 4035 3365
rect 0 3360 4035 3362
rect 0 3304 3974 3360
rect 4030 3304 4035 3360
rect 0 3302 4035 3304
rect 0 3272 480 3302
rect 3969 3299 4035 3302
rect 9673 3362 9739 3365
rect 19333 3362 19399 3365
rect 9673 3360 19399 3362
rect 9673 3304 9678 3360
rect 9734 3304 19338 3360
rect 19394 3304 19399 3360
rect 9673 3302 19399 3304
rect 9673 3299 9739 3302
rect 19333 3299 19399 3302
rect 23013 3362 23079 3365
rect 24945 3362 25011 3365
rect 39520 3362 40000 3392
rect 23013 3360 25011 3362
rect 23013 3304 23018 3360
rect 23074 3304 24950 3360
rect 25006 3304 25011 3360
rect 23013 3302 25011 3304
rect 23013 3299 23079 3302
rect 24945 3299 25011 3302
rect 35574 3302 40000 3362
rect 7610 3296 7930 3297
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7930 3296
rect 7610 3231 7930 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 34277 3296 34597 3297
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 3231 34597 3232
rect 5257 3090 5323 3093
rect 20529 3090 20595 3093
rect 35574 3090 35634 3302
rect 39520 3272 40000 3302
rect 5257 3088 20595 3090
rect 5257 3032 5262 3088
rect 5318 3032 20534 3088
rect 20590 3032 20595 3088
rect 22142 3056 35634 3090
rect 5257 3030 20595 3032
rect 5257 3027 5323 3030
rect 20529 3027 20595 3030
rect 22004 3030 35634 3056
rect 22004 2996 22202 3030
rect 0 2954 480 2984
rect 10317 2954 10383 2957
rect 0 2952 10383 2954
rect 0 2896 10322 2952
rect 10378 2896 10383 2952
rect 0 2894 10383 2896
rect 0 2864 480 2894
rect 10317 2891 10383 2894
rect 18873 2954 18939 2957
rect 22004 2954 22064 2996
rect 18873 2952 22064 2954
rect 18873 2896 18878 2952
rect 18934 2896 22064 2952
rect 18873 2894 22064 2896
rect 27337 2954 27403 2957
rect 28942 2954 28948 2956
rect 27337 2952 28948 2954
rect 27337 2896 27342 2952
rect 27398 2896 28948 2952
rect 27337 2894 28948 2896
rect 18873 2891 18939 2894
rect 27337 2891 27403 2894
rect 28942 2892 28948 2894
rect 29012 2892 29018 2956
rect 35801 2954 35867 2957
rect 39520 2954 40000 2984
rect 35801 2952 40000 2954
rect 35801 2896 35806 2952
rect 35862 2896 40000 2952
rect 35801 2894 40000 2896
rect 35801 2891 35867 2894
rect 39520 2864 40000 2894
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 27610 2752 27930 2753
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2687 27930 2688
rect 6913 2682 6979 2685
rect 2638 2680 6979 2682
rect 2638 2624 6918 2680
rect 6974 2624 6979 2680
rect 2638 2622 6979 2624
rect 0 2546 480 2576
rect 2638 2546 2698 2622
rect 6913 2619 6979 2622
rect 0 2486 2698 2546
rect 4337 2546 4403 2549
rect 14917 2546 14983 2549
rect 4337 2544 14983 2546
rect 4337 2488 4342 2544
rect 4398 2488 14922 2544
rect 14978 2488 14983 2544
rect 4337 2486 14983 2488
rect 0 2456 480 2486
rect 4337 2483 4403 2486
rect 14917 2483 14983 2486
rect 28942 2484 28948 2548
rect 29012 2546 29018 2548
rect 39520 2546 40000 2576
rect 29012 2486 40000 2546
rect 29012 2484 29018 2486
rect 39520 2456 40000 2486
rect 7610 2208 7930 2209
rect 0 2138 480 2168
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7930 2208
rect 7610 2143 7930 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 34277 2208 34597 2209
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2143 34597 2144
rect 3877 2138 3943 2141
rect 0 2136 3943 2138
rect 0 2080 3882 2136
rect 3938 2080 3943 2136
rect 0 2078 3943 2080
rect 0 2048 480 2078
rect 3877 2075 3943 2078
rect 35617 2138 35683 2141
rect 39520 2138 40000 2168
rect 35617 2136 40000 2138
rect 35617 2080 35622 2136
rect 35678 2080 40000 2136
rect 35617 2078 40000 2080
rect 35617 2075 35683 2078
rect 39520 2048 40000 2078
rect 0 1730 480 1760
rect 3141 1730 3207 1733
rect 0 1728 3207 1730
rect 0 1672 3146 1728
rect 3202 1672 3207 1728
rect 0 1670 3207 1672
rect 0 1640 480 1670
rect 3141 1667 3207 1670
rect 25129 1730 25195 1733
rect 39520 1730 40000 1760
rect 25129 1728 40000 1730
rect 25129 1672 25134 1728
rect 25190 1672 40000 1728
rect 25129 1670 40000 1672
rect 25129 1667 25195 1670
rect 39520 1640 40000 1670
rect 17217 1458 17283 1461
rect 35617 1458 35683 1461
rect 17217 1456 35683 1458
rect 17217 1400 17222 1456
rect 17278 1400 35622 1456
rect 35678 1400 35683 1456
rect 17217 1398 35683 1400
rect 17217 1395 17283 1398
rect 35617 1395 35683 1398
rect 0 1322 480 1352
rect 3233 1322 3299 1325
rect 0 1320 3299 1322
rect 0 1264 3238 1320
rect 3294 1264 3299 1320
rect 0 1262 3299 1264
rect 0 1232 480 1262
rect 3233 1259 3299 1262
rect 35341 1322 35407 1325
rect 39520 1322 40000 1352
rect 35341 1320 40000 1322
rect 35341 1264 35346 1320
rect 35402 1264 40000 1320
rect 35341 1262 40000 1264
rect 35341 1259 35407 1262
rect 39520 1232 40000 1262
rect 0 914 480 944
rect 3785 914 3851 917
rect 0 912 3851 914
rect 0 856 3790 912
rect 3846 856 3851 912
rect 0 854 3851 856
rect 0 824 480 854
rect 3785 851 3851 854
rect 34605 914 34671 917
rect 39520 914 40000 944
rect 34605 912 40000 914
rect 34605 856 34610 912
rect 34666 856 40000 912
rect 34605 854 40000 856
rect 34605 851 34671 854
rect 39520 824 40000 854
rect 0 506 480 536
rect 1301 506 1367 509
rect 0 504 1367 506
rect 0 448 1306 504
rect 1362 448 1367 504
rect 0 446 1367 448
rect 0 416 480 446
rect 1301 443 1367 446
rect 35157 506 35223 509
rect 39520 506 40000 536
rect 35157 504 40000 506
rect 35157 448 35162 504
rect 35218 448 40000 504
rect 35157 446 40000 448
rect 35157 443 35223 446
rect 39520 416 40000 446
rect 0 234 480 264
rect 2681 234 2747 237
rect 0 232 2747 234
rect 0 176 2686 232
rect 2742 176 2747 232
rect 0 174 2747 176
rect 0 144 480 174
rect 2681 171 2747 174
rect 34789 234 34855 237
rect 39520 234 40000 264
rect 34789 232 40000 234
rect 34789 176 34794 232
rect 34850 176 40000 232
rect 34789 174 40000 176
rect 34789 171 34855 174
rect 39520 144 40000 174
<< via3 >>
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 27618 13628 27682 13632
rect 27618 13572 27622 13628
rect 27622 13572 27678 13628
rect 27678 13572 27682 13628
rect 27618 13568 27682 13572
rect 27698 13628 27762 13632
rect 27698 13572 27702 13628
rect 27702 13572 27758 13628
rect 27758 13572 27762 13628
rect 27698 13568 27762 13572
rect 27778 13628 27842 13632
rect 27778 13572 27782 13628
rect 27782 13572 27838 13628
rect 27838 13572 27842 13628
rect 27778 13568 27842 13572
rect 27858 13628 27922 13632
rect 27858 13572 27862 13628
rect 27862 13572 27918 13628
rect 27918 13572 27922 13628
rect 27858 13568 27922 13572
rect 7618 13084 7682 13088
rect 7618 13028 7622 13084
rect 7622 13028 7678 13084
rect 7678 13028 7682 13084
rect 7618 13024 7682 13028
rect 7698 13084 7762 13088
rect 7698 13028 7702 13084
rect 7702 13028 7758 13084
rect 7758 13028 7762 13084
rect 7698 13024 7762 13028
rect 7778 13084 7842 13088
rect 7778 13028 7782 13084
rect 7782 13028 7838 13084
rect 7838 13028 7842 13084
rect 7778 13024 7842 13028
rect 7858 13084 7922 13088
rect 7858 13028 7862 13084
rect 7862 13028 7918 13084
rect 7918 13028 7922 13084
rect 7858 13024 7922 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 34285 13084 34349 13088
rect 34285 13028 34289 13084
rect 34289 13028 34345 13084
rect 34345 13028 34349 13084
rect 34285 13024 34349 13028
rect 34365 13084 34429 13088
rect 34365 13028 34369 13084
rect 34369 13028 34425 13084
rect 34425 13028 34429 13084
rect 34365 13024 34429 13028
rect 34445 13084 34509 13088
rect 34445 13028 34449 13084
rect 34449 13028 34505 13084
rect 34505 13028 34509 13084
rect 34445 13024 34509 13028
rect 34525 13084 34589 13088
rect 34525 13028 34529 13084
rect 34529 13028 34585 13084
rect 34585 13028 34589 13084
rect 34525 13024 34589 13028
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 27618 12540 27682 12544
rect 27618 12484 27622 12540
rect 27622 12484 27678 12540
rect 27678 12484 27682 12540
rect 27618 12480 27682 12484
rect 27698 12540 27762 12544
rect 27698 12484 27702 12540
rect 27702 12484 27758 12540
rect 27758 12484 27762 12540
rect 27698 12480 27762 12484
rect 27778 12540 27842 12544
rect 27778 12484 27782 12540
rect 27782 12484 27838 12540
rect 27838 12484 27842 12540
rect 27778 12480 27842 12484
rect 27858 12540 27922 12544
rect 27858 12484 27862 12540
rect 27862 12484 27918 12540
rect 27918 12484 27922 12540
rect 27858 12480 27922 12484
rect 33916 12140 33980 12204
rect 7618 11996 7682 12000
rect 7618 11940 7622 11996
rect 7622 11940 7678 11996
rect 7678 11940 7682 11996
rect 7618 11936 7682 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 34285 11996 34349 12000
rect 34285 11940 34289 11996
rect 34289 11940 34345 11996
rect 34345 11940 34349 11996
rect 34285 11936 34349 11940
rect 34365 11996 34429 12000
rect 34365 11940 34369 11996
rect 34369 11940 34425 11996
rect 34425 11940 34429 11996
rect 34365 11936 34429 11940
rect 34445 11996 34509 12000
rect 34445 11940 34449 11996
rect 34449 11940 34505 11996
rect 34505 11940 34509 11996
rect 34445 11936 34509 11940
rect 34525 11996 34589 12000
rect 34525 11940 34529 11996
rect 34529 11940 34585 11996
rect 34585 11940 34589 11996
rect 34525 11936 34589 11940
rect 4660 11868 4724 11932
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 27618 11452 27682 11456
rect 27618 11396 27622 11452
rect 27622 11396 27678 11452
rect 27678 11396 27682 11452
rect 27618 11392 27682 11396
rect 27698 11452 27762 11456
rect 27698 11396 27702 11452
rect 27702 11396 27758 11452
rect 27758 11396 27762 11452
rect 27698 11392 27762 11396
rect 27778 11452 27842 11456
rect 27778 11396 27782 11452
rect 27782 11396 27838 11452
rect 27838 11396 27842 11452
rect 27778 11392 27842 11396
rect 27858 11452 27922 11456
rect 27858 11396 27862 11452
rect 27862 11396 27918 11452
rect 27918 11396 27922 11452
rect 27858 11392 27922 11396
rect 7618 10908 7682 10912
rect 7618 10852 7622 10908
rect 7622 10852 7678 10908
rect 7678 10852 7682 10908
rect 7618 10848 7682 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 34285 10908 34349 10912
rect 34285 10852 34289 10908
rect 34289 10852 34345 10908
rect 34345 10852 34349 10908
rect 34285 10848 34349 10852
rect 34365 10908 34429 10912
rect 34365 10852 34369 10908
rect 34369 10852 34425 10908
rect 34425 10852 34429 10908
rect 34365 10848 34429 10852
rect 34445 10908 34509 10912
rect 34445 10852 34449 10908
rect 34449 10852 34505 10908
rect 34505 10852 34509 10908
rect 34445 10848 34509 10852
rect 34525 10908 34589 10912
rect 34525 10852 34529 10908
rect 34529 10852 34585 10908
rect 34585 10852 34589 10908
rect 34525 10848 34589 10852
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 27618 10364 27682 10368
rect 27618 10308 27622 10364
rect 27622 10308 27678 10364
rect 27678 10308 27682 10364
rect 27618 10304 27682 10308
rect 27698 10364 27762 10368
rect 27698 10308 27702 10364
rect 27702 10308 27758 10364
rect 27758 10308 27762 10364
rect 27698 10304 27762 10308
rect 27778 10364 27842 10368
rect 27778 10308 27782 10364
rect 27782 10308 27838 10364
rect 27838 10308 27842 10364
rect 27778 10304 27842 10308
rect 27858 10364 27922 10368
rect 27858 10308 27862 10364
rect 27862 10308 27918 10364
rect 27918 10308 27922 10364
rect 27858 10304 27922 10308
rect 7618 9820 7682 9824
rect 7618 9764 7622 9820
rect 7622 9764 7678 9820
rect 7678 9764 7682 9820
rect 7618 9760 7682 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 34285 9820 34349 9824
rect 34285 9764 34289 9820
rect 34289 9764 34345 9820
rect 34345 9764 34349 9820
rect 34285 9760 34349 9764
rect 34365 9820 34429 9824
rect 34365 9764 34369 9820
rect 34369 9764 34425 9820
rect 34425 9764 34429 9820
rect 34365 9760 34429 9764
rect 34445 9820 34509 9824
rect 34445 9764 34449 9820
rect 34449 9764 34505 9820
rect 34505 9764 34509 9820
rect 34445 9760 34509 9764
rect 34525 9820 34589 9824
rect 34525 9764 34529 9820
rect 34529 9764 34585 9820
rect 34585 9764 34589 9820
rect 34525 9760 34589 9764
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 27618 9276 27682 9280
rect 27618 9220 27622 9276
rect 27622 9220 27678 9276
rect 27678 9220 27682 9276
rect 27618 9216 27682 9220
rect 27698 9276 27762 9280
rect 27698 9220 27702 9276
rect 27702 9220 27758 9276
rect 27758 9220 27762 9276
rect 27698 9216 27762 9220
rect 27778 9276 27842 9280
rect 27778 9220 27782 9276
rect 27782 9220 27838 9276
rect 27838 9220 27842 9276
rect 27778 9216 27842 9220
rect 27858 9276 27922 9280
rect 27858 9220 27862 9276
rect 27862 9220 27918 9276
rect 27918 9220 27922 9276
rect 27858 9216 27922 9220
rect 7618 8732 7682 8736
rect 7618 8676 7622 8732
rect 7622 8676 7678 8732
rect 7678 8676 7682 8732
rect 7618 8672 7682 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 34285 8732 34349 8736
rect 34285 8676 34289 8732
rect 34289 8676 34345 8732
rect 34345 8676 34349 8732
rect 34285 8672 34349 8676
rect 34365 8732 34429 8736
rect 34365 8676 34369 8732
rect 34369 8676 34425 8732
rect 34425 8676 34429 8732
rect 34365 8672 34429 8676
rect 34445 8732 34509 8736
rect 34445 8676 34449 8732
rect 34449 8676 34505 8732
rect 34505 8676 34509 8732
rect 34445 8672 34509 8676
rect 34525 8732 34589 8736
rect 34525 8676 34529 8732
rect 34529 8676 34585 8732
rect 34585 8676 34589 8732
rect 34525 8672 34589 8676
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 27618 8188 27682 8192
rect 27618 8132 27622 8188
rect 27622 8132 27678 8188
rect 27678 8132 27682 8188
rect 27618 8128 27682 8132
rect 27698 8188 27762 8192
rect 27698 8132 27702 8188
rect 27702 8132 27758 8188
rect 27758 8132 27762 8188
rect 27698 8128 27762 8132
rect 27778 8188 27842 8192
rect 27778 8132 27782 8188
rect 27782 8132 27838 8188
rect 27838 8132 27842 8188
rect 27778 8128 27842 8132
rect 27858 8188 27922 8192
rect 27858 8132 27862 8188
rect 27862 8132 27918 8188
rect 27918 8132 27922 8188
rect 27858 8128 27922 8132
rect 7618 7644 7682 7648
rect 7618 7588 7622 7644
rect 7622 7588 7678 7644
rect 7678 7588 7682 7644
rect 7618 7584 7682 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 34285 7644 34349 7648
rect 34285 7588 34289 7644
rect 34289 7588 34345 7644
rect 34345 7588 34349 7644
rect 34285 7584 34349 7588
rect 34365 7644 34429 7648
rect 34365 7588 34369 7644
rect 34369 7588 34425 7644
rect 34425 7588 34429 7644
rect 34365 7584 34429 7588
rect 34445 7644 34509 7648
rect 34445 7588 34449 7644
rect 34449 7588 34505 7644
rect 34505 7588 34509 7644
rect 34445 7584 34509 7588
rect 34525 7644 34589 7648
rect 34525 7588 34529 7644
rect 34529 7588 34585 7644
rect 34585 7588 34589 7644
rect 34525 7584 34589 7588
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 27618 7100 27682 7104
rect 27618 7044 27622 7100
rect 27622 7044 27678 7100
rect 27678 7044 27682 7100
rect 27618 7040 27682 7044
rect 27698 7100 27762 7104
rect 27698 7044 27702 7100
rect 27702 7044 27758 7100
rect 27758 7044 27762 7100
rect 27698 7040 27762 7044
rect 27778 7100 27842 7104
rect 27778 7044 27782 7100
rect 27782 7044 27838 7100
rect 27838 7044 27842 7100
rect 27778 7040 27842 7044
rect 27858 7100 27922 7104
rect 27858 7044 27862 7100
rect 27862 7044 27918 7100
rect 27918 7044 27922 7100
rect 27858 7040 27922 7044
rect 7618 6556 7682 6560
rect 7618 6500 7622 6556
rect 7622 6500 7678 6556
rect 7678 6500 7682 6556
rect 7618 6496 7682 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 34285 6556 34349 6560
rect 34285 6500 34289 6556
rect 34289 6500 34345 6556
rect 34345 6500 34349 6556
rect 34285 6496 34349 6500
rect 34365 6556 34429 6560
rect 34365 6500 34369 6556
rect 34369 6500 34425 6556
rect 34425 6500 34429 6556
rect 34365 6496 34429 6500
rect 34445 6556 34509 6560
rect 34445 6500 34449 6556
rect 34449 6500 34505 6556
rect 34505 6500 34509 6556
rect 34445 6496 34509 6500
rect 34525 6556 34589 6560
rect 34525 6500 34529 6556
rect 34529 6500 34585 6556
rect 34585 6500 34589 6556
rect 34525 6496 34589 6500
rect 6316 6488 6380 6492
rect 6316 6432 6330 6488
rect 6330 6432 6380 6488
rect 6316 6428 6380 6432
rect 25452 6488 25516 6492
rect 25452 6432 25466 6488
rect 25466 6432 25516 6488
rect 25452 6428 25516 6432
rect 35940 6428 36004 6492
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 27618 6012 27682 6016
rect 27618 5956 27622 6012
rect 27622 5956 27678 6012
rect 27678 5956 27682 6012
rect 27618 5952 27682 5956
rect 27698 6012 27762 6016
rect 27698 5956 27702 6012
rect 27702 5956 27758 6012
rect 27758 5956 27762 6012
rect 27698 5952 27762 5956
rect 27778 6012 27842 6016
rect 27778 5956 27782 6012
rect 27782 5956 27838 6012
rect 27838 5956 27842 6012
rect 27778 5952 27842 5956
rect 27858 6012 27922 6016
rect 27858 5956 27862 6012
rect 27862 5956 27918 6012
rect 27918 5956 27922 6012
rect 27858 5952 27922 5956
rect 17356 5672 17420 5676
rect 17356 5616 17406 5672
rect 17406 5616 17420 5672
rect 17356 5612 17420 5616
rect 7618 5468 7682 5472
rect 7618 5412 7622 5468
rect 7622 5412 7678 5468
rect 7678 5412 7682 5468
rect 7618 5408 7682 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 34285 5468 34349 5472
rect 34285 5412 34289 5468
rect 34289 5412 34345 5468
rect 34345 5412 34349 5468
rect 34285 5408 34349 5412
rect 34365 5468 34429 5472
rect 34365 5412 34369 5468
rect 34369 5412 34425 5468
rect 34425 5412 34429 5468
rect 34365 5408 34429 5412
rect 34445 5468 34509 5472
rect 34445 5412 34449 5468
rect 34449 5412 34505 5468
rect 34505 5412 34509 5468
rect 34445 5408 34509 5412
rect 34525 5468 34589 5472
rect 34525 5412 34529 5468
rect 34529 5412 34585 5468
rect 34585 5412 34589 5468
rect 34525 5408 34589 5412
rect 18644 5128 18708 5132
rect 18644 5072 18658 5128
rect 18658 5072 18708 5128
rect 18644 5068 18708 5072
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 27618 4924 27682 4928
rect 27618 4868 27622 4924
rect 27622 4868 27678 4924
rect 27678 4868 27682 4924
rect 27618 4864 27682 4868
rect 27698 4924 27762 4928
rect 27698 4868 27702 4924
rect 27702 4868 27758 4924
rect 27758 4868 27762 4924
rect 27698 4864 27762 4868
rect 27778 4924 27842 4928
rect 27778 4868 27782 4924
rect 27782 4868 27838 4924
rect 27838 4868 27842 4924
rect 27778 4864 27842 4868
rect 27858 4924 27922 4928
rect 27858 4868 27862 4924
rect 27862 4868 27918 4924
rect 27918 4868 27922 4924
rect 27858 4864 27922 4868
rect 7618 4380 7682 4384
rect 7618 4324 7622 4380
rect 7622 4324 7678 4380
rect 7678 4324 7682 4380
rect 7618 4320 7682 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 34285 4380 34349 4384
rect 34285 4324 34289 4380
rect 34289 4324 34345 4380
rect 34345 4324 34349 4380
rect 34285 4320 34349 4324
rect 34365 4380 34429 4384
rect 34365 4324 34369 4380
rect 34369 4324 34425 4380
rect 34425 4324 34429 4380
rect 34365 4320 34429 4324
rect 34445 4380 34509 4384
rect 34445 4324 34449 4380
rect 34449 4324 34505 4380
rect 34505 4324 34509 4380
rect 34445 4320 34509 4324
rect 34525 4380 34589 4384
rect 34525 4324 34529 4380
rect 34529 4324 34585 4380
rect 34585 4324 34589 4380
rect 34525 4320 34589 4324
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 27618 3836 27682 3840
rect 27618 3780 27622 3836
rect 27622 3780 27678 3836
rect 27678 3780 27682 3836
rect 27618 3776 27682 3780
rect 27698 3836 27762 3840
rect 27698 3780 27702 3836
rect 27702 3780 27758 3836
rect 27758 3780 27762 3836
rect 27698 3776 27762 3780
rect 27778 3836 27842 3840
rect 27778 3780 27782 3836
rect 27782 3780 27838 3836
rect 27838 3780 27842 3836
rect 27778 3776 27842 3780
rect 27858 3836 27922 3840
rect 27858 3780 27862 3836
rect 27862 3780 27918 3836
rect 27918 3780 27922 3836
rect 27858 3776 27922 3780
rect 30420 3708 30484 3772
rect 7618 3292 7682 3296
rect 7618 3236 7622 3292
rect 7622 3236 7678 3292
rect 7678 3236 7682 3292
rect 7618 3232 7682 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 34285 3292 34349 3296
rect 34285 3236 34289 3292
rect 34289 3236 34345 3292
rect 34345 3236 34349 3292
rect 34285 3232 34349 3236
rect 34365 3292 34429 3296
rect 34365 3236 34369 3292
rect 34369 3236 34425 3292
rect 34425 3236 34429 3292
rect 34365 3232 34429 3236
rect 34445 3292 34509 3296
rect 34445 3236 34449 3292
rect 34449 3236 34505 3292
rect 34505 3236 34509 3292
rect 34445 3232 34509 3236
rect 34525 3292 34589 3296
rect 34525 3236 34529 3292
rect 34529 3236 34585 3292
rect 34585 3236 34589 3292
rect 34525 3232 34589 3236
rect 28948 2892 29012 2956
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 27618 2748 27682 2752
rect 27618 2692 27622 2748
rect 27622 2692 27678 2748
rect 27678 2692 27682 2748
rect 27618 2688 27682 2692
rect 27698 2748 27762 2752
rect 27698 2692 27702 2748
rect 27702 2692 27758 2748
rect 27758 2692 27762 2748
rect 27698 2688 27762 2692
rect 27778 2748 27842 2752
rect 27778 2692 27782 2748
rect 27782 2692 27838 2748
rect 27838 2692 27842 2748
rect 27778 2688 27842 2692
rect 27858 2748 27922 2752
rect 27858 2692 27862 2748
rect 27862 2692 27918 2748
rect 27918 2692 27922 2748
rect 27858 2688 27922 2692
rect 28948 2484 29012 2548
rect 7618 2204 7682 2208
rect 7618 2148 7622 2204
rect 7622 2148 7678 2204
rect 7678 2148 7682 2204
rect 7618 2144 7682 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 34285 2204 34349 2208
rect 34285 2148 34289 2204
rect 34289 2148 34345 2204
rect 34345 2148 34349 2204
rect 34285 2144 34349 2148
rect 34365 2204 34429 2208
rect 34365 2148 34369 2204
rect 34369 2148 34425 2204
rect 34425 2148 34429 2204
rect 34365 2144 34429 2148
rect 34445 2204 34509 2208
rect 34445 2148 34449 2204
rect 34449 2148 34505 2204
rect 34505 2148 34509 2204
rect 34445 2144 34509 2148
rect 34525 2204 34589 2208
rect 34525 2148 34529 2204
rect 34529 2148 34585 2204
rect 34585 2148 34589 2204
rect 34525 2144 34589 2148
<< metal4 >>
rect 7610 13088 7931 13648
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7931 13088
rect 7610 12000 7931 13024
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7931 12000
rect 7610 10912 7931 11936
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7931 10912
rect 7610 9824 7931 10848
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7931 9824
rect 7610 8736 7931 9760
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7931 8736
rect 7610 7648 7931 8672
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7931 7648
rect 7610 6560 7931 7584
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7931 6560
rect 7610 5472 7931 6496
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7931 5472
rect 7610 4384 7931 5408
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7931 4384
rect 7610 3296 7931 4320
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7931 3296
rect 7610 2208 7931 3232
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7931 2208
rect 7610 2128 7931 2144
rect 14277 13632 14597 13648
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 9280 14597 10304
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 20944 13088 21264 13648
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 27610 13632 27930 13648
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 12544 27930 13568
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 11456 27930 12480
rect 34277 13088 34597 13648
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 33915 12204 33981 12205
rect 33915 12140 33916 12204
rect 33980 12140 33981 12204
rect 33915 12139 33981 12140
rect 33918 12018 33978 12139
rect 34277 12000 34597 13024
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 10368 27930 11392
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 9280 27930 10304
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 8192 27930 9216
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 7104 27930 8128
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 17358 5677 17418 6342
rect 17355 5676 17421 5677
rect 17355 5612 17356 5676
rect 17420 5612 17421 5676
rect 17355 5611 17421 5612
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 3840 14597 4864
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 2752 14597 3776
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 27610 6016 27930 7040
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 4928 27930 5952
rect 34277 10912 34597 11936
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 9824 34597 10848
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 8736 34597 9760
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 7648 34597 8672
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 6560 34597 7584
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 5472 34597 6496
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 3840 27930 4864
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 2752 27930 3776
rect 30422 3773 30482 4982
rect 34277 4384 34597 5408
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 30419 3772 30485 3773
rect 30419 3708 30420 3772
rect 30484 3708 30485 3772
rect 30419 3707 30485 3708
rect 34277 3296 34597 4320
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 28947 2956 29013 2957
rect 28947 2892 28948 2956
rect 29012 2892 29013 2956
rect 28947 2891 29013 2892
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2128 27930 2688
rect 28950 2549 29010 2891
rect 28947 2548 29013 2549
rect 28947 2484 28948 2548
rect 29012 2484 29013 2548
rect 28947 2483 29013 2484
rect 34277 2208 34597 3232
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2128 34597 2144
<< via4 >>
rect 4574 11932 4810 12018
rect 4574 11868 4660 11932
rect 4660 11868 4724 11932
rect 4724 11868 4810 11932
rect 4574 11782 4810 11868
rect 6230 6492 6466 6578
rect 6230 6428 6316 6492
rect 6316 6428 6380 6492
rect 6380 6428 6466 6492
rect 6230 6342 6466 6428
rect 17270 6342 17506 6578
rect 33830 11782 34066 12018
rect 25366 6492 25602 6578
rect 25366 6428 25452 6492
rect 25452 6428 25516 6492
rect 25516 6428 25602 6492
rect 25366 6342 25602 6428
rect 18558 5132 18794 5218
rect 18558 5068 18644 5132
rect 18644 5068 18708 5132
rect 18708 5068 18794 5132
rect 18558 4982 18794 5068
rect 35854 6492 36090 6578
rect 35854 6428 35940 6492
rect 35940 6428 36004 6492
rect 36004 6428 36090 6492
rect 35854 6342 36090 6428
rect 30334 4982 30570 5218
<< metal5 >>
rect 4532 12018 34108 12060
rect 4532 11782 4574 12018
rect 4810 11782 33830 12018
rect 34066 11782 34108 12018
rect 4532 11740 34108 11782
rect 6188 6578 17548 6620
rect 6188 6342 6230 6578
rect 6466 6342 17270 6578
rect 17506 6342 17548 6578
rect 6188 6300 17548 6342
rect 25324 6578 36132 6620
rect 25324 6342 25366 6578
rect 25602 6342 35854 6578
rect 36090 6342 36132 6578
rect 25324 6300 36132 6342
rect 18516 5218 30612 5260
rect 18516 4982 18558 5218
rect 18794 4982 30334 5218
rect 30570 4982 30612 5218
rect 18516 4940 30612 4982
use scs8hd_fill_1  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_7
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_3
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_14
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_10
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_18
timestamp 1586364061
transform 1 0 2760 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l1_in_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1786 592
use scs8hd_buf_4  mux_top_ipin_0.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_21
timestamp 1586364061
transform 1 0 3036 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_28 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_51
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_0_59
timestamp 1586364061
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_42
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_46 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5336 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_58
timestamp 1586364061
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_206
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_207
timestamp 1586364061
transform 1 0 20148 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 19872 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_212
timestamp 1586364061
transform 1 0 20608 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_ipin_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 866 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 21620 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_219
timestamp 1586364061
transform 1 0 21252 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_225
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_229
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_241
timestamp 1586364061
transform 1 0 23276 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_256
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_252
timestamp 1586364061
transform 1 0 24288 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_249
timestamp 1586364061
transform 1 0 24012 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 24104 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_260
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_272
timestamp 1586364061
transform 1 0 26128 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_292
timestamp 1586364061
transform 1 0 27968 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_284
timestamp 1586364061
transform 1 0 27232 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_296
timestamp 1586364061
transform 1 0 28336 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_304
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_311
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_304
timestamp 1586364061
transform 1 0 29072 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_323
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_318
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_330
timestamp 1586364061
transform 1 0 31464 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_354
timestamp 1586364061
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_342
timestamp 1586364061
transform 1 0 32568 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_354
timestamp 1586364061
transform 1 0 33672 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_17
timestamp 1586364061
transform 1 0 2668 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_21
timestamp 1586364061
transform 1 0 3036 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_25
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_29
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_36
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_40
timestamp 1586364061
transform 1 0 4784 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_52
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7912 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_72
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_76
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_86
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_90
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 21068 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_2  FILLER_2_210
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_ipin_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 21620 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_219
timestamp 1586364061
transform 1 0 21252 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_ipin_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 24104 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_242
timestamp 1586364061
transform 1 0 23368 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_247
timestamp 1586364061
transform 1 0 23828 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25116 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_259
timestamp 1586364061
transform 1 0 24932 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 27232 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 27600 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_286
timestamp 1586364061
transform 1 0 27416 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_290
timestamp 1586364061
transform 1 0 27784 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 29808 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 30176 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_302
timestamp 1586364061
transform 1 0 28888 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_310
timestamp 1586364061
transform 1 0 29624 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_314
timestamp 1586364061
transform 1 0 29992 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 30544 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_318
timestamp 1586364061
transform 1 0 30360 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_322
timestamp 1586364061
transform 1 0 30728 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_2_334
timestamp 1586364061
transform 1 0 31832 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_337
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_349
timestamp 1586364061
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_361
timestamp 1586364061
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_373
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_385
timestamp 1586364061
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_10
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_23
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_44
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_50
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_54
timestamp 1586364061
transform 1 0 6072 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_58
timestamp 1586364061
transform 1 0 6440 0 1 3808
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_76
timestamp 1586364061
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_80
timestamp 1586364061
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_93
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_105
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_3_117
timestamp 1586364061
transform 1 0 11868 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_121
timestamp 1586364061
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_162
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_166
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_170
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_182
timestamp 1586364061
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_ipin_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_199
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_203
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_207
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_211
timestamp 1586364061
transform 1 0 20516 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_233
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_238
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_ipin_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_242
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_254
timestamp 1586364061
transform 1 0 24472 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 25116 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 26312 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 25484 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_259
timestamp 1586364061
transform 1 0 24932 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_263
timestamp 1586364061
transform 1 0 25300 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_267
timestamp 1586364061
transform 1 0 25668 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_273
timestamp 1586364061
transform 1 0 26220 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_276
timestamp 1586364061
transform 1 0 26496 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l1_in_2_
timestamp 1586364061
transform 1 0 27232 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 27048 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 26680 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_280
timestamp 1586364061
transform 1 0 26864 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_293
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l2_in_3_
timestamp 1586364061
transform 1 0 29808 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 29624 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_301
timestamp 1586364061
transform 1 0 28796 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_306
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 30820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_321
timestamp 1586364061
transform 1 0 30636 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_325
timestamp 1586364061
transform 1 0 31004 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_337
timestamp 1586364061
transform 1 0 32108 0 1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 32844 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 33212 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 33580 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_347
timestamp 1586364061
transform 1 0 33028 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_351
timestamp 1586364061
transform 1 0 33396 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_355
timestamp 1586364061
transform 1 0 33764 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_3_363
timestamp 1586364061
transform 1 0 34500 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_379
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_391
timestamp 1586364061
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2300 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2116 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 3312 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_22
timestamp 1586364061
transform 1 0 3128 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_26
timestamp 1586364061
transform 1 0 3496 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 5980 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_51
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_55
timestamp 1586364061
transform 1 0 6164 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_59
timestamp 1586364061
transform 1 0 6532 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_62
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_75
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10120 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_83
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_86
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_4  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_97
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_104
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_100
timestamp 1586364061
transform 1 0 10304 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_108
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_112
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_116
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_119
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_123
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_135
timestamp 1586364061
transform 1 0 13524 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_147
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_4  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l3_in_1_
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_169
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_177
timestamp 1586364061
transform 1 0 17388 0 -1 4896
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_ipin_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_182
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_196
timestamp 1586364061
transform 1 0 19136 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_2  mux_top_ipin_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23000 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_228
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_236
timestamp 1586364061
transform 1 0 22816 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_ipin_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23184 0 -1 4896
box -38 -48 866 592
use scs8hd_mux2_2  mux_top_ipin_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 24748 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 24564 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_249
timestamp 1586364061
transform 1 0 24012 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_253
timestamp 1586364061
transform 1 0 24380 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25760 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_266
timestamp 1586364061
transform 1 0 25576 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_270
timestamp 1586364061
transform 1 0 25944 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 27232 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 27048 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 26680 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_280
timestamp 1586364061
transform 1 0 26864 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l4_in_0_
timestamp 1586364061
transform 1 0 29716 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 29532 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 29164 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_303
timestamp 1586364061
transform 1 0 28980 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_307
timestamp 1586364061
transform 1 0 29348 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 30728 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 31096 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_320
timestamp 1586364061
transform 1 0 30544 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_324
timestamp 1586364061
transform 1 0 30912 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_328
timestamp 1586364061
transform 1 0 31280 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l2_in_1_
timestamp 1586364061
transform 1 0 32844 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 32292 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 32660 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_341
timestamp 1586364061
transform 1 0 32476 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_354
timestamp 1586364061
transform 1 0 33672 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_366
timestamp 1586364061
transform 1 0 34776 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_378
timestamp 1586364061
transform 1 0 35880 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_4_390
timestamp 1586364061
transform 1 0 36984 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_396
timestamp 1586364061
transform 1 0 37536 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_2  _49_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_11
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_14
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_31
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_44
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_5_50
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_54
timestamp 1586364061
transform 1 0 6072 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_76
timestamp 1586364061
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_80
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_93
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_97
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l4_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 11868 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_100
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_119
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use scs8hd_conb_1  _31_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_126
timestamp 1586364061
transform 1 0 12696 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_130
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_5_138
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_146
timestamp 1586364061
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_142
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_154
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_150
timestamp 1586364061
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_167
timestamp 1586364061
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l2_in_2_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_198
timestamp 1586364061
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_ipin_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 19688 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_211
timestamp 1586364061
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_215
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_ipin_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 22632 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22264 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_228
timestamp 1586364061
transform 1 0 22080 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_ipin_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l2_in_0_
timestamp 1586364061
transform 1 0 25484 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 26496 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 25300 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_262
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_274
timestamp 1586364061
transform 1 0 26312 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l1_in_0_
timestamp 1586364061
transform 1 0 27048 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 26864 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 28428 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 28060 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_278
timestamp 1586364061
transform 1 0 26680 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_291
timestamp 1586364061
transform 1 0 27876 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_295
timestamp 1586364061
transform 1 0 28244 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l3_in_1_
timestamp 1586364061
transform 1 0 29532 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 28796 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_299
timestamp 1586364061
transform 1 0 28612 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_303
timestamp 1586364061
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_306
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_318
timestamp 1586364061
transform 1 0 30360 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 30544 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_322
timestamp 1586364061
transform 1 0 30728 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 30912 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_326
timestamp 1586364061
transform 1 0 31096 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 31280 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_330
timestamp 1586364061
transform 1 0 31464 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_335
timestamp 1586364061
transform 1 0 31924 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 31740 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 32108 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 32292 0 1 4896
box -38 -48 1786 592
use scs8hd_buf_2  _69_
timestamp 1586364061
transform 1 0 35420 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 34224 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 34592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_358
timestamp 1586364061
transform 1 0 34040 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_362
timestamp 1586364061
transform 1 0 34408 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__69__A
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_377
timestamp 1586364061
transform 1 0 35788 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_381
timestamp 1586364061
transform 1 0 36156 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_393
timestamp 1586364061
transform 1 0 37260 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_405
timestamp 1586364061
transform 1 0 38364 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_6_21
timestamp 1586364061
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_29
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_25
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_35
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_36
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4600 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_40
timestamp 1586364061
transform 1 0 4784 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 4968 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l4_in_0_
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l3_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_57
timestamp 1586364061
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7084 0 -1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_61
timestamp 1586364061
transform 1 0 6716 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_85
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_81
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_91
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9936 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10120 0 -1 5984
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l2_in_2_
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l3_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_107
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_113
timestamp 1586364061
transform 1 0 11500 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_126
timestamp 1586364061
transform 1 0 12696 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_134
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_130
timestamp 1586364061
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12604 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_4.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 15088 0 1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_144
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_148
timestamp 1586364061
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_161
timestamp 1586364061
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_172
timestamp 1586364061
transform 1 0 16928 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l2_in_3_
timestamp 1586364061
transform 1 0 17664 0 -1 5984
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_193
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_189
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_201
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 774 592
use scs8hd_decap_6  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_201
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _20_
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_213
timestamp 1586364061
transform 1 0 20700 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_209
timestamp 1586364061
transform 1 0 20332 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20516 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21068 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_ipin_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 22632 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_226
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_232
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l3_in_1_
timestamp 1586364061
transform 1 0 24012 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 23828 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_253
timestamp 1586364061
transform 1 0 24380 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_257
timestamp 1586364061
transform 1 0 24748 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_262
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_258
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_264
timestamp 1586364061
transform 1 0 25392 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_260
timestamp 1586364061
transform 1 0 25024 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25208 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 24840 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 25576 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 25392 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_272
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_268
timestamp 1586364061
transform 1 0 25760 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25944 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 25576 0 1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_7_285
timestamp 1586364061
transform 1 0 27324 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 27508 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 26680 0 -1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l1_in_1_
timestamp 1586364061
transform 1 0 26864 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_297
timestamp 1586364061
transform 1 0 28428 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_293
timestamp 1586364061
transform 1 0 28060 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_289
timestamp 1586364061
transform 1 0 27692 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_293
timestamp 1586364061
transform 1 0 28060 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_289
timestamp 1586364061
transform 1 0 27692 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 27876 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 27876 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l2_in_1_
timestamp 1586364061
transform 1 0 28428 0 -1 5984
box -38 -48 866 592
use scs8hd_conb_1  _25_
timestamp 1586364061
transform 1 0 28152 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_301
timestamp 1586364061
transform 1 0 28796 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_306
timestamp 1586364061
transform 1 0 29256 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 28612 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 28980 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l3_in_0_
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_315
timestamp 1586364061
transform 1 0 30084 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_310
timestamp 1586364061
transform 1 0 29624 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 29808 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 30268 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 29440 0 -1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_12.mux_l2_in_2_
timestamp 1586364061
transform 1 0 29992 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_12.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 31004 0 1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 30820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 31004 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_323
timestamp 1586364061
transform 1 0 30820 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_327
timestamp 1586364061
transform 1 0 31188 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_335
timestamp 1586364061
transform 1 0 31924 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_337
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_319
timestamp 1586364061
transform 1 0 30452 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_344
timestamp 1586364061
transform 1 0 32752 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 32384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 32936 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l2_in_0_
timestamp 1586364061
transform 1 0 32568 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_1  FILLER_7_356
timestamp 1586364061
transform 1 0 33856 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_352
timestamp 1586364061
transform 1 0 33488 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_348
timestamp 1586364061
transform 1 0 33120 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_355
timestamp 1586364061
transform 1 0 33764 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_351
timestamp 1586364061
transform 1 0 33396 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 33580 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 33304 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 33948 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 34132 0 -1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 35236 0 1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 34316 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 35052 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_359
timestamp 1586364061
transform 1 0 34132 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_363
timestamp 1586364061
transform 1 0 34500 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_367
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 36064 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 36432 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 37168 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_378
timestamp 1586364061
transform 1 0 35880 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_382
timestamp 1586364061
transform 1 0 36248 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_386
timestamp 1586364061
transform 1 0 36616 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_394
timestamp 1586364061
transform 1 0 37352 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_390
timestamp 1586364061
transform 1 0 36984 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_394
timestamp 1586364061
transform 1 0 37352 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_406
timestamp 1586364061
transform 1 0 38456 0 1 5984
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 1472 0 -1 7072
box -38 -48 1786 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l2_in_3_
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_40
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_55
timestamp 1586364061
transform 1 0 6164 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_59
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l2_in_2_
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_72
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_76
timestamp 1586364061
transform 1 0 8096 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _30_
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_83
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_87
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11316 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_110
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_4.mux_l2_in_3_
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_120
timestamp 1586364061
transform 1 0 12144 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_124
timestamp 1586364061
transform 1 0 12512 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_127
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_137
timestamp 1586364061
transform 1 0 13708 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_149
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_158
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15732 0 -1 7072
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_182
timestamp 1586364061
transform 1 0 17848 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21068 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_205
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 22264 0 -1 7072
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_8_219
timestamp 1586364061
transform 1 0 21252 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 24564 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_249
timestamp 1586364061
transform 1 0 24012 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_253
timestamp 1586364061
transform 1 0 24380 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_257
timestamp 1586364061
transform 1 0 24748 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l2_in_1_
timestamp 1586364061
transform 1 0 24840 0 -1 7072
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l2_in_2_
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_12.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 25852 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_267
timestamp 1586364061
transform 1 0 25668 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_271
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _24_
timestamp 1586364061
transform 1 0 28060 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 27508 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 27876 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_285
timestamp 1586364061
transform 1 0 27324 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_289
timestamp 1586364061
transform 1 0 27692 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_296
timestamp 1586364061
transform 1 0 28336 0 -1 7072
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_ipin_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 29072 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 28704 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_302
timestamp 1586364061
transform 1 0 28888 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_323
timestamp 1586364061
transform 1 0 30820 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_335
timestamp 1586364061
transform 1 0 31924 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l4_in_0_
timestamp 1586364061
transform 1 0 32752 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 32292 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 33764 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_341
timestamp 1586364061
transform 1 0 32476 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_353
timestamp 1586364061
transform 1 0 33580 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_357
timestamp 1586364061
transform 1 0 33948 0 -1 7072
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l1_in_0_
timestamp 1586364061
transform 1 0 34316 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 35328 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 35696 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_370
timestamp 1586364061
transform 1 0 35144 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_374
timestamp 1586364061
transform 1 0 35512 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l1_in_2_
timestamp 1586364061
transform 1 0 35880 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 36892 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_387
timestamp 1586364061
transform 1 0 36708 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_391
timestamp 1586364061
transform 1 0 37076 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 1786 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 3680 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_26
timestamp 1586364061
transform 1 0 3496 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_30
timestamp 1586364061
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_66
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_88
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_92
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_99
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_116
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_142
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_9_150
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_161
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_172
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_176
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19320 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18952 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 590 592
use scs8hd_fill_2  FILLER_9_192
timestamp 1586364061
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19504 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_209
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_11.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_11.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 24012 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_251
timestamp 1586364061
transform 1 0 24196 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 26496 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_274
timestamp 1586364061
transform 1 0 26312 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l2_in_3_
timestamp 1586364061
transform 1 0 27048 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 26864 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 28060 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_278
timestamp 1586364061
transform 1 0 26680 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_291
timestamp 1586364061
transform 1 0 27876 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_295
timestamp 1586364061
transform 1 0 28244 0 1 7072
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 28980 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 28612 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_301
timestamp 1586364061
transform 1 0 28796 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 32108 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_13.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 31740 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_325
timestamp 1586364061
transform 1 0 31004 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_335
timestamp 1586364061
transform 1 0 31924 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 32292 0 1 7072
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l1_in_1_
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 34592 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 34224 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_358
timestamp 1586364061
transform 1 0 34040 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_362
timestamp 1586364061
transform 1 0 34408 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_376
timestamp 1586364061
transform 1 0 35696 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l2_in_3_
timestamp 1586364061
transform 1 0 36432 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 35880 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 36248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_380
timestamp 1586364061
transform 1 0 36064 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_393
timestamp 1586364061
transform 1 0 37260 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_405
timestamp 1586364061
transform 1 0 38364 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _21_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_10
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l4_in_0_
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_42
timestamp 1586364061
transform 1 0 4968 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_55
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_59
timestamp 1586364061
transform 1 0 6532 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6900 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6716 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 8280 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_72
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_76
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 222 592
use scs8hd_conb_1  _29_
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_89
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_106
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_110
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13800 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_132
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_140
timestamp 1586364061
transform 1 0 13984 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 17296 0 -1 8160
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15732 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_168
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_172
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_195
timestamp 1586364061
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_203
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_199
timestamp 1586364061
transform 1 0 19412 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_207
timestamp 1586364061
transform 1 0 20148 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_211
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_conb_1  _23_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_218
timestamp 1586364061
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 22264 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 21344 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_222
timestamp 1586364061
transform 1 0 21528 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_226
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l3_in_0_
timestamp 1586364061
transform 1 0 24748 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 24564 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_249
timestamp 1586364061
transform 1 0 24012 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_253
timestamp 1586364061
transform 1 0 24380 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_11.mux_l4_in_0_
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 26036 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_266
timestamp 1586364061
transform 1 0 25576 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_270
timestamp 1586364061
transform 1 0 25944 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_273
timestamp 1586364061
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 27508 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 27876 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_285
timestamp 1586364061
transform 1 0 27324 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_289
timestamp 1586364061
transform 1 0 27692 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_293
timestamp 1586364061
transform 1 0 28060 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_297
timestamp 1586364061
transform 1 0 28428 0 -1 8160
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 28704 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 28520 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 30636 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_319
timestamp 1586364061
transform 1 0 30452 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_323
timestamp 1586364061
transform 1 0 30820 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_335
timestamp 1586364061
transform 1 0 31924 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_13.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 32936 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 32292 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 32660 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_341
timestamp 1586364061
transform 1 0 32476 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_345
timestamp 1586364061
transform 1 0 32844 0 -1 8160
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l2_in_2_
timestamp 1586364061
transform 1 0 35420 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 34868 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 35236 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_365
timestamp 1586364061
transform 1 0 34684 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_369
timestamp 1586364061
transform 1 0 35052 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 36432 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 36800 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_382
timestamp 1586364061
transform 1 0 36248 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_386
timestamp 1586364061
transform 1 0 36616 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_390
timestamp 1586364061
transform 1 0 36984 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_396
timestamp 1586364061
transform 1 0 37536 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_buf_2  _53_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 1786 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_35
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l3_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6900 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_72
timestamp 1586364061
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_76
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_100
timestamp 1586364061
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_104
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_108
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_127
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_131
timestamp 1586364061
transform 1 0 13156 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_5.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_151
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use scs8hd_conb_1  _32_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18676 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_182
timestamp 1586364061
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_187
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_206
timestamp 1586364061
transform 1 0 20056 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_210
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 22908 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_233
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l2_in_1_
timestamp 1586364061
transform 1 0 24196 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 24012 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_239
timestamp 1586364061
transform 1 0 23092 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l2_in_3_
timestamp 1586364061
transform 1 0 26036 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_260
timestamp 1586364061
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_264
timestamp 1586364061
transform 1 0 25392 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_268
timestamp 1586364061
transform 1 0 25760 0 1 8160
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l3_in_0_
timestamp 1586364061
transform 1 0 27600 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 27048 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 27416 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_280
timestamp 1586364061
transform 1 0 26864 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_284
timestamp 1586364061
transform 1 0 27232 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_297
timestamp 1586364061
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l4_in_0_
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 30268 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 28980 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 28612 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_301
timestamp 1586364061
transform 1 0 28796 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_315
timestamp 1586364061
transform 1 0 30084 0 1 8160
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_ipin_13.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 31004 0 1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 32108 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 31740 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 30820 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_319
timestamp 1586364061
transform 1 0 30452 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_331
timestamp 1586364061
transform 1 0 31556 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_335
timestamp 1586364061
transform 1 0 31924 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 32292 0 1 8160
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l3_in_1_
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 34224 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_358
timestamp 1586364061
transform 1 0 34040 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_362
timestamp 1586364061
transform 1 0 34408 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_376
timestamp 1586364061
transform 1 0 35696 0 1 8160
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_ipin_15.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 36432 0 1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 35880 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 36248 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 37168 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_380
timestamp 1586364061
transform 1 0 36064 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_390
timestamp 1586364061
transform 1 0 36984 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_394
timestamp 1586364061
transform 1 0 37352 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_406
timestamp 1586364061
transform 1 0 38456 0 1 8160
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_12
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_16
timestamp 1586364061
transform 1 0 2576 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_2  _46_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_20
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_24
timestamp 1586364061
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_28
timestamp 1586364061
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l2_in_3_
timestamp 1586364061
transform 1 0 5520 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_40
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_57
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_61
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_74
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_78
timestamp 1586364061
transform 1 0 8280 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l2_in_2_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_83
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_89
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_107
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_131
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_135
timestamp 1586364061
transform 1 0 13524 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_138
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_142
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_150
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l2_in_2_
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_193
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l3_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l4_in_0_
timestamp 1586364061
transform 1 0 22908 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 22264 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 22724 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_228
timestamp 1586364061
transform 1 0 22080 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_232
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l3_in_0_
timestamp 1586364061
transform 1 0 24472 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_246
timestamp 1586364061
transform 1 0 23736 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_250
timestamp 1586364061
transform 1 0 24104 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_253
timestamp 1586364061
transform 1 0 24380 0 -1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l3_in_1_
timestamp 1586364061
transform 1 0 26588 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 25484 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 26036 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_267
timestamp 1586364061
transform 1 0 25668 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_273
timestamp 1586364061
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 27600 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 27968 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 28336 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_286
timestamp 1586364061
transform 1 0 27416 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_290
timestamp 1586364061
transform 1 0 27784 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_294
timestamp 1586364061
transform 1 0 28152 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 29532 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 29256 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 28888 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_298
timestamp 1586364061
transform 1 0 28520 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_304
timestamp 1586364061
transform 1 0 29072 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_308
timestamp 1586364061
transform 1 0 29440 0 -1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_328
timestamp 1586364061
transform 1 0 31280 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_337
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_13.mux_l3_in_0_
timestamp 1586364061
transform 1 0 32568 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 33580 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 32384 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 33948 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_351
timestamp 1586364061
transform 1 0 33396 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_355
timestamp 1586364061
transform 1 0 33764 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 34132 0 -1 9248
box -38 -48 1786 592
use scs8hd_conb_1  _26_
timestamp 1586364061
transform 1 0 36616 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 36064 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 36432 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_378
timestamp 1586364061
transform 1 0 35880 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_382
timestamp 1586364061
transform 1 0 36248 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_389
timestamp 1586364061
transform 1 0 36892 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_buf_4  mux_bottom_ipin_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 590 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l3_in_1_
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_18
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_14_26
timestamp 1586364061
transform 1 0 3496 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_22
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_38
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_1.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 4508 0 -1 10336
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_13_42
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _47_
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_54
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_50
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_58
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_66
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_60
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_87
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_83
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_90
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_99
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_90
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l2_in_3_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 11316 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l3_in_0_
timestamp 1586364061
transform 1 0 11500 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_126
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_122
timestamp 1586364061
transform 1 0 12328 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_134
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_130
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_146
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_142
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_150
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 16008 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_173
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_177
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_164
timestamp 1586364061
transform 1 0 16192 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_185
timestamp 1586364061
transform 1 0 18124 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_188
timestamp 1586364061
transform 1 0 18400 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_181
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_193
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l1_in_2_
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_204
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_200
timestamp 1586364061
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l2_in_3_
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_210
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 21068 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 21252 0 -1 10336
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_221
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_234
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_14_238
timestamp 1586364061
transform 1 0 23000 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_244
timestamp 1586364061
transform 1 0 23552 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 23368 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 23736 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l2_in_2_
timestamp 1586364061
transform 1 0 23736 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_252
timestamp 1586364061
transform 1 0 24288 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_248
timestamp 1586364061
transform 1 0 23920 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_255
timestamp 1586364061
transform 1 0 24564 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 24472 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l2_in_0_
timestamp 1586364061
transform 1 0 24656 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_265
timestamp 1586364061
transform 1 0 25484 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_259
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 25668 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_273
timestamp 1586364061
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_269
timestamp 1586364061
transform 1 0 25852 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 26036 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_conb_1  _28_
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 25300 0 1 9248
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_14_283
timestamp 1586364061
transform 1 0 27140 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_279
timestamp 1586364061
transform 1 0 26772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_287
timestamp 1586364061
transform 1 0 27508 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_282
timestamp 1586364061
transform 1 0 27048 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 27324 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 26956 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_295
timestamp 1586364061
transform 1 0 28244 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_291
timestamp 1586364061
transform 1 0 27876 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 28060 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 27692 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l2_in_0_
timestamp 1586364061
transform 1 0 27692 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_6  FILLER_14_298
timestamp 1586364061
transform 1 0 28520 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_3  FILLER_13_306
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_301
timestamp 1586364061
transform 1 0 28796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 29072 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 28612 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 28980 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l1_in_0_
timestamp 1586364061
transform 1 0 29256 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_315
timestamp 1586364061
transform 1 0 30084 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_15.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 30268 0 -1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_15.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 29532 0 1 9248
box -38 -48 1786 592
use scs8hd_buf_2  _70_
timestamp 1586364061
transform 1 0 32108 0 1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 31924 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_328
timestamp 1586364061
transform 1 0 31280 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_334
timestamp 1586364061
transform 1 0 31832 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_319
timestamp 1586364061
transform 1 0 30452 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_331
timestamp 1586364061
transform 1 0 31556 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_335
timestamp 1586364061
transform 1 0 31924 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 32660 0 -1 10336
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l1_in_0_
timestamp 1586364061
transform 1 0 33212 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 33028 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__70__A
timestamp 1586364061
transform 1 0 32660 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 32476 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_341
timestamp 1586364061
transform 1 0 32476 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_345
timestamp 1586364061
transform 1 0 32844 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_366
timestamp 1586364061
transform 1 0 34776 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_362
timestamp 1586364061
transform 1 0 34408 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_362
timestamp 1586364061
transform 1 0 34408 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_358
timestamp 1586364061
transform 1 0 34040 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 34224 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_369
timestamp 1586364061
transform 1 0 35052 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_376
timestamp 1586364061
transform 1 0 35696 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 34868 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l2_in_0_
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_ipin_14.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 35144 0 -1 10336
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_13_380
timestamp 1586364061
transform 1 0 36064 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_14.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 35880 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 36248 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _73_
timestamp 1586364061
transform 1 0 36432 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_389
timestamp 1586364061
transform 1 0 36892 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_388
timestamp 1586364061
transform 1 0 36800 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 37076 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__73__A
timestamp 1586364061
transform 1 0 36984 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_393
timestamp 1586364061
transform 1 0 37260 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_392
timestamp 1586364061
transform 1 0 37168 0 1 9248
box -38 -48 406 592
use scs8hd_conb_1  _27_
timestamp 1586364061
transform 1 0 37536 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_399
timestamp 1586364061
transform 1 0 37812 0 1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_conb_1  _22_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_6
timestamp 1586364061
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_10
timestamp 1586364061
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_23
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _45_
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_44
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_52
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_56
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_77
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_80
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_84
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_107
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l4_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 1786 592
use scs8hd_conb_1  _17_
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_168
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_172
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_176
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_188
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_181
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_15_216
timestamp 1586364061
transform 1 0 20976 0 1 10336
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 21712 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_222
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_233
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_237
timestamp 1586364061
transform 1 0 22908 0 1 10336
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_8.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_241
timestamp 1586364061
transform 1 0 23276 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_10.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_10.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_258
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 27140 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 28244 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_281
timestamp 1586364061
transform 1 0 26956 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_285
timestamp 1586364061
transform 1 0 27324 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_293
timestamp 1586364061
transform 1 0 28060 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_297
timestamp 1586364061
transform 1 0 28428 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 28980 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 28612 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_301
timestamp 1586364061
transform 1 0 28796 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _65_
timestamp 1586364061
transform 1 0 32108 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__61__A
timestamp 1586364061
transform 1 0 31188 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 31924 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 31556 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_325
timestamp 1586364061
transform 1 0 31004 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_329
timestamp 1586364061
transform 1 0 31372 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_333
timestamp 1586364061
transform 1 0 31740 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l2_in_1_
timestamp 1586364061
transform 1 0 33212 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 33028 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 32660 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_341
timestamp 1586364061
transform 1 0 32476 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_345
timestamp 1586364061
transform 1 0 32844 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l2_in_2_
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 34592 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 34224 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_358
timestamp 1586364061
transform 1 0 34040 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_362
timestamp 1586364061
transform 1 0 34408 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_376
timestamp 1586364061
transform 1 0 35696 0 1 10336
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l3_in_1_
timestamp 1586364061
transform 1 0 36432 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__72__A
timestamp 1586364061
transform 1 0 36156 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 37444 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_380
timestamp 1586364061
transform 1 0 36064 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_383
timestamp 1586364061
transform 1 0 36340 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_393
timestamp 1586364061
transform 1 0 37260 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_397
timestamp 1586364061
transform 1 0 37628 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_405
timestamp 1586364061
transform 1 0 38364 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _50_
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_45
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_53
timestamp 1586364061
transform 1 0 5980 0 -1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_61
timestamp 1586364061
transform 1 0 6716 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_76
timestamp 1586364061
transform 1 0 8096 0 -1 11424
box -38 -48 406 592
use scs8hd_conb_1  _33_
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_89
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11960 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_114
timestamp 1586364061
transform 1 0 11592 0 -1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_6.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_16_120
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_140
timestamp 1586364061
transform 1 0 13984 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_148
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 590 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l4_in_0_
timestamp 1586364061
transform 1 0 16008 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_171
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_175
timestamp 1586364061
transform 1 0 17204 0 -1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_ipin_7.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 17572 0 -1 11424
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_16_198
timestamp 1586364061
transform 1 0 19320 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 21160 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 21344 0 -1 11424
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_ipin_8.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 23644 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 23276 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_243
timestamp 1586364061
transform 1 0 23460 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 25760 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 26128 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_266
timestamp 1586364061
transform 1 0 25576 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_270
timestamp 1586364061
transform 1 0 25944 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 28428 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_295
timestamp 1586364061
transform 1 0 28244 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_15.mux_l2_in_1_
timestamp 1586364061
transform 1 0 28980 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 29992 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 28796 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_299
timestamp 1586364061
transform 1 0 28612 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_312
timestamp 1586364061
transform 1 0 29808 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_316
timestamp 1586364061
transform 1 0 30176 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _61_
timestamp 1586364061
transform 1 0 30912 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 30360 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 30728 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_320
timestamp 1586364061
transform 1 0 30544 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_328
timestamp 1586364061
transform 1 0 31280 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_337
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l3_in_0_
timestamp 1586364061
transform 1 0 32844 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 33856 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 32660 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 32292 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_341
timestamp 1586364061
transform 1 0 32476 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_354
timestamp 1586364061
transform 1 0 33672 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l2_in_3_
timestamp 1586364061
transform 1 0 34592 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 34408 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 35604 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_358
timestamp 1586364061
transform 1 0 34040 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_373
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _72_
timestamp 1586364061
transform 1 0 36156 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 36708 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_377
timestamp 1586364061
transform 1 0 35788 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_385
timestamp 1586364061
transform 1 0 36524 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_389
timestamp 1586364061
transform 1 0 36892 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_2  _44_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_24
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_28
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _42_
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_41
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_45
timestamp 1586364061
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_ipin_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_68
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_72
timestamp 1586364061
transform 1 0 7728 0 1 11424
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l2_in_2_
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_84
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_96
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_108
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_116
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_120
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l2_in_2_
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_146
timestamp 1586364061
transform 1 0 14536 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_158
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l3_in_1_
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_162
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l2_in_3_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l4_in_0_
timestamp 1586364061
transform 1 0 20792 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 20608 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 19872 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_202
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_206
timestamp 1586364061
transform 1 0 20056 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_210
timestamp 1586364061
transform 1 0 20424 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _18_
timestamp 1586364061
transform 1 0 22356 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 22172 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_223
timestamp 1586364061
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_227
timestamp 1586364061
transform 1 0 21988 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_234
timestamp 1586364061
transform 1 0 22632 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_238
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23920 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_242
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 25484 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 25300 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_261
timestamp 1586364061
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _19_
timestamp 1586364061
transform 1 0 28152 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 27692 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_284
timestamp 1586364061
transform 1 0 27232 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_288
timestamp 1586364061
transform 1 0 27600 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_291
timestamp 1586364061
transform 1 0 27876 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_297
timestamp 1586364061
transform 1 0 28428 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _62_
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__62__A
timestamp 1586364061
transform 1 0 29808 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__60__A
timestamp 1586364061
transform 1 0 30176 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 28612 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 28980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_301
timestamp 1586364061
transform 1 0 28796 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_310
timestamp 1586364061
transform 1 0 29624 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_314
timestamp 1586364061
transform 1 0 29992 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_ipin_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 30360 0 1 11424
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_17_337
timestamp 1586364061
transform 1 0 32108 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_14.mux_l4_in_0_
timestamp 1586364061
transform 1 0 33120 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__58__A
timestamp 1586364061
transform 1 0 32660 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 32292 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_341
timestamp 1586364061
transform 1 0 32476 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_345
timestamp 1586364061
transform 1 0 32844 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_357
timestamp 1586364061
transform 1 0 33948 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _71_
timestamp 1586364061
transform 1 0 35420 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__68__A
timestamp 1586364061
transform 1 0 35236 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 34592 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 34132 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_361
timestamp 1586364061
transform 1 0 34316 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 406 592
use scs8hd_buf_2  _67_
timestamp 1586364061
transform 1 0 36524 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__71__A
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__67__A
timestamp 1586364061
transform 1 0 37076 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__66__A
timestamp 1586364061
transform 1 0 36340 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_377
timestamp 1586364061
transform 1 0 35788 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_381
timestamp 1586364061
transform 1 0 36156 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_389
timestamp 1586364061
transform 1 0 36892 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_393
timestamp 1586364061
transform 1 0 37260 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_405
timestamp 1586364061
transform 1 0 38364 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_9
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _43_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3496 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_20
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_24
timestamp 1586364061
transform 1 0 3312 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_28
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 406 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_18_40
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_18_48
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 774 592
use scs8hd_buf_2  _35_
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_60
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_72
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_ipin_6.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11960 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 130 592
use scs8hd_buf_4  mux_bottom_ipin_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_127
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_131
timestamp 1586364061
transform 1 0 13156 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_151
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l3_in_0_
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_162
timestamp 1586364061
transform 1 0 16008 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_175
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 774 592
use scs8hd_buf_4  mux_bottom_ipin_7.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 17940 0 -1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_189
timestamp 1586364061
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_193
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 590 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l3_in_1_
timestamp 1586364061
transform 1 0 21160 0 -1 12512
box -38 -48 866 592
use scs8hd_buf_4  mux_bottom_ipin_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19504 0 -1 12512
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_199
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_3  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l2_in_2_
timestamp 1586364061
transform 1 0 22724 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 24656 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23920 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_244
timestamp 1586364061
transform 1 0 23552 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_250
timestamp 1586364061
transform 1 0 24104 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_254
timestamp 1586364061
transform 1 0 24472 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 24840 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 25944 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_267
timestamp 1586364061
transform 1 0 25668 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_272
timestamp 1586364061
transform 1 0 26128 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 27692 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 27508 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 26864 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_282
timestamp 1586364061
transform 1 0 27048 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_286
timestamp 1586364061
transform 1 0 27416 0 -1 12512
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l3_in_1_
timestamp 1586364061
transform 1 0 29256 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 30268 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 29072 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 28704 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_298
timestamp 1586364061
transform 1 0 28520 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_302
timestamp 1586364061
transform 1 0 28888 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_315
timestamp 1586364061
transform 1 0 30084 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _60_
timestamp 1586364061
transform 1 0 30912 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 31464 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 30636 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_319
timestamp 1586364061
transform 1 0 30452 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_323
timestamp 1586364061
transform 1 0 30820 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_328
timestamp 1586364061
transform 1 0 31280 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_332
timestamp 1586364061
transform 1 0 31648 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_6  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 590 592
use scs8hd_buf_2  _58_
timestamp 1586364061
transform 1 0 32660 0 -1 12512
box -38 -48 406 592
use scs8hd_buf_4  mux_bottom_ipin_14.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 33764 0 -1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 33580 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_347
timestamp 1586364061
transform 1 0 33028 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_351
timestamp 1586364061
transform 1 0 33396 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _68_
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_361
timestamp 1586364061
transform 1 0 34316 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_2  _66_
timestamp 1586364061
transform 1 0 36524 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_18_377
timestamp 1586364061
transform 1 0 35788 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_18_389
timestamp 1586364061
transform 1 0 36892 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_8
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_16
timestamp 1586364061
transform 1 0 2576 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_1.mux_l2_in_3_
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_28
timestamp 1586364061
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_20
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_25
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_21
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_36
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_35
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_4  mux_bottom_ipin_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 590 592
use scs8hd_buf_2  _40_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 406 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 406 592
use scs8hd_buf_4  mux_bottom_ipin_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_43
timestamp 1586364061
transform 1 0 5060 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_46
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_48
timestamp 1586364061
transform 1 0 5520 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_20_60
timestamp 1586364061
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_66
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_buf_2  _36_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use scs8hd_buf_2  _34_
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_70
timestamp 1586364061
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_79
timestamp 1586364061
transform 1 0 8372 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_67
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_buf_4  mux_bottom_ipin_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_94
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_94
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_103
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_19_119
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use scs8hd_buf_4  mux_bottom_ipin_6.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13340 0 1 12512
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_144
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_139
timestamp 1586364061
transform 1 0 13892 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_5.mux_l4_in_0_
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_150
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_157
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_7.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_162
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_164
timestamp 1586364061
transform 1 0 16192 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 20516 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_213
timestamp 1586364061
transform 1 0 20700 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_217
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_226
timestamp 1586364061
transform 1 0 21896 0 -1 13600
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_8.mux_l2_in_3_
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 866 592
use scs8hd_buf_4  mux_bottom_ipin_10.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21344 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_234
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_230
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_11.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_ipin_11.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22632 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_6  FILLER_19_238
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 590 592
use scs8hd_decap_8  FILLER_20_240
timestamp 1586364061
transform 1 0 23184 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_253
timestamp 1586364061
transform 1 0 24380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_250
timestamp 1586364061
transform 1 0 24104 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23920 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_257
timestamp 1586364061
transform 1 0 24748 0 -1 13600
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_ipin_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_266
timestamp 1586364061
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_262
timestamp 1586364061
transform 1 0 25208 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 24932 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 25392 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_10.mux_l1_in_0_
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_275
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_270
timestamp 1586364061
transform 1 0 25944 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 26588 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 25760 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l4_in_0_
timestamp 1586364061
transform 1 0 25944 0 1 12512
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 27508 0 1 12512
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 26864 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 26772 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 27324 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 26956 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_279
timestamp 1586364061
transform 1 0 26772 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_283
timestamp 1586364061
transform 1 0 27140 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_296
timestamp 1586364061
transform 1 0 28336 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_289
timestamp 1586364061
transform 1 0 27692 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_307
timestamp 1586364061
transform 1 0 29348 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_301
timestamp 1586364061
transform 1 0 28796 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_301
timestamp 1586364061
transform 1 0 28796 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 28612 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 28980 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 29440 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l2_in_3_
timestamp 1586364061
transform 1 0 29532 0 1 12512
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l2_in_2_
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_6  FILLER_20_320
timestamp 1586364061
transform 1 0 30544 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_322
timestamp 1586364061
transform 1 0 30728 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_318
timestamp 1586364061
transform 1 0 30360 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 31096 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 30912 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 30544 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_9.mux_l1_in_2_
timestamp 1586364061
transform 1 0 31096 0 1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_333
timestamp 1586364061
transform 1 0 31740 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_328
timestamp 1586364061
transform 1 0 31280 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_335
timestamp 1586364061
transform 1 0 31924 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__59__A
timestamp 1586364061
transform 1 0 32108 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _59_
timestamp 1586364061
transform 1 0 31372 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_6  FILLER_20_342
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_339
timestamp 1586364061
transform 1 0 32292 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_12.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 32476 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_4  mux_bottom_ipin_12.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 32660 0 1 12512
box -38 -48 590 592
use scs8hd_decap_8  FILLER_20_352
timestamp 1586364061
transform 1 0 33488 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_6  FILLER_19_353
timestamp 1586364061
transform 1 0 33580 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_349
timestamp 1586364061
transform 1 0 33212 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__A
timestamp 1586364061
transform 1 0 33396 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _57_
timestamp 1586364061
transform 1 0 33120 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_364
timestamp 1586364061
transform 1 0 34592 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_19_362
timestamp 1586364061
transform 1 0 34408 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_359
timestamp 1586364061
transform 1 0 34132 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 34224 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _56_
timestamp 1586364061
transform 1 0 34224 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 35236 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_buf_2  _63_
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 406 592
use scs8hd_buf_2  _55_
timestamp 1586364061
transform 1 0 35420 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_377
timestamp 1586364061
transform 1 0 35788 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_381
timestamp 1586364061
transform 1 0 36156 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_377
timestamp 1586364061
transform 1 0 35788 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 36340 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__A
timestamp 1586364061
transform 1 0 35972 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _64_
timestamp 1586364061
transform 1 0 36524 0 1 12512
box -38 -48 406 592
use scs8hd_buf_2  _54_
timestamp 1586364061
transform 1 0 36524 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_389
timestamp 1586364061
transform 1 0 36892 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 37076 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_389
timestamp 1586364061
transform 1 0 36892 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_393
timestamp 1586364061
transform 1 0 37260 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_405
timestamp 1586364061
transform 1 0 38364 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_401
timestamp 1586364061
transform 1 0 37996 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_404
timestamp 1586364061
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal2 s 4986 0 5042 480 6 bottom_grid_pin_0_
port 0 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 ccff_head
port 1 nsew default input
rlabel metal2 s 24950 0 25006 480 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 0 144 480 264 6 chanx_left_in[0]
port 3 nsew default input
rlabel metal3 s 0 4088 480 4208 6 chanx_left_in[10]
port 4 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[11]
port 5 nsew default input
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[12]
port 6 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[13]
port 7 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[14]
port 8 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[15]
port 9 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[16]
port 10 nsew default input
rlabel metal3 s 0 6944 480 7064 6 chanx_left_in[17]
port 11 nsew default input
rlabel metal3 s 0 7352 480 7472 6 chanx_left_in[18]
port 12 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[19]
port 13 nsew default input
rlabel metal3 s 0 416 480 536 6 chanx_left_in[1]
port 14 nsew default input
rlabel metal3 s 0 824 480 944 6 chanx_left_in[2]
port 15 nsew default input
rlabel metal3 s 0 1232 480 1352 6 chanx_left_in[3]
port 16 nsew default input
rlabel metal3 s 0 1640 480 1760 6 chanx_left_in[4]
port 17 nsew default input
rlabel metal3 s 0 2048 480 2168 6 chanx_left_in[5]
port 18 nsew default input
rlabel metal3 s 0 2456 480 2576 6 chanx_left_in[6]
port 19 nsew default input
rlabel metal3 s 0 2864 480 2984 6 chanx_left_in[7]
port 20 nsew default input
rlabel metal3 s 0 3272 480 3392 6 chanx_left_in[8]
port 21 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[9]
port 22 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_out[0]
port 23 nsew default tristate
rlabel metal3 s 0 12112 480 12232 6 chanx_left_out[10]
port 24 nsew default tristate
rlabel metal3 s 0 12520 480 12640 6 chanx_left_out[11]
port 25 nsew default tristate
rlabel metal3 s 0 12928 480 13048 6 chanx_left_out[12]
port 26 nsew default tristate
rlabel metal3 s 0 13336 480 13456 6 chanx_left_out[13]
port 27 nsew default tristate
rlabel metal3 s 0 13744 480 13864 6 chanx_left_out[14]
port 28 nsew default tristate
rlabel metal3 s 0 14152 480 14272 6 chanx_left_out[15]
port 29 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[16]
port 30 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[17]
port 31 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[18]
port 32 nsew default tristate
rlabel metal3 s 0 15784 480 15904 6 chanx_left_out[19]
port 33 nsew default tristate
rlabel metal3 s 0 8440 480 8560 6 chanx_left_out[1]
port 34 nsew default tristate
rlabel metal3 s 0 8848 480 8968 6 chanx_left_out[2]
port 35 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[3]
port 36 nsew default tristate
rlabel metal3 s 0 9664 480 9784 6 chanx_left_out[4]
port 37 nsew default tristate
rlabel metal3 s 0 10072 480 10192 6 chanx_left_out[5]
port 38 nsew default tristate
rlabel metal3 s 0 10480 480 10600 6 chanx_left_out[6]
port 39 nsew default tristate
rlabel metal3 s 0 10888 480 11008 6 chanx_left_out[7]
port 40 nsew default tristate
rlabel metal3 s 0 11296 480 11416 6 chanx_left_out[8]
port 41 nsew default tristate
rlabel metal3 s 0 11704 480 11824 6 chanx_left_out[9]
port 42 nsew default tristate
rlabel metal3 s 39520 144 40000 264 6 chanx_right_in[0]
port 43 nsew default input
rlabel metal3 s 39520 4088 40000 4208 6 chanx_right_in[10]
port 44 nsew default input
rlabel metal3 s 39520 4496 40000 4616 6 chanx_right_in[11]
port 45 nsew default input
rlabel metal3 s 39520 4904 40000 5024 6 chanx_right_in[12]
port 46 nsew default input
rlabel metal3 s 39520 5312 40000 5432 6 chanx_right_in[13]
port 47 nsew default input
rlabel metal3 s 39520 5720 40000 5840 6 chanx_right_in[14]
port 48 nsew default input
rlabel metal3 s 39520 6128 40000 6248 6 chanx_right_in[15]
port 49 nsew default input
rlabel metal3 s 39520 6536 40000 6656 6 chanx_right_in[16]
port 50 nsew default input
rlabel metal3 s 39520 6944 40000 7064 6 chanx_right_in[17]
port 51 nsew default input
rlabel metal3 s 39520 7352 40000 7472 6 chanx_right_in[18]
port 52 nsew default input
rlabel metal3 s 39520 7760 40000 7880 6 chanx_right_in[19]
port 53 nsew default input
rlabel metal3 s 39520 416 40000 536 6 chanx_right_in[1]
port 54 nsew default input
rlabel metal3 s 39520 824 40000 944 6 chanx_right_in[2]
port 55 nsew default input
rlabel metal3 s 39520 1232 40000 1352 6 chanx_right_in[3]
port 56 nsew default input
rlabel metal3 s 39520 1640 40000 1760 6 chanx_right_in[4]
port 57 nsew default input
rlabel metal3 s 39520 2048 40000 2168 6 chanx_right_in[5]
port 58 nsew default input
rlabel metal3 s 39520 2456 40000 2576 6 chanx_right_in[6]
port 59 nsew default input
rlabel metal3 s 39520 2864 40000 2984 6 chanx_right_in[7]
port 60 nsew default input
rlabel metal3 s 39520 3272 40000 3392 6 chanx_right_in[8]
port 61 nsew default input
rlabel metal3 s 39520 3680 40000 3800 6 chanx_right_in[9]
port 62 nsew default input
rlabel metal3 s 39520 8168 40000 8288 6 chanx_right_out[0]
port 63 nsew default tristate
rlabel metal3 s 39520 12112 40000 12232 6 chanx_right_out[10]
port 64 nsew default tristate
rlabel metal3 s 39520 12520 40000 12640 6 chanx_right_out[11]
port 65 nsew default tristate
rlabel metal3 s 39520 12928 40000 13048 6 chanx_right_out[12]
port 66 nsew default tristate
rlabel metal3 s 39520 13336 40000 13456 6 chanx_right_out[13]
port 67 nsew default tristate
rlabel metal3 s 39520 13744 40000 13864 6 chanx_right_out[14]
port 68 nsew default tristate
rlabel metal3 s 39520 14152 40000 14272 6 chanx_right_out[15]
port 69 nsew default tristate
rlabel metal3 s 39520 14560 40000 14680 6 chanx_right_out[16]
port 70 nsew default tristate
rlabel metal3 s 39520 14968 40000 15088 6 chanx_right_out[17]
port 71 nsew default tristate
rlabel metal3 s 39520 15376 40000 15496 6 chanx_right_out[18]
port 72 nsew default tristate
rlabel metal3 s 39520 15784 40000 15904 6 chanx_right_out[19]
port 73 nsew default tristate
rlabel metal3 s 39520 8440 40000 8560 6 chanx_right_out[1]
port 74 nsew default tristate
rlabel metal3 s 39520 8848 40000 8968 6 chanx_right_out[2]
port 75 nsew default tristate
rlabel metal3 s 39520 9256 40000 9376 6 chanx_right_out[3]
port 76 nsew default tristate
rlabel metal3 s 39520 9664 40000 9784 6 chanx_right_out[4]
port 77 nsew default tristate
rlabel metal3 s 39520 10072 40000 10192 6 chanx_right_out[5]
port 78 nsew default tristate
rlabel metal3 s 39520 10480 40000 10600 6 chanx_right_out[6]
port 79 nsew default tristate
rlabel metal3 s 39520 10888 40000 11008 6 chanx_right_out[7]
port 80 nsew default tristate
rlabel metal3 s 39520 11296 40000 11416 6 chanx_right_out[8]
port 81 nsew default tristate
rlabel metal3 s 39520 11704 40000 11824 6 chanx_right_out[9]
port 82 nsew default tristate
rlabel metal2 s 34978 0 35034 480 6 prog_clk
port 83 nsew default input
rlabel metal2 s 1214 15520 1270 16000 6 top_grid_pin_16_
port 84 nsew default tristate
rlabel metal2 s 3698 15520 3754 16000 6 top_grid_pin_17_
port 85 nsew default tristate
rlabel metal2 s 6182 15520 6238 16000 6 top_grid_pin_18_
port 86 nsew default tristate
rlabel metal2 s 8666 15520 8722 16000 6 top_grid_pin_19_
port 87 nsew default tristate
rlabel metal2 s 11150 15520 11206 16000 6 top_grid_pin_20_
port 88 nsew default tristate
rlabel metal2 s 13634 15520 13690 16000 6 top_grid_pin_21_
port 89 nsew default tristate
rlabel metal2 s 16210 15520 16266 16000 6 top_grid_pin_22_
port 90 nsew default tristate
rlabel metal2 s 18694 15520 18750 16000 6 top_grid_pin_23_
port 91 nsew default tristate
rlabel metal2 s 21178 15520 21234 16000 6 top_grid_pin_24_
port 92 nsew default tristate
rlabel metal2 s 23662 15520 23718 16000 6 top_grid_pin_25_
port 93 nsew default tristate
rlabel metal2 s 26146 15520 26202 16000 6 top_grid_pin_26_
port 94 nsew default tristate
rlabel metal2 s 28722 15520 28778 16000 6 top_grid_pin_27_
port 95 nsew default tristate
rlabel metal2 s 31206 15520 31262 16000 6 top_grid_pin_28_
port 96 nsew default tristate
rlabel metal2 s 33690 15520 33746 16000 6 top_grid_pin_29_
port 97 nsew default tristate
rlabel metal2 s 36174 15520 36230 16000 6 top_grid_pin_30_
port 98 nsew default tristate
rlabel metal2 s 38658 15520 38714 16000 6 top_grid_pin_31_
port 99 nsew default tristate
rlabel metal4 s 7611 2128 7931 13648 6 vpwr
port 100 nsew default input
rlabel metal4 s 14277 2128 14597 13648 6 vgnd
port 101 nsew default input
<< properties >>
string FIXED_BBOX 0 0 40000 16000
<< end >>
