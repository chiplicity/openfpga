VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_clb
  CLASS BLOCK ;
  FOREIGN grid_clb ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 85.720 250.000 86.320 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 101.360 250.000 101.960 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 117.000 250.000 117.600 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 132.640 250.000 133.240 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 148.280 250.000 148.880 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 163.920 250.000 164.520 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 179.560 250.000 180.160 ;
    END
  END address[6]
  PIN address[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 195.200 250.000 195.800 ;
    END
  END address[7]
  PIN address[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 210.840 250.000 211.440 ;
    END
  END address[8]
  PIN address[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 226.480 250.000 227.080 ;
    END
  END address[9]
  PIN bottom_width_0_height_0__pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 2.400 ;
    END
  END bottom_width_0_height_0__pin_10_
  PIN bottom_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 2.400 ;
    END
  END bottom_width_0_height_0__pin_14_
  PIN bottom_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 2.400 ;
    END
  END bottom_width_0_height_0__pin_2_
  PIN bottom_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 2.400 ;
    END
  END bottom_width_0_height_0__pin_6_
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 2.400 ;
    END
  END clk
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 242.120 250.000 242.720 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 70.080 250.000 70.680 ;
    END
  END enable
  PIN left_width_0_height_0__pin_11_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 2.400 208.720 ;
    END
  END left_width_0_height_0__pin_11_
  PIN left_width_0_height_0__pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 2.400 42.120 ;
    END
  END left_width_0_height_0__pin_3_
  PIN left_width_0_height_0__pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 2.400 125.080 ;
    END
  END left_width_0_height_0__pin_7_
  PIN reset
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 2.400 ;
    END
  END reset
  PIN right_width_0_height_0__pin_13_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 54.440 250.000 55.040 ;
    END
  END right_width_0_height_0__pin_13_
  PIN right_width_0_height_0__pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 7.520 250.000 8.120 ;
    END
  END right_width_0_height_0__pin_1_
  PIN right_width_0_height_0__pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 23.160 250.000 23.760 ;
    END
  END right_width_0_height_0__pin_5_
  PIN right_width_0_height_0__pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 38.800 250.000 39.400 ;
    END
  END right_width_0_height_0__pin_9_
  PIN set
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 2.400 ;
    END
  END set
  PIN top_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 247.600 31.190 250.000 ;
    END
  END top_width_0_height_0__pin_0_
  PIN top_width_0_height_0__pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 218.130 247.600 218.410 250.000 ;
    END
  END top_width_0_height_0__pin_12_
  PIN top_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.010 247.600 93.290 250.000 ;
    END
  END top_width_0_height_0__pin_4_
  PIN top_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 155.570 247.600 155.850 250.000 ;
    END
  END top_width_0_height_0__pin_8_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 236.880 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 236.880 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 244.260 236.725 ;
      LAYER met1 ;
        RECT 5.520 10.640 247.870 236.880 ;
      LAYER met2 ;
        RECT 17.850 247.320 30.630 247.930 ;
        RECT 31.470 247.320 92.730 247.930 ;
        RECT 93.570 247.320 155.290 247.930 ;
        RECT 156.130 247.320 217.850 247.930 ;
        RECT 218.690 247.320 247.850 247.930 ;
        RECT 17.850 2.680 247.850 247.320 ;
        RECT 18.130 0.270 52.710 2.680 ;
        RECT 53.550 0.270 88.590 2.680 ;
        RECT 89.430 0.270 124.010 2.680 ;
        RECT 124.850 0.270 159.890 2.680 ;
        RECT 160.730 0.270 195.310 2.680 ;
        RECT 196.150 0.270 231.190 2.680 ;
        RECT 232.030 0.270 247.850 2.680 ;
      LAYER met3 ;
        RECT 0.270 241.720 247.200 242.585 ;
        RECT 0.270 227.480 248.130 241.720 ;
        RECT 0.270 226.080 247.200 227.480 ;
        RECT 0.270 211.840 248.130 226.080 ;
        RECT 0.270 210.440 247.200 211.840 ;
        RECT 0.270 209.120 248.130 210.440 ;
        RECT 2.800 207.720 248.130 209.120 ;
        RECT 0.270 196.200 248.130 207.720 ;
        RECT 0.270 194.800 247.200 196.200 ;
        RECT 0.270 180.560 248.130 194.800 ;
        RECT 0.270 179.160 247.200 180.560 ;
        RECT 0.270 164.920 248.130 179.160 ;
        RECT 0.270 163.520 247.200 164.920 ;
        RECT 0.270 149.280 248.130 163.520 ;
        RECT 0.270 147.880 247.200 149.280 ;
        RECT 0.270 133.640 248.130 147.880 ;
        RECT 0.270 132.240 247.200 133.640 ;
        RECT 0.270 125.480 248.130 132.240 ;
        RECT 2.800 124.080 248.130 125.480 ;
        RECT 0.270 118.000 248.130 124.080 ;
        RECT 0.270 116.600 247.200 118.000 ;
        RECT 0.270 102.360 248.130 116.600 ;
        RECT 0.270 100.960 247.200 102.360 ;
        RECT 0.270 86.720 248.130 100.960 ;
        RECT 0.270 85.320 247.200 86.720 ;
        RECT 0.270 71.080 248.130 85.320 ;
        RECT 0.270 69.680 247.200 71.080 ;
        RECT 0.270 55.440 248.130 69.680 ;
        RECT 0.270 54.040 247.200 55.440 ;
        RECT 0.270 42.520 248.130 54.040 ;
        RECT 2.800 41.120 248.130 42.520 ;
        RECT 0.270 39.800 248.130 41.120 ;
        RECT 0.270 38.400 247.200 39.800 ;
        RECT 0.270 24.160 248.130 38.400 ;
        RECT 0.270 22.760 247.200 24.160 ;
        RECT 0.270 8.520 248.130 22.760 ;
        RECT 0.270 8.120 247.200 8.520 ;
      LAYER met4 ;
        RECT 0.295 10.640 20.640 236.880 ;
        RECT 23.040 10.640 97.440 236.880 ;
        RECT 99.840 10.640 248.105 236.880 ;
  END
END grid_clb
END LIBRARY

