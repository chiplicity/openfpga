* NGSPICE file created from sb_3__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

.subckt sb_3__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_13_ bottom_right_grid_pin_11_ bottom_right_grid_pin_13_
+ bottom_right_grid_pin_15_ bottom_right_grid_pin_1_ bottom_right_grid_pin_3_ bottom_right_grid_pin_5_
+ bottom_right_grid_pin_7_ bottom_right_grid_pin_9_ chanx_left_in[0] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ left_bottom_grid_pin_12_ left_top_grid_pin_10_ top_left_grid_pin_13_ top_right_grid_pin_11_
+ top_right_grid_pin_13_ top_right_grid_pin_15_ top_right_grid_pin_1_ top_right_grid_pin_3_
+ top_right_grid_pin_5_ top_right_grid_pin_7_ top_right_grid_pin_9_ vpwr vgnd
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_137 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_1_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _218_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_18_225 vgnd vpwr scs8hd_fill_1
XFILLER_18_269 vgnd vpwr scs8hd_decap_6
XANTENNA__124__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vpwr vgnd scs8hd_fill_2
XFILLER_24_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _208_/HI mem_bottom_track_17.LATCH_2_.latch/Q
+ mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _189_/A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
X_200_ _200_/A _200_/Y vgnd vpwr scs8hd_inv_8
X_131_ _131_/A _132_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_97 vpwr vgnd scs8hd_fill_2
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XANTENNA__110__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__119__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_77 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_17.LATCH_2_.latch data_in mem_bottom_track_17.LATCH_2_.latch/Q _160_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _235_/A vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_97 vgnd vpwr scs8hd_decap_3
XFILLER_34_85 vgnd vpwr scs8hd_decap_6
XFILLER_11_253 vpwr vgnd scs8hd_fill_2
XFILLER_11_275 vpwr vgnd scs8hd_fill_2
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
X_114_ _134_/A address[4] _134_/C _114_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _203_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_6_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__121__B _120_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XANTENNA__222__A _222_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _216_/HI _193_/Y mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[7] mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_23 vgnd vpwr scs8hd_decap_8
XANTENNA__116__B _177_/C vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_194 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_0_230 vgnd vpwr scs8hd_decap_3
XFILLER_0_241 vgnd vpwr scs8hd_decap_6
XFILLER_31_145 vpwr vgnd scs8hd_fill_2
XFILLER_31_134 vpwr vgnd scs8hd_fill_2
XFILLER_16_186 vgnd vpwr scs8hd_decap_6
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A _127_/A vgnd vpwr scs8hd_diode_2
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _208_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_112 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_149 vgnd vpwr scs8hd_decap_4
XFILLER_13_178 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[0] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_171 vgnd vpwr scs8hd_decap_12
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _210_/HI _190_/Y mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_259 vpwr vgnd scs8hd_fill_2
XFILLER_10_148 vgnd vpwr scs8hd_decap_4
XFILLER_12_22 vgnd vpwr scs8hd_decap_4
XFILLER_12_55 vgnd vpwr scs8hd_decap_3
XANTENNA__230__A _230_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _205_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_204 vpwr vgnd scs8hd_fill_2
Xmux_left_track_13.tap_buf4_0_.scs8hd_inv_1 mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _224_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _140_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_15_207 vpwr vgnd scs8hd_fill_2
XFILLER_23_32 vpwr vgnd scs8hd_fill_2
X_130_ _140_/A _132_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_87 vgnd vpwr scs8hd_fill_1
XANTENNA__225__A _225_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_144 vpwr vgnd scs8hd_fill_2
XANTENNA__119__B _120_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_58 vgnd vpwr scs8hd_decap_4
XFILLER_0_69 vpwr vgnd scs8hd_fill_2
XFILLER_9_12 vpwr vgnd scs8hd_fill_2
XANTENNA__135__A _134_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_34 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_232 vgnd vpwr scs8hd_decap_12
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_5.tap_buf4_0_.scs8hd_inv_1 mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _228_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _196_/Y vgnd vpwr
+ scs8hd_diode_2
X_113_ address[3] _134_/A vgnd vpwr scs8hd_inv_8
XFILLER_11_210 vgnd vpwr scs8hd_decap_4
XFILLER_11_221 vpwr vgnd scs8hd_fill_2
XFILLER_11_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_20_11 vgnd vpwr scs8hd_fill_1
XFILLER_20_99 vgnd vpwr scs8hd_decap_4
XFILLER_6_35 vgnd vpwr scs8hd_decap_6
Xmux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _192_/A mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__132__B _132_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_184 vgnd vpwr scs8hd_fill_1
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
Xmem_left_track_5.LATCH_1_.latch data_in _193_/A _174_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_187 vpwr vgnd scs8hd_fill_2
XFILLER_25_121 vgnd vpwr scs8hd_fill_1
XANTENNA__233__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[7] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vpwr vgnd scs8hd_fill_2
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_9 vpwr vgnd scs8hd_fill_2
XFILLER_26_32 vpwr vgnd scs8hd_fill_2
XFILLER_26_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__228__A _228_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_157 vpwr vgnd scs8hd_fill_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _231_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A _128_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _196_/Y mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_8_194 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_127 vpwr vgnd scs8hd_fill_2
XFILLER_12_89 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _198_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_6 vpwr vgnd scs8hd_fill_2
XFILLER_37_31 vgnd vpwr scs8hd_decap_12
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_271 vgnd vpwr scs8hd_decap_4
XFILLER_5_153 vpwr vgnd scs8hd_fill_2
XFILLER_5_197 vpwr vgnd scs8hd_fill_2
XFILLER_38_6 vgnd vpwr scs8hd_decap_12
XANTENNA__140__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
XFILLER_23_11 vpwr vgnd scs8hd_fill_2
XANTENNA__241__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_15 vgnd vpwr scs8hd_decap_4
X_189_ _189_/A _189_/Y vgnd vpwr scs8hd_inv_8
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A _140_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_11 vpwr vgnd scs8hd_fill_2
XFILLER_18_22 vgnd vpwr scs8hd_fill_1
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_88 vpwr vgnd scs8hd_fill_2
XANTENNA__236__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
X_112_ _099_/A _133_/A _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__A _155_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_5_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_23 vgnd vpwr scs8hd_decap_4
XFILLER_20_45 vpwr vgnd scs8hd_fill_2
XFILLER_20_89 vgnd vpwr scs8hd_decap_3
XFILLER_29_65 vpwr vgnd scs8hd_fill_2
XFILLER_28_174 vgnd vpwr scs8hd_decap_12
XFILLER_28_163 vgnd vpwr scs8hd_decap_3
XFILLER_6_14 vgnd vpwr scs8hd_decap_3
XFILLER_3_262 vgnd vpwr scs8hd_decap_12
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_177 vpwr vgnd scs8hd_fill_2
XFILLER_15_12 vpwr vgnd scs8hd_fill_2
XFILLER_15_34 vpwr vgnd scs8hd_fill_2
XFILLER_31_55 vgnd vpwr scs8hd_decap_3
XFILLER_31_44 vgnd vpwr scs8hd_decap_4
XFILLER_31_22 vgnd vpwr scs8hd_decap_3
XFILLER_31_11 vgnd vpwr scs8hd_decap_4
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_258 vpwr vgnd scs8hd_fill_2
XFILLER_39_225 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_125 vgnd vpwr scs8hd_decap_6
XFILLER_22_169 vpwr vgnd scs8hd_fill_2
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_136 vgnd vpwr scs8hd_decap_4
XANTENNA__244__A _244_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_59 vpwr vgnd scs8hd_fill_2
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_4_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__138__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_151 vpwr vgnd scs8hd_fill_2
XFILLER_12_180 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.INVTX1_1_.scs8hd_inv_1 chany_top_in[8] mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_68 vpwr vgnd scs8hd_fill_2
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_43 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__239__A _239_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_121 vgnd vpwr scs8hd_fill_1
Xmem_left_track_15.LATCH_0_.latch data_in _204_/A _186_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_132 vpwr vgnd scs8hd_fill_2
XFILLER_5_176 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _112_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__149__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_track_17.LATCH_3_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_220 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB _184_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_168 vgnd vpwr scs8hd_decap_3
XFILLER_2_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_0_49 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
X_188_ _172_/A _163_/A _166_/C _167_/A _188_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__151__B _153_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_190 vgnd vpwr scs8hd_decap_12
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A bottom_right_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
X_111_ _110_/X _133_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_245 vgnd vpwr scs8hd_decap_8
XANTENNA__162__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_81 vpwr vgnd scs8hd_fill_2
XFILLER_4_208 vgnd vpwr scs8hd_decap_6
XFILLER_29_11 vpwr vgnd scs8hd_fill_2
XFILLER_20_79 vpwr vgnd scs8hd_fill_2
XFILLER_29_88 vpwr vgnd scs8hd_fill_2
XFILLER_29_55 vgnd vpwr scs8hd_decap_4
XFILLER_28_186 vgnd vpwr scs8hd_decap_12
XFILLER_28_120 vgnd vpwr scs8hd_decap_6
XANTENNA__247__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_3_241 vgnd vpwr scs8hd_decap_3
XFILLER_3_274 vgnd vpwr scs8hd_decap_3
XFILLER_20_7 vpwr vgnd scs8hd_fill_2
XFILLER_19_131 vpwr vgnd scs8hd_fill_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__157__A _128_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_2_.latch data_in mem_bottom_track_1.LATCH_2_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_25_156 vpwr vgnd scs8hd_fill_2
XFILLER_25_145 vpwr vgnd scs8hd_fill_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_16_134 vgnd vpwr scs8hd_decap_4
XFILLER_16_145 vgnd vpwr scs8hd_decap_8
XFILLER_31_126 vpwr vgnd scs8hd_fill_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB _181_/Y vgnd vpwr scs8hd_diode_2
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _191_/Y mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _206_/Y vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_1.LATCH_1_.latch data_in _189_/A _166_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_67 vpwr vgnd scs8hd_fill_2
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__154__B _153_/B vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_107 vpwr vgnd scs8hd_fill_2
XFILLER_12_14 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_55 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_218 vgnd vpwr scs8hd_decap_4
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_37_88 vpwr vgnd scs8hd_fill_2
XFILLER_26_251 vgnd vpwr scs8hd_decap_4
XANTENNA__149__B _153_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_240 vgnd vpwr scs8hd_decap_4
XFILLER_17_273 vgnd vpwr scs8hd_decap_4
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_70 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_79 vpwr vgnd scs8hd_fill_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_23_24 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_136 vgnd vpwr scs8hd_decap_6
XFILLER_2_125 vpwr vgnd scs8hd_fill_2
Xmux_left_track_13.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[6] mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_39 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _172_/A _163_/A _166_/C _165_/A _187_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_1_180 vgnd vpwr scs8hd_decap_3
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_9.INVTX1_3_.scs8hd_inv_1 bottom_right_grid_pin_9_ mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_56 vgnd vpwr scs8hd_fill_1
X_110_ address[1] address[2] address[0] _110_/X vgnd vpwr scs8hd_or3_4
XFILLER_7_206 vpwr vgnd scs8hd_fill_2
X_239_ _239_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__B _162_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_34 vpwr vgnd scs8hd_fill_2
XFILLER_28_198 vgnd vpwr scs8hd_decap_12
XFILLER_3_253 vpwr vgnd scs8hd_fill_2
XFILLER_34_124 vgnd vpwr scs8hd_decap_12
XFILLER_19_198 vpwr vgnd scs8hd_fill_2
XANTENNA__157__B _162_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _211_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__173__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_25_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _178_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XFILLER_31_79 vpwr vgnd scs8hd_fill_2
XFILLER_31_149 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_102 vpwr vgnd scs8hd_fill_2
XFILLER_16_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__168__A _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_190 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _190_/A mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_26_57 vgnd vpwr scs8hd_fill_1
XFILLER_13_116 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_171 vpwr vgnd scs8hd_fill_2
XFILLER_21_160 vpwr vgnd scs8hd_fill_2
XFILLER_3_39 vgnd vpwr scs8hd_fill_1
XFILLER_16_90 vpwr vgnd scs8hd_fill_2
XANTENNA__170__B _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _195_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_208 vgnd vpwr scs8hd_decap_6
Xmem_top_track_8.LATCH_1_.latch data_in mem_top_track_8.LATCH_1_.latch/Q _122_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__181__A _180_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _194_/Y mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__091__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_2_148 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_16 vpwr vgnd scs8hd_fill_2
XFILLER_9_49 vpwr vgnd scs8hd_fill_2
X_186_ _180_/X _163_/A _177_/C _167_/A _186_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__176__A _172_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_247 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_11.LATCH_0_.latch data_in _200_/A _182_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_1.INVTX1_6_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_25 vpwr vgnd scs8hd_fill_2
XFILLER_34_68 vpwr vgnd scs8hd_fill_2
XANTENNA__086__A _107_/C vgnd vpwr scs8hd_diode_2
XFILLER_11_214 vgnd vpwr scs8hd_fill_1
XFILLER_11_225 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_5_.scs8hd_inv_1 chanx_left_in[2] mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_238_ chany_top_in[0] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
X_169_ _169_/A _163_/X _169_/C _165_/X _169_/Y vgnd vpwr scs8hd_nor4_4
Xmux_left_track_11.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[5] mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_251 vgnd vpwr scs8hd_decap_12
XFILLER_37_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_133 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_81 vpwr vgnd scs8hd_fill_2
XFILLER_19_90 vgnd vpwr scs8hd_decap_3
XFILLER_19_144 vpwr vgnd scs8hd_fill_2
XFILLER_19_155 vpwr vgnd scs8hd_fill_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_34_136 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_9.LATCH_3_.latch data_in mem_bottom_track_9.LATCH_3_.latch/Q _151_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _197_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_213 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_158 vgnd vpwr scs8hd_fill_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_206 vpwr vgnd scs8hd_fill_2
XANTENNA__168__B _163_/X vgnd vpwr scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__184__A _180_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_47 vpwr vgnd scs8hd_fill_2
XANTENNA__094__A _094_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_143 vpwr vgnd scs8hd_fill_2
XFILLER_8_154 vpwr vgnd scs8hd_fill_2
XANTENNA__170__C _169_/C vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _172_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_12_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__089__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_113 vpwr vgnd scs8hd_fill_2
XFILLER_5_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__181__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_4_190 vgnd vpwr scs8hd_decap_3
XFILLER_23_245 vgnd vpwr scs8hd_decap_12
XFILLER_3_7 vgnd vpwr scs8hd_decap_12
XANTENNA__091__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_19 vgnd vpwr scs8hd_fill_1
XFILLER_14_201 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
X_185_ _180_/X _163_/A _177_/C _165_/A _185_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_1_160 vpwr vgnd scs8hd_fill_2
XFILLER_20_215 vpwr vgnd scs8hd_fill_2
XFILLER_20_204 vpwr vgnd scs8hd_fill_2
XANTENNA__176__B _175_/B vgnd vpwr scs8hd_diode_2
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_259 vgnd vpwr scs8hd_decap_12
XFILLER_18_59 vpwr vgnd scs8hd_fill_2
XFILLER_11_237 vgnd vpwr scs8hd_decap_6
XFILLER_11_259 vpwr vgnd scs8hd_fill_2
X_237_ chany_top_in[1] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_24_80 vpwr vgnd scs8hd_fill_2
X_168_ _169_/A _163_/X _166_/C _167_/X _168_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
X_099_ _099_/A _119_/A _099_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XFILLER_1_62 vpwr vgnd scs8hd_fill_2
XANTENNA__187__A _172_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_27 vgnd vpwr scs8hd_fill_1
XFILLER_20_49 vgnd vpwr scs8hd_decap_3
XFILLER_29_69 vpwr vgnd scs8hd_fill_2
XFILLER_28_145 vgnd vpwr scs8hd_decap_8
XANTENNA__097__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_148 vgnd vpwr scs8hd_decap_4
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_25_126 vpwr vgnd scs8hd_fill_2
XFILLER_15_16 vgnd vpwr scs8hd_decap_3
XFILLER_0_247 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_17.LATCH_3_.latch data_in mem_bottom_track_17.LATCH_3_.latch/Q _159_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_118 vgnd vpwr scs8hd_decap_4
XFILLER_24_192 vgnd vpwr scs8hd_decap_12
XFILLER_24_181 vpwr vgnd scs8hd_fill_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_229 vgnd vpwr scs8hd_decap_12
XFILLER_39_218 vgnd vpwr scs8hd_decap_3
Xmux_left_track_5.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__168__C _166_/C vgnd vpwr scs8hd_diode_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__184__B _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_251 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_184 vpwr vgnd scs8hd_fill_2
XFILLER_3_19 vgnd vpwr scs8hd_decap_12
XFILLER_29_262 vgnd vpwr scs8hd_decap_12
XFILLER_8_122 vpwr vgnd scs8hd_fill_2
XANTENNA__170__D _167_/X vgnd vpwr scs8hd_diode_2
XANTENNA__179__B _175_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XANTENNA__195__A _195_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_3.INVTX1_2_.scs8hd_inv_1_A left_bottom_grid_pin_12_ vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _189_/Y mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__089__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_136 vpwr vgnd scs8hd_fill_2
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XANTENNA__181__C _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_213 vgnd vpwr scs8hd_decap_4
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
XFILLER_23_224 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_106 vgnd vpwr scs8hd_decap_4
XANTENNA__091__C _134_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_29 vgnd vpwr scs8hd_decap_3
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
XFILLER_14_224 vgnd vpwr scs8hd_decap_12
X_184_ _180_/X _163_/X _184_/C _167_/A _184_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_29_7 vpwr vgnd scs8hd_fill_2
XFILLER_1_172 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_5_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__176__C _177_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_167_ _167_/A _167_/X vgnd vpwr scs8hd_buf_1
X_236_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
X_098_ _098_/A _119_/A vgnd vpwr scs8hd_buf_1
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
XFILLER_1_85 vpwr vgnd scs8hd_fill_2
XANTENNA__187__B _163_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _205_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_15 vgnd vpwr scs8hd_decap_8
XFILLER_28_168 vgnd vpwr scs8hd_decap_3
XFILLER_28_102 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__097__B _084_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
XFILLER_35_91 vpwr vgnd scs8hd_fill_2
XFILLER_35_80 vpwr vgnd scs8hd_fill_2
X_219_ _219_/HI _219_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_149 vpwr vgnd scs8hd_fill_2
XFILLER_15_28 vgnd vpwr scs8hd_decap_4
XFILLER_31_27 vpwr vgnd scs8hd_fill_2
XFILLER_0_237 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_108 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _220_/HI mem_top_track_16.LATCH_2_.latch/Q
+ mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_108 vgnd vpwr scs8hd_decap_6
XANTENNA__168__D _167_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XANTENNA__184__C _184_/C vgnd vpwr scs8hd_diode_2
XFILLER_30_163 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_84 vpwr vgnd scs8hd_fill_2
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XFILLER_26_27 vpwr vgnd scs8hd_fill_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_274 vgnd vpwr scs8hd_decap_3
XFILLER_16_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_167 vpwr vgnd scs8hd_fill_2
XFILLER_12_141 vgnd vpwr scs8hd_fill_1
XFILLER_12_163 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A top_right_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__179__C _166_/C vgnd vpwr scs8hd_diode_2
XFILLER_12_18 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_26_200 vgnd vpwr scs8hd_decap_12
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_104 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _230_/A vgnd vpwr scs8hd_inv_1
XANTENNA__181__D _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_74 vgnd vpwr scs8hd_fill_1
XFILLER_4_30 vgnd vpwr scs8hd_fill_1
XFILLER_23_236 vgnd vpwr scs8hd_decap_8
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XFILLER_23_28 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_236 vgnd vpwr scs8hd_decap_8
XFILLER_14_247 vgnd vpwr scs8hd_decap_8
XFILLER_13_83 vpwr vgnd scs8hd_fill_2
XFILLER_13_94 vpwr vgnd scs8hd_fill_2
X_183_ _180_/X _163_/X _184_/C _165_/A _183_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_1_184 vgnd vpwr scs8hd_decap_4
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XANTENNA__176__D _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_217 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 top_right_grid_pin_9_ mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_6 vpwr vgnd scs8hd_fill_2
XFILLER_24_93 vgnd vpwr scs8hd_decap_3
X_235_ _235_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_40_81 vgnd vpwr scs8hd_decap_8
Xmux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _192_/Y mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_166_ _169_/A _163_/X _166_/C _165_/X _166_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_097_ address[1] _084_/Y _167_/A _098_/A vgnd vpwr scs8hd_or3_4
XFILLER_37_147 vgnd vpwr scs8hd_decap_12
XFILLER_1_31 vpwr vgnd scs8hd_fill_2
XFILLER_1_42 vgnd vpwr scs8hd_decap_4
XFILLER_1_53 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _198_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__187__C _166_/C vgnd vpwr scs8hd_diode_2
XFILLER_29_38 vpwr vgnd scs8hd_fill_2
XANTENNA__097__C _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_60 vgnd vpwr scs8hd_fill_1
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
X_218_ _218_/HI _218_/LO vgnd vpwr scs8hd_conb_1
X_149_ _128_/A _153_/B _149_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _212_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_117 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_191 vpwr vgnd scs8hd_fill_2
XFILLER_0_249 vgnd vpwr scs8hd_decap_12
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_106 vgnd vpwr scs8hd_decap_4
XFILLER_16_117 vpwr vgnd scs8hd_fill_2
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_94 vgnd vpwr scs8hd_decap_3
XFILLER_21_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_161 vgnd vpwr scs8hd_decap_3
XANTENNA__184__D _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_175 vgnd vpwr scs8hd_decap_12
XFILLER_7_30 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _209_/HI mem_bottom_track_9.LATCH_2_.latch/Q
+ mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_197 vpwr vgnd scs8hd_fill_2
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_253 vpwr vgnd scs8hd_fill_2
XFILLER_29_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_102 vgnd vpwr scs8hd_decap_3
XFILLER_12_120 vgnd vpwr scs8hd_decap_3
XFILLER_32_93 vpwr vgnd scs8hd_fill_2
XFILLER_12_186 vpwr vgnd scs8hd_fill_2
XFILLER_12_197 vgnd vpwr scs8hd_decap_4
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XANTENNA__179__D _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_212 vpwr vgnd scs8hd_fill_2
XFILLER_5_149 vpwr vgnd scs8hd_fill_2
XFILLER_17_212 vgnd vpwr scs8hd_decap_3
XFILLER_17_223 vpwr vgnd scs8hd_fill_2
XFILLER_17_245 vgnd vpwr scs8hd_decap_4
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_97 vpwr vgnd scs8hd_fill_2
XFILLER_4_53 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_119 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_3_.scs8hd_inv_1 bottom_right_grid_pin_7_ mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_182_ _180_/X address[5] _169_/C _167_/X _182_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_14_259 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_13_ mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_18 vgnd vpwr scs8hd_decap_4
XFILLER_18_29 vpwr vgnd scs8hd_fill_2
X_165_ _165_/A _165_/X vgnd vpwr scs8hd_buf_1
X_234_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
XFILLER_34_7 vgnd vpwr scs8hd_decap_12
X_096_ address[0] _167_/A vgnd vpwr scs8hd_buf_1
XFILLER_37_159 vgnd vpwr scs8hd_decap_12
XFILLER_37_104 vgnd vpwr scs8hd_decap_12
XFILLER_1_10 vpwr vgnd scs8hd_fill_2
XFILLER_1_98 vpwr vgnd scs8hd_fill_2
XANTENNA__187__D _165_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _109_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_left_track_15.LATCH_1_.latch data_in _203_/A _185_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_126 vgnd vpwr scs8hd_fill_1
XFILLER_3_258 vpwr vgnd scs8hd_fill_2
XFILLER_10_41 vpwr vgnd scs8hd_fill_2
XFILLER_10_85 vpwr vgnd scs8hd_fill_2
XFILLER_19_126 vgnd vpwr scs8hd_decap_3
XFILLER_19_148 vpwr vgnd scs8hd_fill_2
XFILLER_19_159 vgnd vpwr scs8hd_decap_3
XFILLER_34_107 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd vpwr
+ scs8hd_diode_2
X_148_ _147_/X _153_/B vgnd vpwr scs8hd_buf_1
X_217_ _217_/HI _217_/LO vgnd vpwr scs8hd_conb_1
XFILLER_18_181 vgnd vpwr scs8hd_decap_4
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XFILLER_31_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB _175_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_162 vpwr vgnd scs8hd_fill_2
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _099_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_187 vgnd vpwr scs8hd_decap_12
XFILLER_30_132 vpwr vgnd scs8hd_fill_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_151 vgnd vpwr scs8hd_decap_8
XFILLER_15_184 vgnd vpwr scs8hd_decap_4
XFILLER_7_42 vpwr vgnd scs8hd_fill_2
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_154 vgnd vpwr scs8hd_decap_4
XFILLER_29_232 vgnd vpwr scs8hd_decap_12
XFILLER_32_72 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_147 vpwr vgnd scs8hd_fill_2
XANTENNA__103__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_4_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_180 vgnd vpwr scs8hd_fill_1
XFILLER_5_117 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_3_.latch data_in mem_bottom_track_1.LATCH_3_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_257 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_205 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A bottom_right_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
X_181_ _180_/X address[5] _169_/C _165_/X _181_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_1_131 vpwr vgnd scs8hd_fill_2
XFILLER_38_93 vgnd vpwr scs8hd_decap_3
XFILLER_1_164 vpwr vgnd scs8hd_fill_2
XFILLER_20_219 vgnd vpwr scs8hd_decap_4
XFILLER_20_208 vgnd vpwr scs8hd_decap_6
Xmux_top_track_0.INVTX1_5_.scs8hd_inv_1 chanx_left_in[0] mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
X_233_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_24_84 vpwr vgnd scs8hd_fill_2
X_164_ _126_/B _166_/C vgnd vpwr scs8hd_buf_1
XFILLER_6_201 vgnd vpwr scs8hd_decap_12
XFILLER_10_230 vgnd vpwr scs8hd_decap_12
XFILLER_10_274 vgnd vpwr scs8hd_fill_1
X_095_ _128_/A _099_/A _095_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_7 vpwr vgnd scs8hd_fill_2
XFILLER_37_116 vgnd vpwr scs8hd_decap_6
XFILLER_1_66 vgnd vpwr scs8hd_decap_4
XANTENNA__111__A _110_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_64 vgnd vpwr scs8hd_decap_3
XFILLER_27_160 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_62 vgnd vpwr scs8hd_decap_4
XFILLER_19_95 vpwr vgnd scs8hd_fill_2
X_216_ _216_/HI _216_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__106__A _099_/A vgnd vpwr scs8hd_diode_2
X_147_ _169_/A _163_/A _184_/C _147_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_141 vgnd vpwr scs8hd_decap_12
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XFILLER_24_141 vpwr vgnd scs8hd_fill_2
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_199 vgnd vpwr scs8hd_decap_12
XFILLER_30_100 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_65 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _205_/A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_126 vpwr vgnd scs8hd_fill_2
XFILLER_12_100 vgnd vpwr scs8hd_decap_3
XFILLER_12_144 vpwr vgnd scs8hd_fill_2
XFILLER_16_74 vpwr vgnd scs8hd_fill_2
XFILLER_32_84 vgnd vpwr scs8hd_decap_8
XANTENNA__103__B _140_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_84 vgnd vpwr scs8hd_decap_8
XFILLER_17_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_66 vpwr vgnd scs8hd_fill_2
XANTENNA__114__A _134_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_180_ _172_/A _180_/X vgnd vpwr scs8hd_buf_1
XFILLER_22_261 vgnd vpwr scs8hd_decap_12
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_176 vpwr vgnd scs8hd_fill_2
XFILLER_1_143 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_243 vgnd vpwr scs8hd_fill_1
XANTENNA__109__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_19 vgnd vpwr scs8hd_decap_12
X_232_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
X_163_ _163_/A _163_/X vgnd vpwr scs8hd_buf_1
XFILLER_6_213 vgnd vpwr scs8hd_fill_1
XFILLER_10_242 vgnd vpwr scs8hd_decap_12
X_094_ _094_/A _099_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _221_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _188_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_2_.latch data_in mem_top_track_8.LATCH_2_.latch/Q _121_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_205 vgnd vpwr scs8hd_decap_12
XFILLER_10_10 vpwr vgnd scs8hd_fill_2
XFILLER_10_76 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
Xmux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_150 vgnd vpwr scs8hd_decap_4
XFILLER_19_52 vpwr vgnd scs8hd_fill_2
XFILLER_35_95 vgnd vpwr scs8hd_decap_4
XFILLER_35_84 vpwr vgnd scs8hd_fill_2
XFILLER_35_62 vgnd vpwr scs8hd_decap_6
X_215_ _215_/HI _215_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
X_146_ _155_/B _163_/A vgnd vpwr scs8hd_buf_1
XANTENNA__122__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA__106__B _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_153 vgnd vpwr scs8hd_decap_12
XFILLER_18_161 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _190_/Y mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_24_175 vgnd vpwr scs8hd_decap_4
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_left_track_11.LATCH_1_.latch data_in _199_/A _181_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_120 vpwr vgnd scs8hd_fill_2
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XFILLER_30_145 vgnd vpwr scs8hd_decap_8
XFILLER_7_88 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _116_/X vgnd vpwr scs8hd_diode_2
X_129_ _119_/A _132_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_21_123 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_8
XFILLER_16_53 vpwr vgnd scs8hd_fill_2
XFILLER_16_86 vpwr vgnd scs8hd_fill_2
XFILLER_12_167 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_19 vgnd vpwr scs8hd_decap_12
XFILLER_26_259 vgnd vpwr scs8hd_decap_12
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB _185_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_108 vgnd vpwr scs8hd_decap_3
Xmem_bottom_track_9.LATCH_4_.latch data_in mem_bottom_track_9.LATCH_4_.latch/Q _150_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _200_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
Xmem_left_track_7.LATCH_0_.latch data_in _196_/A _177_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__114__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA__130__A _140_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_196 vgnd vpwr scs8hd_decap_12
XFILLER_4_185 vgnd vpwr scs8hd_decap_3
XFILLER_4_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _197_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_273 vpwr vgnd scs8hd_fill_2
XFILLER_13_43 vpwr vgnd scs8hd_fill_2
XFILLER_13_98 vgnd vpwr scs8hd_decap_3
XANTENNA__109__B _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA__125__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_6_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_170 vgnd vpwr scs8hd_fill_1
X_231_ _231_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
X_162_ _133_/A _162_/B _162_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_30 vgnd vpwr scs8hd_fill_1
XFILLER_10_254 vgnd vpwr scs8hd_decap_12
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
X_093_ _136_/A _184_/C _094_/A vgnd vpwr scs8hd_or2_4
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_35 vpwr vgnd scs8hd_fill_2
XFILLER_28_129 vgnd vpwr scs8hd_decap_4
XFILLER_28_107 vpwr vgnd scs8hd_fill_2
XFILLER_3_217 vgnd vpwr scs8hd_decap_12
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XFILLER_27_173 vpwr vgnd scs8hd_fill_2
XFILLER_19_86 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_214_ _214_/HI _214_/LO vgnd vpwr scs8hd_conb_1
X_145_ address[5] _155_/B vgnd vpwr scs8hd_inv_8
XANTENNA__122__B _120_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_165 vgnd vpwr scs8hd_decap_12
XFILLER_33_121 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _213_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_209 vpwr vgnd scs8hd_fill_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_6
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__223__A _223_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_113 vgnd vpwr scs8hd_decap_12
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_132 vpwr vgnd scs8hd_fill_2
XFILLER_30_157 vgnd vpwr scs8hd_decap_4
XANTENNA__133__A _133_/A vgnd vpwr scs8hd_diode_2
X_128_ _128_/A _132_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_34 vgnd vpwr scs8hd_decap_4
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_190 vgnd vpwr scs8hd_decap_3
XFILLER_8_139 vpwr vgnd scs8hd_fill_2
XANTENNA__128__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_172 vpwr vgnd scs8hd_fill_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_17_249 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
XFILLER_27_97 vpwr vgnd scs8hd_fill_2
XANTENNA__114__C _134_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_track_17.LATCH_4_.latch data_in mem_bottom_track_17.LATCH_4_.latch/Q _158_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__130__B _132_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_271 vgnd vpwr scs8hd_decap_4
XFILLER_13_22 vpwr vgnd scs8hd_fill_2
XFILLER_38_30 vgnd vpwr scs8hd_fill_1
XANTENNA__231__A _231_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _189_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_223 vgnd vpwr scs8hd_decap_12
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XANTENNA__125__B _134_/B vgnd vpwr scs8hd_diode_2
XANTENNA__141__A _131_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_182 vgnd vpwr scs8hd_fill_1
X_230_ _230_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_24_32 vgnd vpwr scs8hd_decap_4
XFILLER_24_21 vgnd vpwr scs8hd_decap_4
XANTENNA__226__A _226_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
X_161_ _161_/A _162_/B _161_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_266 vgnd vpwr scs8hd_decap_8
X_092_ _092_/A _184_/C vgnd vpwr scs8hd_buf_1
XFILLER_1_14 vgnd vpwr scs8hd_decap_12
XANTENNA__136__A _136_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_229 vgnd vpwr scs8hd_decap_12
XFILLER_10_23 vpwr vgnd scs8hd_fill_2
XFILLER_10_45 vpwr vgnd scs8hd_fill_2
XFILLER_10_89 vgnd vpwr scs8hd_decap_3
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_144_ address[6] _169_/A vgnd vpwr scs8hd_buf_1
Xmux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _221_/HI mem_top_track_8.LATCH_2_.latch/Q
+ mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_213_ _213_/HI _213_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_177 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_111 vgnd vpwr scs8hd_decap_4
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_99 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA__133__B _132_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_13 vpwr vgnd scs8hd_fill_2
XFILLER_7_46 vpwr vgnd scs8hd_fill_2
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
X_127_ _127_/A _132_/B vgnd vpwr scs8hd_buf_1
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _239_/A vgnd vpwr scs8hd_inv_1
Xmux_top_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[4] mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
XFILLER_29_258 vpwr vgnd scs8hd_fill_2
XFILLER_8_107 vgnd vpwr scs8hd_decap_6
XFILLER_12_125 vgnd vpwr scs8hd_decap_3
XFILLER_32_32 vgnd vpwr scs8hd_decap_3
XANTENNA__234__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__144__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _132_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_140 vpwr vgnd scs8hd_fill_2
XFILLER_7_184 vpwr vgnd scs8hd_fill_2
XFILLER_7_195 vpwr vgnd scs8hd_fill_2
XFILLER_34_250 vgnd vpwr scs8hd_decap_12
XFILLER_26_239 vgnd vpwr scs8hd_decap_12
XANTENNA__229__A _229_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_65 vpwr vgnd scs8hd_fill_2
XFILLER_27_32 vgnd vpwr scs8hd_decap_4
XFILLER_17_217 vgnd vpwr scs8hd_decap_4
XFILLER_4_154 vgnd vpwr scs8hd_fill_1
XFILLER_4_143 vpwr vgnd scs8hd_fill_2
XFILLER_4_132 vgnd vpwr scs8hd_decap_8
XFILLER_4_110 vgnd vpwr scs8hd_decap_8
XFILLER_4_36 vgnd vpwr scs8hd_decap_4
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XFILLER_23_209 vpwr vgnd scs8hd_fill_2
XANTENNA__139__A _119_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _203_/A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_13_12 vpwr vgnd scs8hd_fill_2
XFILLER_1_102 vpwr vgnd scs8hd_fill_2
XFILLER_1_113 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_135 vgnd vpwr scs8hd_decap_4
XANTENNA__125__C _134_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_235 vgnd vpwr scs8hd_decap_8
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
Xmem_left_track_3.LATCH_0_.latch data_in _192_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__141__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_190 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_150 vpwr vgnd scs8hd_fill_2
XFILLER_5_90 vgnd vpwr scs8hd_fill_1
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_88 vpwr vgnd scs8hd_fill_2
XFILLER_24_55 vpwr vgnd scs8hd_fill_2
X_091_ address[3] address[4] _134_/C _092_/A vgnd vpwr scs8hd_or3_4
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
X_160_ _131_/A _162_/B _160_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_76 vpwr vgnd scs8hd_fill_2
XANTENNA__242__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_1_26 vpwr vgnd scs8hd_fill_2
XFILLER_1_48 vpwr vgnd scs8hd_fill_2
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XANTENNA__136__B _169_/C vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_131 vpwr vgnd scs8hd_fill_2
XFILLER_19_44 vpwr vgnd scs8hd_fill_2
XFILLER_19_66 vgnd vpwr scs8hd_fill_1
XFILLER_19_99 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XANTENNA__237__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
X_212_ _212_/HI _212_/LO vgnd vpwr scs8hd_conb_1
X_143_ _133_/A _140_/B _143_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_7 vpwr vgnd scs8hd_fill_2
XANTENNA__147__A _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_2_91 vgnd vpwr scs8hd_fill_1
XFILLER_24_145 vgnd vpwr scs8hd_decap_8
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_45 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_101 vpwr vgnd scs8hd_fill_2
XFILLER_15_112 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_69 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[8] mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_126_ _136_/A _126_/B _127_/A vgnd vpwr scs8hd_or2_4
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_30_6 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_137 vpwr vgnd scs8hd_fill_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_12_137 vgnd vpwr scs8hd_decap_4
XFILLER_12_148 vgnd vpwr scs8hd_decap_3
XFILLER_16_78 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_170 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__160__A _131_/A vgnd vpwr scs8hd_diode_2
X_109_ _099_/A _161_/A _109_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_262 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_11 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XANTENNA__245__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_166 vgnd vpwr scs8hd_decap_8
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XANTENNA__155__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__139__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_13_79 vpwr vgnd scs8hd_fill_2
XFILLER_1_147 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_210 vgnd vpwr scs8hd_decap_4
XFILLER_13_221 vpwr vgnd scs8hd_fill_2
XFILLER_13_243 vgnd vpwr scs8hd_fill_1
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_184 vgnd vpwr scs8hd_decap_12
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
X_090_ enable _134_/C vgnd vpwr scs8hd_inv_8
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__152__B _153_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _206_/A mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_23 vpwr vgnd scs8hd_fill_2
XFILLER_19_56 vpwr vgnd scs8hd_fill_2
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
X_142_ _161_/A _140_/B _142_/Y vgnd vpwr scs8hd_nor2_4
X_211_ _211_/HI _211_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.tap_buf4_0_.scs8hd_inv_1 mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _223_/A vgnd vpwr scs8hd_inv_1
XANTENNA__147__B _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_132 vpwr vgnd scs8hd_fill_2
XFILLER_18_187 vpwr vgnd scs8hd_fill_2
XANTENNA__163__A _163_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_70 vpwr vgnd scs8hd_fill_2
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XFILLER_24_124 vpwr vgnd scs8hd_fill_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_79 vpwr vgnd scs8hd_fill_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_21_24 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _199_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__248__A _248_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_26 vpwr vgnd scs8hd_fill_2
X_125_ address[3] _134_/B _134_/C _126_/B vgnd vpwr scs8hd_or3_4
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XANTENNA__158__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_67 vgnd vpwr scs8hd_decap_3
XFILLER_32_56 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _106_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_105 vpwr vgnd scs8hd_fill_2
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.tap_buf4_0_.scs8hd_inv_1 mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _227_/A vgnd vpwr scs8hd_inv_1
X_108_ _107_/X _161_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_153 vpwr vgnd scs8hd_fill_2
XFILLER_11_193 vpwr vgnd scs8hd_fill_2
XFILLER_21_3 vgnd vpwr scs8hd_fill_1
XANTENNA__160__B _162_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_274 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _244_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_49 vpwr vgnd scs8hd_fill_2
XFILLER_16_241 vgnd vpwr scs8hd_decap_12
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__155__B _155_/B vgnd vpwr scs8hd_diode_2
XANTENNA__171__A _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_3_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_47 vgnd vpwr scs8hd_decap_4
XFILLER_38_99 vgnd vpwr scs8hd_decap_12
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
Xmux_left_track_15.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_204 vpwr vgnd scs8hd_fill_2
XFILLER_9_215 vpwr vgnd scs8hd_fill_2
XANTENNA__166__A _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_270 vgnd vpwr scs8hd_decap_4
XFILLER_39_196 vgnd vpwr scs8hd_decap_6
XFILLER_39_174 vpwr vgnd scs8hd_fill_2
XFILLER_24_13 vpwr vgnd scs8hd_fill_2
XFILLER_40_89 vgnd vpwr scs8hd_decap_3
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.LATCH_4_.latch data_in mem_bottom_track_1.LATCH_4_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XFILLER_10_59 vgnd vpwr scs8hd_decap_3
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_27_177 vgnd vpwr scs8hd_decap_6
X_210_ _210_/HI _210_/LO vgnd vpwr scs8hd_conb_1
X_141_ _131_/A _140_/B _141_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_111 vpwr vgnd scs8hd_fill_2
XANTENNA__147__C _184_/C vgnd vpwr scs8hd_diode_2
XFILLER_18_166 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _214_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _192_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_128 vpwr vgnd scs8hd_fill_2
XFILLER_15_136 vpwr vgnd scs8hd_fill_2
XFILLER_7_38 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_124_ address[4] _134_/B vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_7 vpwr vgnd scs8hd_fill_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_5_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__158__B _162_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__174__A _172_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_14 vgnd vpwr scs8hd_decap_3
XANTENNA__084__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_20_150 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A bottom_right_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_132 vpwr vgnd scs8hd_fill_2
XFILLER_7_176 vgnd vpwr scs8hd_decap_4
X_107_ address[1] address[2] _107_/C _107_/X vgnd vpwr scs8hd_or3_4
XANTENNA__169__A _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_81 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB _182_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A bottom_right_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_253 vpwr vgnd scs8hd_fill_2
XFILLER_16_253 vpwr vgnd scs8hd_fill_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XANTENNA__155__C _177_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_127 vpwr vgnd scs8hd_fill_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XFILLER_13_245 vpwr vgnd scs8hd_fill_2
XFILLER_0_171 vpwr vgnd scs8hd_fill_2
XFILLER_0_160 vpwr vgnd scs8hd_fill_2
XANTENNA__166__B _163_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A bottom_right_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__182__A _180_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_82 vpwr vgnd scs8hd_fill_2
XFILLER_5_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.INVTX1_2_.scs8hd_inv_1 left_bottom_grid_pin_12_ mux_left_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _201_/A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_8
XANTENNA__092__A _092_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_13.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XANTENNA__177__A _172_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
XFILLER_10_49 vgnd vpwr scs8hd_fill_1
XFILLER_27_101 vpwr vgnd scs8hd_fill_2
XFILLER_19_14 vpwr vgnd scs8hd_fill_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_35_68 vgnd vpwr scs8hd_fill_1
XFILLER_27_156 vpwr vgnd scs8hd_fill_2
XFILLER_27_123 vgnd vpwr scs8hd_fill_1
XANTENNA__087__A address[1] vgnd vpwr scs8hd_diode_2
X_140_ _140_/A _140_/B _140_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.INVTX1_2_.scs8hd_inv_1 bottom_right_grid_pin_3_ mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_211 vgnd vpwr scs8hd_decap_3
XFILLER_18_145 vgnd vpwr scs8hd_decap_8
XFILLER_33_137 vpwr vgnd scs8hd_fill_2
XFILLER_33_126 vgnd vpwr scs8hd_decap_8
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_15 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _214_/HI _205_/Y mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[2] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_123_ _133_/A _120_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_92 vgnd vpwr scs8hd_fill_1
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA__174__B _175_/B vgnd vpwr scs8hd_diode_2
XANTENNA__190__A _190_/A vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_3_.latch data_in mem_top_track_8.LATCH_3_.latch/Q _120_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _179_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_151 vpwr vgnd scs8hd_fill_2
XFILLER_11_173 vpwr vgnd scs8hd_fill_2
XFILLER_7_199 vpwr vgnd scs8hd_fill_2
X_106_ _099_/A _131_/A _106_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__169__B _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_240 vpwr vgnd scs8hd_fill_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _180_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_60 vpwr vgnd scs8hd_fill_2
XFILLER_27_69 vpwr vgnd scs8hd_fill_2
XFILLER_27_36 vgnd vpwr scs8hd_fill_1
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XFILLER_25_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__095__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_147 vgnd vpwr scs8hd_decap_4
XFILLER_4_18 vgnd vpwr scs8hd_decap_12
XFILLER_16_210 vgnd vpwr scs8hd_decap_4
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XFILLER_22_213 vgnd vpwr scs8hd_fill_1
XFILLER_13_16 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_1_117 vgnd vpwr scs8hd_decap_3
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
XFILLER_0_194 vgnd vpwr scs8hd_decap_12
XFILLER_0_150 vgnd vpwr scs8hd_decap_4
XANTENNA__166__C _166_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__182__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_39_143 vgnd vpwr scs8hd_decap_3
XFILLER_39_121 vgnd vpwr scs8hd_fill_1
XFILLER_39_154 vgnd vpwr scs8hd_decap_12
XFILLER_24_59 vpwr vgnd scs8hd_fill_2
XFILLER_6_6 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.LATCH_5_.latch data_in mem_bottom_track_9.LATCH_5_.latch/Q _149_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XFILLER_30_91 vgnd vpwr scs8hd_fill_1
XFILLER_36_113 vgnd vpwr scs8hd_decap_12
XFILLER_36_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB _176_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_track_7.LATCH_1_.latch data_in _195_/A _176_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__177__B _175_/B vgnd vpwr scs8hd_diode_2
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _200_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_48 vpwr vgnd scs8hd_fill_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_27_146 vpwr vgnd scs8hd_fill_2
XANTENNA__087__B _084_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_105 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_5_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 left_top_grid_pin_10_ mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_157 vpwr vgnd scs8hd_fill_2
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ _199_/A _199_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_2_84 vgnd vpwr scs8hd_decap_4
XANTENNA__188__A _172_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_4_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_49 vpwr vgnd scs8hd_fill_2
Xmux_left_track_11.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_8.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[5] mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__098__A _098_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_105 vgnd vpwr scs8hd_decap_4
XFILLER_15_116 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_71 vpwr vgnd scs8hd_fill_2
X_122_ _161_/A _120_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _204_/A mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_182 vpwr vgnd scs8hd_fill_2
XANTENNA__174__C _184_/C vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _128_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_263 vgnd vpwr scs8hd_decap_12
XFILLER_29_208 vgnd vpwr scs8hd_decap_12
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_16_49 vpwr vgnd scs8hd_fill_2
XFILLER_20_185 vgnd vpwr scs8hd_decap_3
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
XFILLER_7_101 vpwr vgnd scs8hd_fill_2
XFILLER_7_112 vpwr vgnd scs8hd_fill_2
X_105_ _105_/A _131_/A vgnd vpwr scs8hd_buf_1
XANTENNA__169__C _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_19_252 vgnd vpwr scs8hd_decap_12
XANTENNA__185__B _163_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__B _099_/A vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_70 vpwr vgnd scs8hd_fill_2
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _202_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_225 vgnd vpwr scs8hd_decap_12
XFILLER_22_203 vpwr vgnd scs8hd_fill_2
XFILLER_13_214 vgnd vpwr scs8hd_fill_1
XFILLER_13_225 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__166__D _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_251 vgnd vpwr scs8hd_decap_4
XANTENNA__182__C _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_39_166 vgnd vpwr scs8hd_decap_4
XFILLER_24_27 vpwr vgnd scs8hd_fill_2
XFILLER_10_206 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_125 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__177__C _177_/C vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_5_.latch data_in mem_bottom_track_17.LATCH_5_.latch/Q _157_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XANTENNA__087__C _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_33_117 vgnd vpwr scs8hd_decap_4
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _207_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ _198_/A _198_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__188__B _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_74 vgnd vpwr scs8hd_fill_1
XFILLER_2_30 vgnd vpwr scs8hd_fill_1
XFILLER_32_150 vgnd vpwr scs8hd_decap_3
XFILLER_24_128 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_180 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _189_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_150 vpwr vgnd scs8hd_fill_2
X_121_ _131_/A _120_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_50 vpwr vgnd scs8hd_fill_2
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__174__D _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_275 vpwr vgnd scs8hd_fill_2
XFILLER_37_253 vpwr vgnd scs8hd_fill_2
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_142 vgnd vpwr scs8hd_decap_8
Xmem_left_track_17.LATCH_0_.latch data_in _206_/A _188_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_93 vpwr vgnd scs8hd_fill_2
XFILLER_22_71 vgnd vpwr scs8hd_decap_4
XFILLER_22_60 vpwr vgnd scs8hd_fill_2
XFILLER_7_157 vpwr vgnd scs8hd_fill_2
X_104_ _104_/A address[2] _167_/A _105_/A vgnd vpwr scs8hd_or3_4
XFILLER_11_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__169__D _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_264 vgnd vpwr scs8hd_decap_12
XANTENNA__185__C _177_/C vgnd vpwr scs8hd_diode_2
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_49 vpwr vgnd scs8hd_fill_2
XFILLER_25_245 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_92 vpwr vgnd scs8hd_fill_2
XFILLER_3_193 vgnd vpwr scs8hd_decap_12
XFILLER_22_215 vgnd vpwr scs8hd_fill_1
XFILLER_22_237 vgnd vpwr scs8hd_decap_12
XFILLER_9_208 vgnd vpwr scs8hd_decap_4
XFILLER_9_219 vpwr vgnd scs8hd_fill_2
XFILLER_13_237 vgnd vpwr scs8hd_decap_6
XFILLER_0_185 vgnd vpwr scs8hd_fill_1
XFILLER_12_270 vgnd vpwr scs8hd_decap_4
XANTENNA__182__D _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_274 vgnd vpwr scs8hd_fill_1
XFILLER_39_178 vgnd vpwr scs8hd_decap_4
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _191_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_17 vpwr vgnd scs8hd_fill_2
XFILLER_10_218 vgnd vpwr scs8hd_decap_12
XFILLER_36_137 vgnd vpwr scs8hd_decap_12
XANTENNA__177__D _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XFILLER_2_203 vgnd vpwr scs8hd_decap_8
XFILLER_18_115 vgnd vpwr scs8hd_decap_4
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_25_60 vgnd vpwr scs8hd_fill_1
Xmux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _199_/A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
X_197_ _197_/A _197_/Y vgnd vpwr scs8hd_inv_8
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _240_/A vgnd vpwr scs8hd_inv_1
XFILLER_24_107 vpwr vgnd scs8hd_fill_2
XANTENNA__188__C _166_/C vgnd vpwr scs8hd_diode_2
XFILLER_2_53 vpwr vgnd scs8hd_fill_2
Xmem_left_track_3.LATCH_1_.latch data_in _191_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_173 vgnd vpwr scs8hd_decap_4
X_120_ _140_/A _120_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_95 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_154 vgnd vpwr scs8hd_decap_3
XFILLER_28_210 vgnd vpwr scs8hd_decap_4
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_11_132 vpwr vgnd scs8hd_fill_2
XFILLER_7_136 vpwr vgnd scs8hd_fill_2
X_103_ _099_/A _140_/A _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_19_276 vgnd vpwr scs8hd_fill_1
XFILLER_19_232 vgnd vpwr scs8hd_decap_8
Xmux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _213_/HI _203_/Y mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__185__D _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_39 vgnd vpwr scs8hd_fill_1
XFILLER_27_17 vgnd vpwr scs8hd_decap_4
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_202 vpwr vgnd scs8hd_fill_2
XFILLER_16_224 vgnd vpwr scs8hd_decap_3
XFILLER_17_83 vpwr vgnd scs8hd_fill_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_71 vgnd vpwr scs8hd_fill_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_161 vgnd vpwr scs8hd_decap_3
XFILLER_22_249 vgnd vpwr scs8hd_decap_12
XFILLER_1_109 vpwr vgnd scs8hd_fill_2
XFILLER_13_249 vgnd vpwr scs8hd_decap_6
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _210_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_175 vpwr vgnd scs8hd_fill_2
XFILLER_0_164 vgnd vpwr scs8hd_decap_4
XFILLER_5_86 vgnd vpwr scs8hd_decap_4
XFILLER_5_75 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_39_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
XFILLER_5_201 vpwr vgnd scs8hd_fill_2
XFILLER_5_212 vgnd vpwr scs8hd_decap_12
XFILLER_14_73 vpwr vgnd scs8hd_fill_2
XFILLER_14_84 vpwr vgnd scs8hd_fill_2
XFILLER_30_83 vgnd vpwr scs8hd_decap_8
XFILLER_30_72 vpwr vgnd scs8hd_fill_2
XFILLER_30_50 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XFILLER_39_81 vpwr vgnd scs8hd_fill_2
XFILLER_36_149 vgnd vpwr scs8hd_decap_4
XANTENNA__101__A _104_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_19_18 vgnd vpwr scs8hd_decap_3
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_127 vpwr vgnd scs8hd_fill_2
XFILLER_4_6 vgnd vpwr scs8hd_decap_12
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_26_171 vpwr vgnd scs8hd_fill_2
XFILLER_25_94 vpwr vgnd scs8hd_fill_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
X_196_ _196_/A _196_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_3_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_3
XANTENNA__188__D _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_19 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _207_/HI mem_bottom_track_1.LATCH_2_.latch/Q
+ mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_163 vgnd vpwr scs8hd_decap_3
X_248_ _248_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
X_179_ _172_/X _175_/B _166_/C _167_/X _179_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_16_19 vpwr vgnd scs8hd_fill_2
XFILLER_20_166 vpwr vgnd scs8hd_fill_2
XFILLER_11_155 vpwr vgnd scs8hd_fill_2
XFILLER_22_84 vgnd vpwr scs8hd_decap_8
XFILLER_22_51 vgnd vpwr scs8hd_decap_3
XFILLER_22_40 vpwr vgnd scs8hd_fill_2
X_102_ _102_/A _140_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_177 vgnd vpwr scs8hd_decap_4
XFILLER_19_211 vpwr vgnd scs8hd_fill_2
XFILLER_8_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_203 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _202_/A mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_4_118 vgnd vpwr scs8hd_fill_1
XFILLER_17_62 vgnd vpwr scs8hd_fill_1
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_151 vgnd vpwr scs8hd_decap_4
XANTENNA__104__A _104_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _199_/Y vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_13.LATCH_0_.latch data_in _202_/A _184_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_217 vgnd vpwr scs8hd_fill_1
XFILLER_28_50 vgnd vpwr scs8hd_decap_8
XFILLER_0_154 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_10 vpwr vgnd scs8hd_fill_2
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _103_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_bottom_track_9.LATCH_0_.latch data_in mem_bottom_track_9.LATCH_0_.latch/Q _154_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _206_/Y mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_11.tap_buf4_0_.scs8hd_inv_1 mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _225_/A vgnd vpwr scs8hd_inv_1
XFILLER_30_40 vgnd vpwr scs8hd_fill_1
XFILLER_5_224 vgnd vpwr scs8hd_decap_12
XFILLER_14_52 vgnd vpwr scs8hd_decap_4
XFILLER_14_96 vgnd vpwr scs8hd_decap_8
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XFILLER_39_93 vpwr vgnd scs8hd_fill_2
XFILLER_36_106 vgnd vpwr scs8hd_decap_4
XANTENNA__101__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 bottom_right_grid_pin_1_ mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 top_right_grid_pin_7_ mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_109 vgnd vpwr scs8hd_decap_6
XFILLER_18_128 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vpwr vgnd scs8hd_fill_2
XFILLER_25_51 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ _195_/A _195_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_66 vpwr vgnd scs8hd_fill_2
XANTENNA__112__A _099_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vgnd vpwr scs8hd_fill_1
XFILLER_17_172 vpwr vgnd scs8hd_fill_2
XFILLER_32_142 vgnd vpwr scs8hd_decap_8
Xmux_left_track_3.tap_buf4_0_.scs8hd_inv_1 mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _229_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_197 vgnd vpwr scs8hd_decap_8
XFILLER_11_75 vpwr vgnd scs8hd_fill_2
X_247_ chany_bottom_in[0] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__107__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_14_186 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _201_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_178_ _172_/X _175_/B _166_/C _165_/X _178_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_37_245 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_1.LATCH_5_.latch data_in mem_bottom_track_1.LATCH_5_.latch/Q _138_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_101_ _104_/A address[2] _165_/A _102_/A vgnd vpwr scs8hd_or3_4
XFILLER_7_105 vpwr vgnd scs8hd_fill_2
XFILLER_7_116 vgnd vpwr scs8hd_decap_4
XFILLER_11_101 vpwr vgnd scs8hd_fill_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vpwr vgnd scs8hd_fill_2
XFILLER_8_43 vpwr vgnd scs8hd_fill_2
XFILLER_8_87 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_7_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_259 vgnd vpwr scs8hd_decap_12
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_84 vpwr vgnd scs8hd_fill_2
XFILLER_33_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _192_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__104__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _140_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
XFILLER_22_207 vgnd vpwr scs8hd_decap_6
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _197_/A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_38_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_262 vgnd vpwr scs8hd_decap_12
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
XANTENNA__115__A _114_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_17.LATCH_0_.latch data_in mem_bottom_track_17.LATCH_0_.latch/Q _162_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_8.LATCH_4_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_5_236 vgnd vpwr scs8hd_decap_8
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_39_50 vgnd vpwr scs8hd_decap_8
XFILLER_30_96 vpwr vgnd scs8hd_fill_2
XANTENNA__101__C _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[4] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _194_/A _194_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__112__B _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_32_121 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_140 vpwr vgnd scs8hd_fill_2
XFILLER_17_195 vpwr vgnd scs8hd_fill_2
XFILLER_23_154 vpwr vgnd scs8hd_fill_2
XFILLER_23_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A bottom_right_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_54 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _194_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_121 vpwr vgnd scs8hd_fill_2
X_246_ chany_bottom_in[1] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__107__B address[2] vgnd vpwr scs8hd_diode_2
X_177_ _172_/X _175_/B _177_/C _167_/X _177_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__123__A _133_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_124 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
X_100_ address[1] _104_/A vgnd vpwr scs8hd_inv_8
XFILLER_11_168 vgnd vpwr scs8hd_decap_3
XFILLER_34_238 vgnd vpwr scs8hd_decap_12
XFILLER_34_227 vgnd vpwr scs8hd_decap_8
XANTENNA__118__A _128_/A vgnd vpwr scs8hd_diode_2
X_229_ _229_/A chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_6_150 vgnd vpwr scs8hd_decap_3
XFILLER_8_77 vpwr vgnd scs8hd_fill_2
XFILLER_25_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_33_74 vgnd vpwr scs8hd_fill_1
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XANTENNA__104__C _167_/A vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _120_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _212_/HI _201_/Y mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _192_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_274 vgnd vpwr scs8hd_decap_3
XFILLER_0_134 vgnd vpwr scs8hd_decap_8
Xmux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_74 vgnd vpwr scs8hd_decap_12
XFILLER_12_274 vgnd vpwr scs8hd_fill_1
Xmem_top_track_8.LATCH_4_.latch data_in mem_top_track_8.LATCH_4_.latch/Q _119_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_34 vpwr vgnd scs8hd_fill_2
XFILLER_5_23 vpwr vgnd scs8hd_fill_2
XANTENNA__131__A _131_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_5_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_29_182 vgnd vpwr scs8hd_fill_1
XANTENNA__126__A _136_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_25_20 vpwr vgnd scs8hd_fill_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_25_75 vpwr vgnd scs8hd_fill_2
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_193_ _193_/A _193_/Y vgnd vpwr scs8hd_inv_8
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_17_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_6 vgnd vpwr scs8hd_decap_12
XFILLER_11_33 vpwr vgnd scs8hd_fill_2
XFILLER_11_88 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_3_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_245_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__107__C _107_/C vgnd vpwr scs8hd_diode_2
X_176_ _172_/X _175_/B _177_/C _165_/X _176_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__123__B _120_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vpwr vgnd scs8hd_fill_2
XFILLER_22_10 vpwr vgnd scs8hd_fill_2
XFILLER_11_136 vpwr vgnd scs8hd_fill_2
XANTENNA__224__A _224_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_12 vgnd vpwr scs8hd_decap_4
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XANTENNA__118__B _120_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_184 vpwr vgnd scs8hd_fill_2
X_159_ _140_/A _162_/B _159_/Y vgnd vpwr scs8hd_nor2_4
X_228_ _228_/A chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__134__A _134_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_3 vpwr vgnd scs8hd_fill_2
XFILLER_25_239 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_206 vpwr vgnd scs8hd_fill_2
XFILLER_17_32 vpwr vgnd scs8hd_fill_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_53 vpwr vgnd scs8hd_fill_2
XFILLER_33_42 vpwr vgnd scs8hd_fill_2
XFILLER_33_31 vgnd vpwr scs8hd_decap_8
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_87 vpwr vgnd scs8hd_fill_2
XANTENNA__129__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_179 vgnd vpwr scs8hd_decap_6
XFILLER_0_146 vpwr vgnd scs8hd_fill_2
Xmux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _200_/A mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_28_86 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _215_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB _186_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XANTENNA__131__B _132_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XFILLER_14_88 vpwr vgnd scs8hd_fill_2
XANTENNA__232__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_30_76 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_8
XFILLER_39_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__126__B _126_/B vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_5_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_175 vgnd vpwr scs8hd_decap_4
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_32 vpwr vgnd scs8hd_fill_2
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XANTENNA__227__A _227_/A vgnd vpwr scs8hd_diode_2
XPHY_32 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _202_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/A _192_/Y vgnd vpwr scs8hd_inv_8
XFILLER_25_98 vgnd vpwr scs8hd_decap_4
Xmux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _204_/Y mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XANTENNA__137__A _136_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_112 vgnd vpwr scs8hd_decap_3
XFILLER_11_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_244_ _244_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_14_134 vgnd vpwr scs8hd_decap_6
XFILLER_14_145 vgnd vpwr scs8hd_decap_8
X_175_ _172_/X _175_/B _184_/C _167_/X _175_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_37_259 vpwr vgnd scs8hd_fill_2
XFILLER_9_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB _183_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XANTENNA__240__A _240_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_248 vpwr vgnd scs8hd_fill_2
XFILLER_19_215 vpwr vgnd scs8hd_fill_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
X_227_ _227_/A chanx_left_out[3] vgnd vpwr scs8hd_buf_2
X_158_ _119_/A _162_/B _158_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_130 vgnd vpwr scs8hd_decap_8
XFILLER_6_141 vgnd vpwr scs8hd_decap_3
XANTENNA__134__B _134_/B vgnd vpwr scs8hd_diode_2
X_089_ address[6] address[5] _136_/A vgnd vpwr scs8hd_or2_4
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__150__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_229 vgnd vpwr scs8hd_decap_3
XFILLER_17_66 vpwr vgnd scs8hd_fill_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_251 vgnd vpwr scs8hd_decap_12
XANTENNA__235__A _235_/A vgnd vpwr scs8hd_diode_2
XANTENNA__129__B _132_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _204_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_103 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_3
XFILLER_0_114 vpwr vgnd scs8hd_fill_2
XFILLER_8_258 vgnd vpwr scs8hd_decap_12
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_14 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_6 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_1_.latch data_in _205_/A _187_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _195_/A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_12 vpwr vgnd scs8hd_fill_2
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_14_56 vgnd vpwr scs8hd_fill_1
XFILLER_39_97 vgnd vpwr scs8hd_decap_12
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XFILLER_29_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__142__B _140_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_110 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _219_/HI mem_top_track_0.LATCH_2_.latch/Q
+ mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vgnd vpwr scs8hd_decap_6
XFILLER_26_132 vpwr vgnd scs8hd_fill_2
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
X_191_ _191_/A _191_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__243__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_17_165 vgnd vpwr scs8hd_decap_4
XFILLER_17_176 vgnd vpwr scs8hd_decap_4
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_46 vpwr vgnd scs8hd_fill_2
XFILLER_36_76 vgnd vpwr scs8hd_fill_1
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XANTENNA__238__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_0_.latch data_in mem_bottom_track_1.LATCH_0_.latch/Q _143_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _191_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_190 vgnd vpwr scs8hd_decap_4
X_243_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_14_168 vgnd vpwr scs8hd_decap_3
X_174_ _172_/X _175_/B _184_/C _165_/X _174_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_28_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ _192_/A mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__148__A _147_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_105 vpwr vgnd scs8hd_fill_2
XFILLER_20_116 vgnd vpwr scs8hd_decap_8
XFILLER_20_138 vpwr vgnd scs8hd_fill_2
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XFILLER_22_23 vpwr vgnd scs8hd_fill_2
XFILLER_22_67 vpwr vgnd scs8hd_fill_2
XFILLER_22_56 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_4_.scs8hd_inv_1 bottom_right_grid_pin_15_ mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[4] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_226_ _226_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_8_36 vgnd vpwr scs8hd_decap_4
XFILLER_8_47 vgnd vpwr scs8hd_decap_4
X_157_ _128_/A _162_/B _157_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__C _134_/C vgnd vpwr scs8hd_diode_2
XFILLER_40_6 vgnd vpwr scs8hd_decap_12
XANTENNA__150__B _153_/B vgnd vpwr scs8hd_diode_2
X_088_ _088_/A _128_/A vgnd vpwr scs8hd_buf_1
XFILLER_19_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_263 vgnd vpwr scs8hd_decap_12
XFILLER_17_12 vpwr vgnd scs8hd_fill_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_88 vpwr vgnd scs8hd_fill_2
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.INVTX1_5_.scs8hd_inv_1 chanx_left_in[1] mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_134 vpwr vgnd scs8hd_fill_2
XFILLER_30_211 vgnd vpwr scs8hd_decap_3
XFILLER_15_252 vgnd vpwr scs8hd_decap_3
X_209_ _209_/HI _209_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_22 vgnd vpwr scs8hd_decap_3
XFILLER_28_11 vpwr vgnd scs8hd_fill_2
XANTENNA__246__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_12_211 vgnd vpwr scs8hd_decap_3
XFILLER_12_222 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__156__A _155_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_35 vpwr vgnd scs8hd_fill_2
XFILLER_30_23 vgnd vpwr scs8hd_decap_8
XFILLER_39_65 vpwr vgnd scs8hd_fill_2
XFILLER_39_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _193_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
XFILLER_29_174 vgnd vpwr scs8hd_decap_8
Xmux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _211_/HI _199_/Y mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 top_right_grid_pin_5_ mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_12 vpwr vgnd scs8hd_fill_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
X_190_ _190_/A _190_/Y vgnd vpwr scs8hd_inv_8
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_188 vgnd vpwr scs8hd_decap_12
XFILLER_25_56 vpwr vgnd scs8hd_fill_2
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_2_49 vpwr vgnd scs8hd_fill_2
XFILLER_2_38 vgnd vpwr scs8hd_decap_6
XFILLER_17_100 vpwr vgnd scs8hd_fill_2
XFILLER_17_144 vgnd vpwr scs8hd_fill_1
XFILLER_17_199 vpwr vgnd scs8hd_fill_2
XANTENNA__153__B _153_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_169 vpwr vgnd scs8hd_fill_2
XFILLER_23_136 vgnd vpwr scs8hd_decap_3
XFILLER_11_58 vgnd vpwr scs8hd_fill_1
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
X_242_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
X_173_ address[5] _175_/B vgnd vpwr scs8hd_buf_1
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _198_/A mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__164__A _126_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_162 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _216_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_81 vpwr vgnd scs8hd_fill_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_228 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_1.INVTX1_7_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_156_ _155_/X _162_/B vgnd vpwr scs8hd_buf_1
XFILLER_6_110 vgnd vpwr scs8hd_decap_3
XFILLER_6_154 vpwr vgnd scs8hd_fill_2
XFILLER_6_165 vpwr vgnd scs8hd_fill_2
X_087_ address[1] _084_/Y _165_/A _088_/A vgnd vpwr scs8hd_or3_4
XFILLER_10_161 vpwr vgnd scs8hd_fill_2
X_225_ _225_/A chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XANTENNA__159__A _140_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[5] mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XFILLER_33_67 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_220 vpwr vgnd scs8hd_fill_2
XFILLER_15_231 vpwr vgnd scs8hd_fill_2
X_208_ _208_/HI _208_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__161__B _162_/B vgnd vpwr scs8hd_diode_2
X_139_ _119_/A _140_/B _139_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_track_7.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[8] mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_201 vpwr vgnd scs8hd_fill_2
XFILLER_21_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_205 vgnd vpwr scs8hd_decap_8
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XFILLER_12_234 vgnd vpwr scs8hd_decap_12
XFILLER_5_38 vpwr vgnd scs8hd_fill_2
XFILLER_5_27 vpwr vgnd scs8hd_fill_2
XFILLER_39_109 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _172_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A left_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_69 vpwr vgnd scs8hd_fill_2
XFILLER_5_208 vpwr vgnd scs8hd_fill_2
XFILLER_39_77 vgnd vpwr scs8hd_fill_1
XFILLER_29_153 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XANTENNA__167__A _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_70 vgnd vpwr scs8hd_decap_3
XFILLER_26_145 vpwr vgnd scs8hd_fill_2
XFILLER_25_24 vgnd vpwr scs8hd_fill_1
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
Xmem_left_track_13.LATCH_1_.latch data_in _201_/A _183_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_32_104 vgnd vpwr scs8hd_decap_8
XFILLER_17_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_181 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _099_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_bottom_track_9.LATCH_1_.latch data_in mem_bottom_track_9.LATCH_1_.latch/Q _153_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_104 vpwr vgnd scs8hd_fill_2
X_172_ _172_/A _172_/X vgnd vpwr scs8hd_buf_1
X_241_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_170 vpwr vgnd scs8hd_fill_2
XANTENNA__180__A _172_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_71 vgnd vpwr scs8hd_decap_4
Xmux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _202_/Y mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XFILLER_22_36 vpwr vgnd scs8hd_fill_2
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A enable vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_0_.latch data_in _198_/A _179_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_16 vgnd vpwr scs8hd_fill_1
XFILLER_8_27 vpwr vgnd scs8hd_fill_2
X_224_ _224_/A chanx_left_out[6] vgnd vpwr scs8hd_buf_2
X_086_ _107_/C _165_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_188 vpwr vgnd scs8hd_fill_2
XFILLER_10_195 vgnd vpwr scs8hd_decap_6
X_155_ address[6] _155_/B _177_/C _155_/X vgnd vpwr scs8hd_or3_4
XFILLER_33_7 vgnd vpwr scs8hd_decap_12
XFILLER_26_6 vpwr vgnd scs8hd_fill_2
XFILLER_33_243 vgnd vpwr scs8hd_fill_1
XFILLER_33_232 vgnd vpwr scs8hd_decap_3
XANTENNA__159__B _162_/B vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _172_/X vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_57 vpwr vgnd scs8hd_fill_2
XFILLER_33_46 vgnd vpwr scs8hd_decap_4
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XANTENNA__085__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_103 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_243 vgnd vpwr scs8hd_fill_1
X_207_ _207_/HI _207_/LO vgnd vpwr scs8hd_conb_1
X_138_ _128_/A _140_/B _138_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_191 vgnd vpwr scs8hd_decap_12
XFILLER_2_180 vpwr vgnd scs8hd_fill_2
XFILLER_21_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _201_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XFILLER_12_246 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
XFILLER_14_59 vgnd vpwr scs8hd_fill_1
XFILLER_30_58 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_5.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[7] mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_2_.scs8hd_inv_1 bottom_right_grid_pin_5_ mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
XANTENNA__183__A _180_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _248_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_25_47 vpwr vgnd scs8hd_fill_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XANTENNA__093__A _136_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_12
XFILLER_2_18 vgnd vpwr scs8hd_decap_12
XFILLER_32_138 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _193_/A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_31_90 vpwr vgnd scs8hd_fill_2
XANTENNA__178__A _172_/X vgnd vpwr scs8hd_diode_2
XFILLER_11_16 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A _088_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_8
X_240_ _240_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_171_ _169_/A _172_/A vgnd vpwr scs8hd_inv_8
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_17.LATCH_1_.latch data_in mem_bottom_track_17.LATCH_1_.latch/Q _161_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_153 vgnd vpwr scs8hd_fill_1
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_193 vpwr vgnd scs8hd_fill_2
XFILLER_9_197 vpwr vgnd scs8hd_fill_2
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _203_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_27_263 vgnd vpwr scs8hd_decap_12
X_223_ _223_/A chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_10_152 vgnd vpwr scs8hd_fill_1
X_154_ _133_/A _153_/B _154_/Y vgnd vpwr scs8hd_nor2_4
X_085_ address[0] _107_/C vgnd vpwr scs8hd_inv_8
Xmux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _218_/HI _197_/Y mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__175__B _175_/B vgnd vpwr scs8hd_diode_2
XANTENNA__191__A _191_/A vgnd vpwr scs8hd_diode_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ _190_/A mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_206_ _206_/A _206_/Y vgnd vpwr scs8hd_inv_8
X_137_ _136_/X _140_/B vgnd vpwr scs8hd_buf_1
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_258 vpwr vgnd scs8hd_fill_2
XFILLER_0_84 vpwr vgnd scs8hd_fill_2
XANTENNA__186__A _180_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _222_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _194_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_107 vgnd vpwr scs8hd_decap_4
XFILLER_0_118 vgnd vpwr scs8hd_decap_4
XFILLER_28_58 vgnd vpwr scs8hd_decap_3
XANTENNA__096__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_12_203 vgnd vpwr scs8hd_decap_8
Xmux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_top_track_8.LATCH_5_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_12_258 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A top_right_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_111 vgnd vpwr scs8hd_decap_12
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_16 vpwr vgnd scs8hd_fill_2
XFILLER_14_27 vpwr vgnd scs8hd_fill_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
XFILLER_35_114 vgnd vpwr scs8hd_decap_8
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _226_/A vgnd vpwr scs8hd_inv_1
XANTENNA__183__B _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_61 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A bottom_right_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__B _184_/C vgnd vpwr scs8hd_diode_2
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XFILLER_1_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_136 vpwr vgnd scs8hd_fill_2
XFILLER_17_169 vgnd vpwr scs8hd_fill_1
XFILLER_25_191 vgnd vpwr scs8hd_decap_12
Xmux_left_track_3.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[3] mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _192_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__194__A _194_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_117 vgnd vpwr scs8hd_decap_3
XANTENNA__178__B _175_/B vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_5_.latch data_in mem_top_track_8.LATCH_5_.latch/Q _118_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_161 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
X_170_ _169_/A _163_/X _169_/C _167_/X _170_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_22_150 vgnd vpwr scs8hd_decap_3
XFILLER_14_117 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_132 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _196_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_27 vpwr vgnd scs8hd_fill_2
XANTENNA__099__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_275 vpwr vgnd scs8hd_fill_2
XFILLER_27_253 vpwr vgnd scs8hd_fill_2
XFILLER_27_220 vgnd vpwr scs8hd_decap_12
X_222_ _222_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_6_102 vgnd vpwr scs8hd_decap_8
XFILLER_10_131 vgnd vpwr scs8hd_decap_4
X_153_ _161_/A _153_/B _153_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_146 vpwr vgnd scs8hd_fill_2
XFILLER_12_60 vpwr vgnd scs8hd_fill_2
X_084_ address[2] _084_/Y vgnd vpwr scs8hd_inv_8
XFILLER_12_82 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_15_ mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
XANTENNA__175__C _184_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _196_/A mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_212 vpwr vgnd scs8hd_fill_2
XFILLER_17_16 vgnd vpwr scs8hd_decap_3
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_205_ _205_/A _205_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_136_ _136_/A _169_/C _136_/X vgnd vpwr scs8hd_or2_4
Xmem_left_track_5.LATCH_0_.latch data_in _194_/A _175_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_63 vgnd vpwr scs8hd_decap_4
XANTENNA__186__B _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_226 vgnd vpwr scs8hd_decap_12
XFILLER_9_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _219_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_91 vgnd vpwr scs8hd_fill_1
X_119_ _119_/A _120_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_123 vgnd vpwr scs8hd_decap_12
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_39 vpwr vgnd scs8hd_fill_2
XFILLER_39_14 vgnd vpwr scs8hd_decap_12
XFILLER_39_69 vgnd vpwr scs8hd_decap_8
XFILLER_39_58 vgnd vpwr scs8hd_decap_3
XFILLER_29_123 vpwr vgnd scs8hd_fill_2
XFILLER_29_112 vpwr vgnd scs8hd_fill_2
XFILLER_29_101 vpwr vgnd scs8hd_fill_2
XFILLER_20_71 vpwr vgnd scs8hd_fill_2
XFILLER_20_93 vgnd vpwr scs8hd_decap_3
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XANTENNA__183__C _184_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XFILLER_26_104 vpwr vgnd scs8hd_fill_2
XFILLER_25_16 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_269 vgnd vpwr scs8hd_decap_8
XFILLER_1_214 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_4_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_104 vpwr vgnd scs8hd_fill_2
XFILLER_17_148 vpwr vgnd scs8hd_fill_2
XFILLER_25_181 vpwr vgnd scs8hd_fill_2
XFILLER_15_82 vpwr vgnd scs8hd_fill_2
XANTENNA__178__C _166_/C vgnd vpwr scs8hd_diode_2
XFILLER_16_181 vgnd vpwr scs8hd_decap_3
XFILLER_16_192 vgnd vpwr scs8hd_fill_1
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_31_173 vgnd vpwr scs8hd_decap_8
XFILLER_11_29 vpwr vgnd scs8hd_fill_2
XFILLER_39_262 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_173 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.INVTX1_4_.scs8hd_inv_1 bottom_right_grid_pin_13_ mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _217_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__B _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_232 vgnd vpwr scs8hd_decap_12
X_152_ _131_/A _153_/B _152_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_19 vgnd vpwr scs8hd_fill_1
XFILLER_10_165 vpwr vgnd scs8hd_fill_2
XFILLER_12_72 vgnd vpwr scs8hd_fill_1
X_221_ _221_/HI _221_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_8.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[1] mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_169 vgnd vpwr scs8hd_decap_4
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XANTENNA__175__D _167_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_28 vpwr vgnd scs8hd_fill_2
Xmux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _200_/Y mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
X_204_ _204_/A _204_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_224 vpwr vgnd scs8hd_fill_2
XFILLER_15_235 vgnd vpwr scs8hd_decap_8
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
XFILLER_23_93 vpwr vgnd scs8hd_fill_2
X_135_ _134_/X _169_/C vgnd vpwr scs8hd_buf_1
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_7 vpwr vgnd scs8hd_fill_2
XANTENNA__186__C _177_/C vgnd vpwr scs8hd_diode_2
XFILLER_21_238 vgnd vpwr scs8hd_decap_6
XFILLER_9_62 vgnd vpwr scs8hd_decap_4
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_93 vpwr vgnd scs8hd_fill_2
XFILLER_34_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB _174_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_242 vpwr vgnd scs8hd_fill_2
XFILLER_7_253 vpwr vgnd scs8hd_fill_2
X_118_ _128_/A _120_/B _118_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_135 vgnd vpwr scs8hd_decap_12
XFILLER_39_26 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_41 vgnd vpwr scs8hd_fill_1
XANTENNA__183__D _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_149 vgnd vpwr scs8hd_decap_4
XFILLER_26_116 vgnd vpwr scs8hd_decap_3
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_28 vpwr vgnd scs8hd_fill_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_226 vgnd vpwr scs8hd_decap_12
XFILLER_25_160 vpwr vgnd scs8hd_fill_2
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XFILLER_31_60 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _204_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__178__D _165_/X vgnd vpwr scs8hd_diode_2
XFILLER_31_130 vpwr vgnd scs8hd_fill_2
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
XFILLER_39_241 vgnd vpwr scs8hd_decap_3
XFILLER_39_274 vgnd vpwr scs8hd_decap_3
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_71 vpwr vgnd scs8hd_fill_2
XFILLER_13_174 vpwr vgnd scs8hd_fill_2
XFILLER_9_156 vgnd vpwr scs8hd_decap_4
XFILLER_3_53 vgnd vpwr scs8hd_decap_4
XFILLER_3_42 vpwr vgnd scs8hd_fill_2
XFILLER_3_31 vgnd vpwr scs8hd_decap_8
Xmux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _191_/A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_220_ _220_/HI _220_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
X_151_ _140_/A _153_/B _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_115 vgnd vpwr scs8hd_decap_4
XFILLER_10_111 vgnd vpwr scs8hd_decap_3
XFILLER_10_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _220_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[3] mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_92 vpwr vgnd scs8hd_fill_2
XFILLER_18_222 vgnd vpwr scs8hd_fill_1
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_107 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_203 vpwr vgnd scs8hd_fill_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_203_ _203_/A _203_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
XFILLER_23_83 vgnd vpwr scs8hd_decap_4
X_134_ _134_/A _134_/B _134_/C _134_/X vgnd vpwr scs8hd_or3_4
Xmem_bottom_track_1.LATCH_1_.latch data_in mem_bottom_track_1.LATCH_1_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_184 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_4
XFILLER_0_43 vgnd vpwr scs8hd_decap_6
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XANTENNA__186__D _167_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _217_/HI _195_/Y mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_34_93 vgnd vpwr scs8hd_decap_3
XFILLER_34_60 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _206_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_210 vgnd vpwr scs8hd_decap_12
X_117_ _116_/X _120_/B vgnd vpwr scs8hd_buf_1
XFILLER_38_147 vgnd vpwr scs8hd_decap_6
Xmem_left_track_1.LATCH_0_.latch data_in _190_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_18 vpwr vgnd scs8hd_fill_2
XFILLER_39_38 vgnd vpwr scs8hd_decap_12
XFILLER_29_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_84 vgnd vpwr scs8hd_decap_3
XFILLER_6_64 vgnd vpwr scs8hd_decap_4
XFILLER_26_128 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_1_238 vgnd vpwr scs8hd_decap_6
XFILLER_15_62 vgnd vpwr scs8hd_decap_3
XFILLER_31_94 vgnd vpwr scs8hd_decap_3
XFILLER_31_83 vpwr vgnd scs8hd_fill_2
XANTENNA__102__A _102_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _215_/HI _192_/Y mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_253 vpwr vgnd scs8hd_fill_2
XFILLER_22_142 vgnd vpwr scs8hd_decap_8
XFILLER_22_186 vpwr vgnd scs8hd_fill_2
XFILLER_9_102 vgnd vpwr scs8hd_decap_3
XFILLER_13_153 vpwr vgnd scs8hd_fill_2
XFILLER_13_197 vpwr vgnd scs8hd_fill_2
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_98 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _193_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_8
X_150_ _119_/A _153_/B _150_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_178 vgnd vpwr scs8hd_decap_6
XFILLER_12_96 vpwr vgnd scs8hd_fill_2
XFILLER_37_82 vpwr vgnd scs8hd_fill_2
XFILLER_33_237 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A top_right_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XFILLER_24_204 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _187_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_248 vpwr vgnd scs8hd_fill_2
X_133_ _133_/A _132_/B _133_/Y vgnd vpwr scs8hd_nor2_4
X_202_ _202_/A _202_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_163 vgnd vpwr scs8hd_decap_3
XANTENNA__110__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_0_88 vgnd vpwr scs8hd_decap_3
XFILLER_9_53 vgnd vpwr scs8hd_decap_6
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_218 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _194_/A mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_18_84 vpwr vgnd scs8hd_fill_2
XFILLER_7_222 vgnd vpwr scs8hd_decap_12
XANTENNA__105__A _105_/A vgnd vpwr scs8hd_diode_2
X_116_ _136_/A _177_/C _116_/X vgnd vpwr scs8hd_or2_4
XFILLER_20_30 vgnd vpwr scs8hd_fill_1
XFILLER_20_41 vpwr vgnd scs8hd_fill_2
XFILLER_6_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _195_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_0_.latch data_in mem_top_track_8.LATCH_0_.latch/Q _123_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_173 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vgnd vpwr scs8hd_decap_6
XFILLER_31_51 vpwr vgnd scs8hd_fill_2
XFILLER_31_40 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _198_/Y mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_261 vgnd vpwr scs8hd_decap_12
XFILLER_16_162 vgnd vpwr scs8hd_decap_8
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_210 vgnd vpwr scs8hd_decap_8
XFILLER_22_154 vpwr vgnd scs8hd_fill_2
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_84 vgnd vpwr scs8hd_decap_8
XFILLER_26_51 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_77 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_10_102 vgnd vpwr scs8hd_decap_3
XFILLER_10_157 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_42 vpwr vgnd scs8hd_fill_2
XFILLER_12_64 vpwr vgnd scs8hd_fill_2
XFILLER_12_86 vgnd vpwr scs8hd_fill_1
XFILLER_18_235 vgnd vpwr scs8hd_decap_8
XFILLER_18_246 vgnd vpwr scs8hd_decap_8
XFILLER_18_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__108__A _107_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_172 vpwr vgnd scs8hd_fill_2
XFILLER_24_227 vgnd vpwr scs8hd_decap_12
XFILLER_33_19 vgnd vpwr scs8hd_decap_12
X_132_ _161_/A _132_/B _132_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _095_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_201_ _201_/A _201_/Y vgnd vpwr scs8hd_inv_8
Xmem_bottom_track_9.LATCH_2_.latch data_in mem_bottom_track_9.LATCH_2_.latch/Q _152_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_21_208 vgnd vpwr scs8hd_decap_3
XFILLER_14_271 vgnd vpwr scs8hd_decap_4
XFILLER_9_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_63 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_7_234 vgnd vpwr scs8hd_decap_8
XFILLER_7_245 vgnd vpwr scs8hd_decap_8
XFILLER_11_263 vgnd vpwr scs8hd_decap_12
X_115_ _114_/X _177_/C vgnd vpwr scs8hd_buf_1
XFILLER_22_6 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_1_.latch data_in _197_/A _178_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__121__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_116 vgnd vpwr scs8hd_decap_4
XFILLER_29_105 vpwr vgnd scs8hd_fill_2
XFILLER_37_171 vgnd vpwr scs8hd_decap_12
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XFILLER_29_51 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_20_75 vpwr vgnd scs8hd_fill_2
XFILLER_29_84 vpwr vgnd scs8hd_fill_2
XANTENNA__116__A _136_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_55 vgnd vpwr scs8hd_decap_6
XFILLER_6_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_108 vgnd vpwr scs8hd_decap_8
XFILLER_20_3 vpwr vgnd scs8hd_fill_2
XFILLER_34_152 vgnd vpwr scs8hd_fill_1
XFILLER_25_130 vpwr vgnd scs8hd_fill_2
XFILLER_17_108 vgnd vpwr scs8hd_decap_3
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_86 vpwr vgnd scs8hd_fill_2
XFILLER_0_273 vgnd vpwr scs8hd_decap_4
XFILLER_16_130 vpwr vgnd scs8hd_fill_2
XFILLER_16_141 vpwr vgnd scs8hd_fill_2
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _209_/HI vgnd vpwr
+ scs8hd_diode_2
.ends

