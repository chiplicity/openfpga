magic
tech sky130A
magscale 1 2
timestamp 1604669046
<< locali >>
rect 10609 11679 10643 11849
rect 9505 11543 9539 11645
rect 10609 11543 10643 11645
rect 11989 10523 12023 10625
rect 2421 9503 2455 9605
rect 2513 9367 2547 9469
rect 4077 6171 4111 6409
rect 10333 6239 10367 6341
rect 15945 3927 15979 4029
rect 6745 2295 6779 2601
<< viali >>
rect 24777 23273 24811 23307
rect 24593 23137 24627 23171
rect 1593 22729 1627 22763
rect 1409 22525 1443 22559
rect 1961 22525 1995 22559
rect 24593 22389 24627 22423
rect 23765 22185 23799 22219
rect 23581 22049 23615 22083
rect 24593 22049 24627 22083
rect 24777 21913 24811 21947
rect 24777 21641 24811 21675
rect 23857 21437 23891 21471
rect 24593 21437 24627 21471
rect 25145 21437 25179 21471
rect 24409 21301 24443 21335
rect 1777 21097 1811 21131
rect 1593 20961 1627 20995
rect 1593 20553 1627 20587
rect 13369 20417 13403 20451
rect 1409 20349 1443 20383
rect 13277 20281 13311 20315
rect 13636 20281 13670 20315
rect 1961 20213 1995 20247
rect 2421 20213 2455 20247
rect 14749 20213 14783 20247
rect 1593 20009 1627 20043
rect 1409 19873 1443 19907
rect 13369 19669 13403 19703
rect 1409 19261 1443 19295
rect 13553 19261 13587 19295
rect 2421 19193 2455 19227
rect 13820 19193 13854 19227
rect 1593 19125 1627 19159
rect 2053 19125 2087 19159
rect 13369 19125 13403 19159
rect 14933 19125 14967 19159
rect 1777 18921 1811 18955
rect 1593 18785 1627 18819
rect 12817 18785 12851 18819
rect 12909 18717 12943 18751
rect 13093 18717 13127 18751
rect 14013 18717 14047 18751
rect 12449 18649 12483 18683
rect 12357 18581 12391 18615
rect 13645 18581 13679 18615
rect 1593 18377 1627 18411
rect 2421 18377 2455 18411
rect 11529 18377 11563 18411
rect 1409 18173 1443 18207
rect 12449 18173 12483 18207
rect 12716 18105 12750 18139
rect 2053 18037 2087 18071
rect 11805 18037 11839 18071
rect 12265 18037 12299 18071
rect 13829 18037 13863 18071
rect 1593 17833 1627 17867
rect 13553 17833 13587 17867
rect 13921 17833 13955 17867
rect 14657 17833 14691 17867
rect 24777 17833 24811 17867
rect 1409 17697 1443 17731
rect 11325 17697 11359 17731
rect 24593 17697 24627 17731
rect 11069 17629 11103 17663
rect 14013 17629 14047 17663
rect 14105 17629 14139 17663
rect 15301 17629 15335 17663
rect 12449 17561 12483 17595
rect 13093 17561 13127 17595
rect 10793 17493 10827 17527
rect 13369 17493 13403 17527
rect 1593 17289 1627 17323
rect 2329 17289 2363 17323
rect 12449 17289 12483 17323
rect 24777 17289 24811 17323
rect 14197 17221 14231 17255
rect 11161 17153 11195 17187
rect 11345 17153 11379 17187
rect 13001 17153 13035 17187
rect 14381 17153 14415 17187
rect 1409 17085 1443 17119
rect 10609 17085 10643 17119
rect 12909 17085 12943 17119
rect 24593 17085 24627 17119
rect 25145 17085 25179 17119
rect 9873 17017 9907 17051
rect 14648 17017 14682 17051
rect 2053 16949 2087 16983
rect 10149 16949 10183 16983
rect 10701 16949 10735 16983
rect 11069 16949 11103 16983
rect 11713 16949 11747 16983
rect 12265 16949 12299 16983
rect 12817 16949 12851 16983
rect 13553 16949 13587 16983
rect 15761 16949 15795 16983
rect 24409 16949 24443 16983
rect 1593 16745 1627 16779
rect 11897 16745 11931 16779
rect 12541 16745 12575 16779
rect 13001 16745 13035 16779
rect 14013 16745 14047 16779
rect 15025 16745 15059 16779
rect 17049 16745 17083 16779
rect 23765 16745 23799 16779
rect 24777 16745 24811 16779
rect 14381 16677 14415 16711
rect 1409 16609 1443 16643
rect 10773 16609 10807 16643
rect 13369 16609 13403 16643
rect 15669 16609 15703 16643
rect 16865 16609 16899 16643
rect 23581 16609 23615 16643
rect 24593 16609 24627 16643
rect 10517 16541 10551 16575
rect 13461 16541 13495 16575
rect 13645 16541 13679 16575
rect 15761 16541 15795 16575
rect 15853 16541 15887 16575
rect 12909 16473 12943 16507
rect 15301 16473 15335 16507
rect 8769 16405 8803 16439
rect 10333 16405 10367 16439
rect 2697 16201 2731 16235
rect 10241 16201 10275 16235
rect 14289 16201 14323 16235
rect 14749 16201 14783 16235
rect 16773 16201 16807 16235
rect 24685 16201 24719 16235
rect 1593 16133 1627 16167
rect 9781 16133 9815 16167
rect 13277 16133 13311 16167
rect 18245 16133 18279 16167
rect 9229 16065 9263 16099
rect 10701 16065 10735 16099
rect 10793 16065 10827 16099
rect 13921 16065 13955 16099
rect 14841 16065 14875 16099
rect 1409 15997 1443 16031
rect 2505 15997 2539 16031
rect 10149 15997 10183 16031
rect 15108 15997 15142 16031
rect 18061 15997 18095 16031
rect 18521 15997 18555 16031
rect 23857 15997 23891 16031
rect 3065 15929 3099 15963
rect 8585 15929 8619 15963
rect 10609 15929 10643 15963
rect 11621 15929 11655 15963
rect 12725 15929 12759 15963
rect 13645 15929 13679 15963
rect 2053 15861 2087 15895
rect 2421 15861 2455 15895
rect 8217 15861 8251 15895
rect 8677 15861 8711 15895
rect 9045 15861 9079 15895
rect 9137 15861 9171 15895
rect 11253 15861 11287 15895
rect 12173 15861 12207 15895
rect 13093 15861 13127 15895
rect 13737 15861 13771 15895
rect 16221 15861 16255 15895
rect 17141 15861 17175 15895
rect 24225 15861 24259 15895
rect 1593 15657 1627 15691
rect 7941 15657 7975 15691
rect 8401 15657 8435 15691
rect 14105 15657 14139 15691
rect 14841 15657 14875 15691
rect 16313 15657 16347 15691
rect 19625 15657 19659 15691
rect 24777 15657 24811 15691
rect 10609 15589 10643 15623
rect 10946 15589 10980 15623
rect 12633 15589 12667 15623
rect 15669 15589 15703 15623
rect 1409 15521 1443 15555
rect 8493 15521 8527 15555
rect 14013 15521 14047 15555
rect 15761 15521 15795 15555
rect 17233 15521 17267 15555
rect 18429 15521 18463 15555
rect 19441 15521 19475 15555
rect 23581 15521 23615 15555
rect 24593 15521 24627 15555
rect 8585 15453 8619 15487
rect 9689 15453 9723 15487
rect 10701 15453 10735 15487
rect 13277 15453 13311 15487
rect 14289 15453 14323 15487
rect 15853 15453 15887 15487
rect 17325 15453 17359 15487
rect 17417 15453 17451 15487
rect 22569 15453 22603 15487
rect 8033 15385 8067 15419
rect 13645 15385 13679 15419
rect 4261 15317 4295 15351
rect 12081 15317 12115 15351
rect 15301 15317 15335 15351
rect 16773 15317 16807 15351
rect 16865 15317 16899 15351
rect 18613 15317 18647 15351
rect 23765 15317 23799 15351
rect 2053 15113 2087 15147
rect 7481 15113 7515 15147
rect 9873 15113 9907 15147
rect 13553 15113 13587 15147
rect 13921 15113 13955 15147
rect 16037 15113 16071 15147
rect 16405 15113 16439 15147
rect 17325 15113 17359 15147
rect 24777 15113 24811 15147
rect 10793 15045 10827 15079
rect 19349 15045 19383 15079
rect 3801 14977 3835 15011
rect 4445 14977 4479 15011
rect 11345 14977 11379 15011
rect 11897 14977 11931 15011
rect 13001 14977 13035 15011
rect 14013 14977 14047 15011
rect 1869 14909 1903 14943
rect 4261 14909 4295 14943
rect 7941 14909 7975 14943
rect 11161 14909 11195 14943
rect 16497 14909 16531 14943
rect 19165 14909 19199 14943
rect 19625 14909 19659 14943
rect 20361 14909 20395 14943
rect 20821 14909 20855 14943
rect 22569 14909 22603 14943
rect 24593 14909 24627 14943
rect 25145 14909 25179 14943
rect 4353 14841 4387 14875
rect 8208 14841 8242 14875
rect 10241 14841 10275 14875
rect 12265 14841 12299 14875
rect 12817 14841 12851 14875
rect 12909 14841 12943 14875
rect 14258 14841 14292 14875
rect 16957 14841 16991 14875
rect 18521 14841 18555 14875
rect 19993 14841 20027 14875
rect 1685 14773 1719 14807
rect 2513 14773 2547 14807
rect 3341 14773 3375 14807
rect 3893 14773 3927 14807
rect 6929 14773 6963 14807
rect 7757 14773 7791 14807
rect 9321 14773 9355 14807
rect 10701 14773 10735 14807
rect 11253 14773 11287 14807
rect 12449 14773 12483 14807
rect 15393 14773 15427 14807
rect 16681 14773 16715 14807
rect 17693 14773 17727 14807
rect 18061 14773 18095 14807
rect 20545 14773 20579 14807
rect 21557 14773 21591 14807
rect 22753 14773 22787 14807
rect 23121 14773 23155 14807
rect 23949 14773 23983 14807
rect 24409 14773 24443 14807
rect 1593 14569 1627 14603
rect 2697 14569 2731 14603
rect 4077 14569 4111 14603
rect 11069 14569 11103 14603
rect 11621 14569 11655 14603
rect 13737 14569 13771 14603
rect 14657 14569 14691 14603
rect 15025 14569 15059 14603
rect 15761 14569 15795 14603
rect 17325 14569 17359 14603
rect 18613 14569 18647 14603
rect 24777 14569 24811 14603
rect 5886 14501 5920 14535
rect 14105 14501 14139 14535
rect 15669 14501 15703 14535
rect 1409 14433 1443 14467
rect 2421 14433 2455 14467
rect 2513 14433 2547 14467
rect 4445 14433 4479 14467
rect 4537 14433 4571 14467
rect 5641 14433 5675 14467
rect 9956 14433 9990 14467
rect 12541 14433 12575 14467
rect 14197 14433 14231 14467
rect 17233 14433 17267 14467
rect 18429 14433 18463 14467
rect 19533 14433 19567 14467
rect 20913 14433 20947 14467
rect 22569 14433 22603 14467
rect 23581 14433 23615 14467
rect 24593 14433 24627 14467
rect 4721 14365 4755 14399
rect 8217 14365 8251 14399
rect 9689 14365 9723 14399
rect 12633 14365 12667 14399
rect 12725 14365 12759 14399
rect 13277 14365 13311 14399
rect 15853 14365 15887 14399
rect 17417 14365 17451 14399
rect 3801 14297 3835 14331
rect 5089 14297 5123 14331
rect 8033 14297 8067 14331
rect 15301 14297 15335 14331
rect 1961 14229 1995 14263
rect 3157 14229 3191 14263
rect 3433 14229 3467 14263
rect 7021 14229 7055 14263
rect 8677 14229 8711 14263
rect 11989 14229 12023 14263
rect 12173 14229 12207 14263
rect 14381 14229 14415 14263
rect 16405 14229 16439 14263
rect 16681 14229 16715 14263
rect 16865 14229 16899 14263
rect 18153 14229 18187 14263
rect 19073 14229 19107 14263
rect 19717 14229 19751 14263
rect 21097 14229 21131 14263
rect 22753 14229 22787 14263
rect 23765 14229 23799 14263
rect 2329 14025 2363 14059
rect 3801 14025 3835 14059
rect 5641 14025 5675 14059
rect 6561 14025 6595 14059
rect 9689 14025 9723 14059
rect 10517 14025 10551 14059
rect 12265 14025 12299 14059
rect 15393 14025 15427 14059
rect 15761 14025 15795 14059
rect 17233 14025 17267 14059
rect 18061 14025 18095 14059
rect 19441 14025 19475 14059
rect 21189 14025 21223 14059
rect 23397 14025 23431 14059
rect 1593 13957 1627 13991
rect 4169 13957 4203 13991
rect 12633 13957 12667 13991
rect 16129 13957 16163 13991
rect 24777 13957 24811 13991
rect 4261 13889 4295 13923
rect 9413 13889 9447 13923
rect 10977 13889 11011 13923
rect 11161 13889 11195 13923
rect 11805 13889 11839 13923
rect 16681 13889 16715 13923
rect 18613 13889 18647 13923
rect 19073 13889 19107 13923
rect 1409 13821 1443 13855
rect 2053 13821 2087 13855
rect 2513 13821 2547 13855
rect 2973 13821 3007 13855
rect 4517 13821 4551 13855
rect 6285 13821 6319 13855
rect 7113 13821 7147 13855
rect 7205 13821 7239 13855
rect 7461 13821 7495 13855
rect 10057 13821 10091 13855
rect 13093 13821 13127 13855
rect 13360 13821 13394 13855
rect 16589 13821 16623 13855
rect 17601 13821 17635 13855
rect 18521 13821 18555 13855
rect 20177 13821 20211 13855
rect 21005 13821 21039 13855
rect 21833 13821 21867 13855
rect 22569 13821 22603 13855
rect 23029 13821 23063 13855
rect 23857 13821 23891 13855
rect 24593 13821 24627 13855
rect 25145 13821 25179 13855
rect 10885 13753 10919 13787
rect 16497 13753 16531 13787
rect 19625 13753 19659 13787
rect 2697 13685 2731 13719
rect 3433 13685 3467 13719
rect 8585 13685 8619 13719
rect 14473 13685 14507 13719
rect 18429 13685 18463 13719
rect 21465 13685 21499 13719
rect 22753 13685 22787 13719
rect 24409 13685 24443 13719
rect 2053 13481 2087 13515
rect 5641 13481 5675 13515
rect 7297 13481 7331 13515
rect 7573 13481 7607 13515
rect 10149 13481 10183 13515
rect 10793 13481 10827 13515
rect 12265 13481 12299 13515
rect 13093 13481 13127 13515
rect 13553 13481 13587 13515
rect 14565 13481 14599 13515
rect 15117 13481 15151 13515
rect 15853 13481 15887 13515
rect 17417 13481 17451 13515
rect 23765 13481 23799 13515
rect 24777 13481 24811 13515
rect 8033 13413 8067 13447
rect 12357 13413 12391 13447
rect 1409 13345 1443 13379
rect 2513 13345 2547 13379
rect 3433 13345 3467 13379
rect 4261 13345 4295 13379
rect 4528 13345 4562 13379
rect 6929 13345 6963 13379
rect 7941 13345 7975 13379
rect 10057 13345 10091 13379
rect 13921 13345 13955 13379
rect 14013 13345 14047 13379
rect 16293 13345 16327 13379
rect 18889 13345 18923 13379
rect 23581 13345 23615 13379
rect 24593 13345 24627 13379
rect 8125 13277 8159 13311
rect 10241 13277 10275 13311
rect 12541 13277 12575 13311
rect 14197 13277 14231 13311
rect 16037 13277 16071 13311
rect 18981 13277 19015 13311
rect 19073 13277 19107 13311
rect 20913 13277 20947 13311
rect 22569 13277 22603 13311
rect 2421 13209 2455 13243
rect 11897 13209 11931 13243
rect 1593 13141 1627 13175
rect 2697 13141 2731 13175
rect 3065 13141 3099 13175
rect 3893 13141 3927 13175
rect 8585 13141 8619 13175
rect 9413 13141 9447 13175
rect 9689 13141 9723 13175
rect 11345 13141 11379 13175
rect 11805 13141 11839 13175
rect 15577 13141 15611 13175
rect 18153 13141 18187 13175
rect 18521 13141 18555 13175
rect 19625 13141 19659 13175
rect 20085 13141 20119 13175
rect 1593 12937 1627 12971
rect 3065 12937 3099 12971
rect 6653 12937 6687 12971
rect 8125 12937 8159 12971
rect 9137 12937 9171 12971
rect 9505 12937 9539 12971
rect 11161 12937 11195 12971
rect 11989 12937 12023 12971
rect 13645 12937 13679 12971
rect 14657 12937 14691 12971
rect 15209 12937 15243 12971
rect 16221 12937 16255 12971
rect 16589 12937 16623 12971
rect 16957 12937 16991 12971
rect 19625 12937 19659 12971
rect 20729 12937 20763 12971
rect 21005 12937 21039 12971
rect 23857 12937 23891 12971
rect 24777 12937 24811 12971
rect 4629 12869 4663 12903
rect 22753 12869 22787 12903
rect 24409 12869 24443 12903
rect 3525 12801 3559 12835
rect 3617 12801 3651 12835
rect 5181 12801 5215 12835
rect 5641 12801 5675 12835
rect 8677 12801 8711 12835
rect 10241 12801 10275 12835
rect 14289 12801 14323 12835
rect 15761 12801 15795 12835
rect 17509 12801 17543 12835
rect 18613 12801 18647 12835
rect 20177 12801 20211 12835
rect 1409 12733 1443 12767
rect 2053 12733 2087 12767
rect 3433 12733 3467 12767
rect 7113 12733 7147 12767
rect 7665 12733 7699 12767
rect 8493 12733 8527 12767
rect 11345 12733 11379 12767
rect 12633 12733 12667 12767
rect 13553 12733 13587 12767
rect 14013 12733 14047 12767
rect 16773 12733 16807 12767
rect 18521 12733 18555 12767
rect 22569 12733 22603 12767
rect 23029 12733 23063 12767
rect 24593 12733 24627 12767
rect 25145 12733 25179 12767
rect 2329 12665 2363 12699
rect 2973 12665 3007 12699
rect 4537 12665 4571 12699
rect 4997 12665 5031 12699
rect 5089 12665 5123 12699
rect 15117 12665 15151 12699
rect 15577 12665 15611 12699
rect 17785 12665 17819 12699
rect 19073 12665 19107 12699
rect 19533 12665 19567 12699
rect 19993 12665 20027 12699
rect 4169 12597 4203 12631
rect 7297 12597 7331 12631
rect 8033 12597 8067 12631
rect 8585 12597 8619 12631
rect 9689 12597 9723 12631
rect 10057 12597 10091 12631
rect 10149 12597 10183 12631
rect 10701 12597 10735 12631
rect 11529 12597 11563 12631
rect 12817 12597 12851 12631
rect 13185 12597 13219 12631
rect 14105 12597 14139 12631
rect 15669 12597 15703 12631
rect 18061 12597 18095 12631
rect 18429 12597 18463 12631
rect 20085 12597 20119 12631
rect 21189 12597 21223 12631
rect 2421 12393 2455 12427
rect 2789 12393 2823 12427
rect 4261 12393 4295 12427
rect 7757 12393 7791 12427
rect 8861 12393 8895 12427
rect 11805 12393 11839 12427
rect 12449 12393 12483 12427
rect 14197 12393 14231 12427
rect 14565 12393 14599 12427
rect 15301 12393 15335 12427
rect 15853 12393 15887 12427
rect 18521 12393 18555 12427
rect 19073 12393 19107 12427
rect 21833 12393 21867 12427
rect 24777 12393 24811 12427
rect 4813 12325 4847 12359
rect 7665 12325 7699 12359
rect 10692 12325 10726 12359
rect 13645 12325 13679 12359
rect 14933 12325 14967 12359
rect 1409 12257 1443 12291
rect 2881 12257 2915 12291
rect 5641 12257 5675 12291
rect 8125 12257 8159 12291
rect 13553 12257 13587 12291
rect 16856 12257 16890 12291
rect 19441 12257 19475 12291
rect 20453 12257 20487 12291
rect 22017 12257 22051 12291
rect 22284 12257 22318 12291
rect 24593 12257 24627 12291
rect 2329 12189 2363 12223
rect 3065 12189 3099 12223
rect 5733 12189 5767 12223
rect 5917 12189 5951 12223
rect 8217 12189 8251 12223
rect 8309 12189 8343 12223
rect 9505 12189 9539 12223
rect 10241 12189 10275 12223
rect 10425 12189 10459 12223
rect 13093 12189 13127 12223
rect 13829 12189 13863 12223
rect 16589 12189 16623 12223
rect 19533 12189 19567 12223
rect 19625 12189 19659 12223
rect 20913 12189 20947 12223
rect 1593 12121 1627 12155
rect 5273 12121 5307 12155
rect 13185 12121 13219 12155
rect 20085 12121 20119 12155
rect 1961 12053 1995 12087
rect 3433 12053 3467 12087
rect 3893 12053 3927 12087
rect 5181 12053 5215 12087
rect 6285 12053 6319 12087
rect 6653 12053 6687 12087
rect 7205 12053 7239 12087
rect 9965 12053 9999 12087
rect 16129 12053 16163 12087
rect 17969 12053 18003 12087
rect 18981 12053 19015 12087
rect 21465 12053 21499 12087
rect 23397 12053 23431 12087
rect 24041 12053 24075 12087
rect 2237 11849 2271 11883
rect 3341 11849 3375 11883
rect 5181 11849 5215 11883
rect 6469 11849 6503 11883
rect 9689 11849 9723 11883
rect 10609 11849 10643 11883
rect 13185 11849 13219 11883
rect 16129 11849 16163 11883
rect 17509 11849 17543 11883
rect 22845 11849 22879 11883
rect 23397 11849 23431 11883
rect 1777 11781 1811 11815
rect 2789 11713 2823 11747
rect 10333 11713 10367 11747
rect 15025 11781 15059 11815
rect 11345 11713 11379 11747
rect 15669 11713 15703 11747
rect 16773 11713 16807 11747
rect 22385 11713 22419 11747
rect 23673 11713 23707 11747
rect 3709 11645 3743 11679
rect 3801 11645 3835 11679
rect 7205 11645 7239 11679
rect 7297 11645 7331 11679
rect 7564 11645 7598 11679
rect 9505 11645 9539 11679
rect 2697 11577 2731 11611
rect 4068 11577 4102 11611
rect 5825 11577 5859 11611
rect 10609 11645 10643 11679
rect 13645 11645 13679 11679
rect 13912 11645 13946 11679
rect 16589 11645 16623 11679
rect 19349 11645 19383 11679
rect 21373 11645 21407 11679
rect 10149 11577 10183 11611
rect 10793 11577 10827 11611
rect 19594 11577 19628 11611
rect 21649 11577 21683 11611
rect 22201 11577 22235 11611
rect 23940 11577 23974 11611
rect 2145 11509 2179 11543
rect 2605 11509 2639 11543
rect 6193 11509 6227 11543
rect 8677 11509 8711 11543
rect 9321 11509 9355 11543
rect 9505 11509 9539 11543
rect 9781 11509 9815 11543
rect 10241 11509 10275 11543
rect 10609 11509 10643 11543
rect 11253 11509 11287 11543
rect 11805 11509 11839 11543
rect 12173 11509 12207 11543
rect 12633 11509 12667 11543
rect 15945 11509 15979 11543
rect 16497 11509 16531 11543
rect 17233 11509 17267 11543
rect 18153 11509 18187 11543
rect 18797 11509 18831 11543
rect 19257 11509 19291 11543
rect 20729 11509 20763 11543
rect 21833 11509 21867 11543
rect 22293 11509 22327 11543
rect 25053 11509 25087 11543
rect 1593 11305 1627 11339
rect 2329 11305 2363 11339
rect 2697 11305 2731 11339
rect 4077 11305 4111 11339
rect 4445 11305 4479 11339
rect 7021 11305 7055 11339
rect 7389 11305 7423 11339
rect 8033 11305 8067 11339
rect 9689 11305 9723 11339
rect 12081 11305 12115 11339
rect 13001 11305 13035 11339
rect 13185 11305 13219 11339
rect 14657 11305 14691 11339
rect 15117 11305 15151 11339
rect 16681 11305 16715 11339
rect 17233 11305 17267 11339
rect 19441 11305 19475 11339
rect 20729 11305 20763 11339
rect 22293 11305 22327 11339
rect 23397 11305 23431 11339
rect 23857 11305 23891 11339
rect 25237 11305 25271 11339
rect 4537 11237 4571 11271
rect 7849 11237 7883 11271
rect 8401 11237 8435 11271
rect 9137 11237 9171 11271
rect 10946 11237 10980 11271
rect 12725 11237 12759 11271
rect 13553 11237 13587 11271
rect 15546 11237 15580 11271
rect 23949 11237 23983 11271
rect 1409 11169 1443 11203
rect 2501 11169 2535 11203
rect 6009 11169 6043 11203
rect 8493 11169 8527 11203
rect 13645 11169 13679 11203
rect 18328 11169 18362 11203
rect 20913 11169 20947 11203
rect 21169 11169 21203 11203
rect 25053 11169 25087 11203
rect 4629 11101 4663 11135
rect 6101 11101 6135 11135
rect 6193 11101 6227 11135
rect 8677 11101 8711 11135
rect 10701 11101 10735 11135
rect 13829 11101 13863 11135
rect 14289 11101 14323 11135
rect 15301 11101 15335 11135
rect 18061 11101 18095 11135
rect 24041 11101 24075 11135
rect 24593 11101 24627 11135
rect 3433 11033 3467 11067
rect 3893 11033 3927 11067
rect 5549 11033 5583 11067
rect 9505 11033 9539 11067
rect 10241 11033 10275 11067
rect 20361 11033 20395 11067
rect 23029 11033 23063 11067
rect 3157 10965 3191 10999
rect 5181 10965 5215 10999
rect 5641 10965 5675 10999
rect 10609 10965 10643 10999
rect 17969 10965 18003 10999
rect 23489 10965 23523 10999
rect 1593 10761 1627 10795
rect 3985 10761 4019 10795
rect 4629 10761 4663 10795
rect 6469 10761 6503 10795
rect 8953 10761 8987 10795
rect 13553 10761 13587 10795
rect 14197 10761 14231 10795
rect 16865 10761 16899 10795
rect 18245 10761 18279 10795
rect 20637 10761 20671 10795
rect 22661 10761 22695 10795
rect 24685 10761 24719 10795
rect 25053 10761 25087 10795
rect 25421 10761 25455 10795
rect 10333 10693 10367 10727
rect 20545 10693 20579 10727
rect 2053 10625 2087 10659
rect 5733 10625 5767 10659
rect 10241 10625 10275 10659
rect 10885 10625 10919 10659
rect 11897 10625 11931 10659
rect 11989 10625 12023 10659
rect 12265 10625 12299 10659
rect 13001 10625 13035 10659
rect 17509 10625 17543 10659
rect 18797 10625 18831 10659
rect 21097 10625 21131 10659
rect 21281 10625 21315 10659
rect 24317 10625 24351 10659
rect 1409 10557 1443 10591
rect 2605 10557 2639 10591
rect 4997 10557 5031 10591
rect 5457 10557 5491 10591
rect 7573 10557 7607 10591
rect 7840 10557 7874 10591
rect 10701 10557 10735 10591
rect 12817 10557 12851 10591
rect 15025 10557 15059 10591
rect 15485 10557 15519 10591
rect 15752 10557 15786 10591
rect 21005 10557 21039 10591
rect 22477 10557 22511 10591
rect 23029 10557 23063 10591
rect 24041 10557 24075 10591
rect 25237 10557 25271 10591
rect 25789 10557 25823 10591
rect 2872 10489 2906 10523
rect 7113 10489 7147 10523
rect 11989 10489 12023 10523
rect 12909 10489 12943 10523
rect 13921 10489 13955 10523
rect 18613 10489 18647 10523
rect 19625 10489 19659 10523
rect 21741 10489 21775 10523
rect 23489 10489 23523 10523
rect 24133 10489 24167 10523
rect 2329 10421 2363 10455
rect 5089 10421 5123 10455
rect 5549 10421 5583 10455
rect 6193 10421 6227 10455
rect 7481 10421 7515 10455
rect 9597 10421 9631 10455
rect 10793 10421 10827 10455
rect 11345 10421 11379 10455
rect 12449 10421 12483 10455
rect 14473 10421 14507 10455
rect 15393 10421 15427 10455
rect 17785 10421 17819 10455
rect 18705 10421 18739 10455
rect 19349 10421 19383 10455
rect 20177 10421 20211 10455
rect 22385 10421 22419 10455
rect 23673 10421 23707 10455
rect 2421 10217 2455 10251
rect 7573 10217 7607 10251
rect 8677 10217 8711 10251
rect 9321 10217 9355 10251
rect 11161 10217 11195 10251
rect 11621 10217 11655 10251
rect 14473 10217 14507 10251
rect 15117 10217 15151 10251
rect 18153 10217 18187 10251
rect 20545 10217 20579 10251
rect 20913 10217 20947 10251
rect 21281 10217 21315 10251
rect 21373 10217 21407 10251
rect 22109 10217 22143 10251
rect 23121 10217 23155 10251
rect 2329 10149 2363 10183
rect 8953 10149 8987 10183
rect 13185 10149 13219 10183
rect 15761 10149 15795 10183
rect 18061 10149 18095 10183
rect 18521 10149 18555 10183
rect 22845 10149 22879 10183
rect 1409 10081 1443 10115
rect 2789 10081 2823 10115
rect 3525 10081 3559 10115
rect 4537 10081 4571 10115
rect 4804 10081 4838 10115
rect 7941 10081 7975 10115
rect 8033 10081 8067 10115
rect 11069 10081 11103 10115
rect 11529 10081 11563 10115
rect 13093 10081 13127 10115
rect 15669 10081 15703 10115
rect 18613 10081 18647 10115
rect 19809 10081 19843 10115
rect 23572 10081 23606 10115
rect 2881 10013 2915 10047
rect 3065 10013 3099 10047
rect 8217 10013 8251 10047
rect 10149 10013 10183 10047
rect 11713 10013 11747 10047
rect 13277 10013 13311 10047
rect 15853 10013 15887 10047
rect 16681 10013 16715 10047
rect 17141 10013 17175 10047
rect 18705 10013 18739 10047
rect 21465 10013 21499 10047
rect 23305 10013 23339 10047
rect 1869 9945 1903 9979
rect 3801 9945 3835 9979
rect 7481 9945 7515 9979
rect 12725 9945 12759 9979
rect 15301 9945 15335 9979
rect 19993 9945 20027 9979
rect 1593 9877 1627 9911
rect 4445 9877 4479 9911
rect 5917 9877 5951 9911
rect 6469 9877 6503 9911
rect 6929 9877 6963 9911
rect 9965 9877 9999 9911
rect 10701 9877 10735 9911
rect 12541 9877 12575 9911
rect 13829 9877 13863 9911
rect 14105 9877 14139 9911
rect 16405 9877 16439 9911
rect 17601 9877 17635 9911
rect 24685 9877 24719 9911
rect 9321 9673 9355 9707
rect 13461 9673 13495 9707
rect 19441 9673 19475 9707
rect 19993 9673 20027 9707
rect 20361 9673 20395 9707
rect 21465 9673 21499 9707
rect 23305 9673 23339 9707
rect 1593 9605 1627 9639
rect 2421 9605 2455 9639
rect 2789 9605 2823 9639
rect 4353 9605 4387 9639
rect 10517 9605 10551 9639
rect 12173 9605 12207 9639
rect 12449 9605 12483 9639
rect 14289 9605 14323 9639
rect 17141 9605 17175 9639
rect 17509 9605 17543 9639
rect 17785 9605 17819 9639
rect 20729 9605 20763 9639
rect 23673 9605 23707 9639
rect 25421 9605 25455 9639
rect 3433 9537 3467 9571
rect 4997 9537 5031 9571
rect 6653 9537 6687 9571
rect 11069 9537 11103 9571
rect 13001 9537 13035 9571
rect 14013 9537 14047 9571
rect 15025 9537 15059 9571
rect 16681 9537 16715 9571
rect 18061 9537 18095 9571
rect 21189 9537 21223 9571
rect 22477 9537 22511 9571
rect 22661 9537 22695 9571
rect 24317 9537 24351 9571
rect 1409 9469 1443 9503
rect 2421 9469 2455 9503
rect 2513 9469 2547 9503
rect 3157 9469 3191 9503
rect 4813 9469 4847 9503
rect 7941 9469 7975 9503
rect 8208 9469 8242 9503
rect 12817 9469 12851 9503
rect 12909 9469 12943 9503
rect 14841 9469 14875 9503
rect 15577 9469 15611 9503
rect 20545 9469 20579 9503
rect 21925 9469 21959 9503
rect 22385 9469 22419 9503
rect 24041 9469 24075 9503
rect 25237 9469 25271 9503
rect 25789 9469 25823 9503
rect 2329 9401 2363 9435
rect 3801 9401 3835 9435
rect 4261 9401 4295 9435
rect 4721 9401 4755 9435
rect 6837 9401 6871 9435
rect 10977 9401 11011 9435
rect 14933 9401 14967 9435
rect 16497 9401 16531 9435
rect 18306 9401 18340 9435
rect 24133 9401 24167 9435
rect 25053 9401 25087 9435
rect 2513 9333 2547 9367
rect 2605 9333 2639 9367
rect 3249 9333 3283 9367
rect 5365 9333 5399 9367
rect 5733 9333 5767 9367
rect 6193 9333 6227 9367
rect 7573 9333 7607 9367
rect 9965 9333 9999 9367
rect 10333 9333 10367 9367
rect 10885 9333 10919 9367
rect 11621 9333 11655 9367
rect 14473 9333 14507 9367
rect 15853 9333 15887 9367
rect 16037 9333 16071 9367
rect 16405 9333 16439 9367
rect 22017 9333 22051 9367
rect 24777 9333 24811 9367
rect 1593 9129 1627 9163
rect 2329 9129 2363 9163
rect 7205 9129 7239 9163
rect 8953 9129 8987 9163
rect 11621 9129 11655 9163
rect 12449 9129 12483 9163
rect 15025 9129 15059 9163
rect 16681 9129 16715 9163
rect 17601 9129 17635 9163
rect 18061 9129 18095 9163
rect 20269 9129 20303 9163
rect 21281 9129 21315 9163
rect 21373 9129 21407 9163
rect 22109 9129 22143 9163
rect 23305 9129 23339 9163
rect 2789 9061 2823 9095
rect 7665 9061 7699 9095
rect 15568 9061 15602 9095
rect 24032 9061 24066 9095
rect 1409 8993 1443 9027
rect 4344 8993 4378 9027
rect 7573 8993 7607 9027
rect 8309 8993 8343 9027
rect 10508 8993 10542 9027
rect 12992 8993 13026 9027
rect 15301 8993 15335 9027
rect 18429 8993 18463 9027
rect 19717 8993 19751 9027
rect 23765 8993 23799 9027
rect 2881 8925 2915 8959
rect 2973 8925 3007 8959
rect 4077 8925 4111 8959
rect 7757 8925 7791 8959
rect 8677 8925 8711 8959
rect 10241 8925 10275 8959
rect 12725 8925 12759 8959
rect 18521 8925 18555 8959
rect 18613 8925 18647 8959
rect 20729 8925 20763 8959
rect 21465 8925 21499 8959
rect 22753 8925 22787 8959
rect 2421 8857 2455 8891
rect 9321 8857 9355 8891
rect 14749 8857 14783 8891
rect 1961 8789 1995 8823
rect 3433 8789 3467 8823
rect 3893 8789 3927 8823
rect 5457 8789 5491 8823
rect 6009 8789 6043 8823
rect 6377 8789 6411 8823
rect 7113 8789 7147 8823
rect 9873 8789 9907 8823
rect 14105 8789 14139 8823
rect 17969 8789 18003 8823
rect 19073 8789 19107 8823
rect 19441 8789 19475 8823
rect 19901 8789 19935 8823
rect 20913 8789 20947 8823
rect 25145 8789 25179 8823
rect 2145 8585 2179 8619
rect 5181 8585 5215 8619
rect 7205 8585 7239 8619
rect 10149 8585 10183 8619
rect 11069 8585 11103 8619
rect 17509 8585 17543 8619
rect 19441 8585 19475 8619
rect 20177 8585 20211 8619
rect 20545 8585 20579 8619
rect 24869 8585 24903 8619
rect 25237 8585 25271 8619
rect 25605 8585 25639 8619
rect 4261 8517 4295 8551
rect 8585 8517 8619 8551
rect 16405 8517 16439 8551
rect 17877 8517 17911 8551
rect 22017 8517 22051 8551
rect 1777 8449 1811 8483
rect 5825 8449 5859 8483
rect 6193 8449 6227 8483
rect 7757 8449 7791 8483
rect 8309 8449 8343 8483
rect 10701 8449 10735 8483
rect 11897 8449 11931 8483
rect 24501 8449 24535 8483
rect 2237 8381 2271 8415
rect 5549 8381 5583 8415
rect 8769 8381 8803 8415
rect 12173 8381 12207 8415
rect 12449 8381 12483 8415
rect 12716 8381 12750 8415
rect 15025 8381 15059 8415
rect 18061 8381 18095 8415
rect 20637 8381 20671 8415
rect 23121 8381 23155 8415
rect 24317 8381 24351 8415
rect 25421 8381 25455 8415
rect 25973 8381 26007 8415
rect 2482 8313 2516 8347
rect 4537 8313 4571 8347
rect 5089 8313 5123 8347
rect 5641 8313 5675 8347
rect 6561 8313 6595 8347
rect 7665 8313 7699 8347
rect 9014 8313 9048 8347
rect 14565 8313 14599 8347
rect 15292 8313 15326 8347
rect 17141 8313 17175 8347
rect 18328 8313 18362 8347
rect 20882 8313 20916 8347
rect 23489 8313 23523 8347
rect 24225 8313 24259 8347
rect 3617 8245 3651 8279
rect 7021 8245 7055 8279
rect 7573 8245 7607 8279
rect 11253 8245 11287 8279
rect 13829 8245 13863 8279
rect 14841 8245 14875 8279
rect 22569 8245 22603 8279
rect 23857 8245 23891 8279
rect 2329 8041 2363 8075
rect 2789 8041 2823 8075
rect 5273 8041 5307 8075
rect 7849 8041 7883 8075
rect 10149 8041 10183 8075
rect 12081 8041 12115 8075
rect 12817 8041 12851 8075
rect 13093 8041 13127 8075
rect 13645 8041 13679 8075
rect 14013 8041 14047 8075
rect 14749 8041 14783 8075
rect 15117 8041 15151 8075
rect 16589 8041 16623 8075
rect 17693 8041 17727 8075
rect 18061 8041 18095 8075
rect 19165 8041 19199 8075
rect 19625 8041 19659 8075
rect 22293 8041 22327 8075
rect 22845 8041 22879 8075
rect 23765 8041 23799 8075
rect 2237 7973 2271 8007
rect 2697 7973 2731 8007
rect 8401 7973 8435 8007
rect 11621 7973 11655 8007
rect 14105 7973 14139 8007
rect 15485 7973 15519 8007
rect 18705 7973 18739 8007
rect 20361 7973 20395 8007
rect 21180 7973 21214 8007
rect 24216 7973 24250 8007
rect 5816 7905 5850 7939
rect 8493 7905 8527 7939
rect 10517 7905 10551 7939
rect 16497 7905 16531 7939
rect 17601 7905 17635 7939
rect 19717 7905 19751 7939
rect 23949 7905 23983 7939
rect 2881 7837 2915 7871
rect 4077 7837 4111 7871
rect 5549 7837 5583 7871
rect 8677 7837 8711 7871
rect 10609 7837 10643 7871
rect 10701 7837 10735 7871
rect 12173 7837 12207 7871
rect 12265 7837 12299 7871
rect 13553 7837 13587 7871
rect 14197 7837 14231 7871
rect 16773 7837 16807 7871
rect 18153 7837 18187 7871
rect 18245 7837 18279 7871
rect 19809 7837 19843 7871
rect 20729 7837 20763 7871
rect 20913 7837 20947 7871
rect 3709 7769 3743 7803
rect 16129 7769 16163 7803
rect 19257 7769 19291 7803
rect 1593 7701 1627 7735
rect 3341 7701 3375 7735
rect 4537 7701 4571 7735
rect 6929 7701 6963 7735
rect 7573 7701 7607 7735
rect 8033 7701 8067 7735
rect 9045 7701 9079 7735
rect 9413 7701 9447 7735
rect 10057 7701 10091 7735
rect 11253 7701 11287 7735
rect 11713 7701 11747 7735
rect 16037 7701 16071 7735
rect 17141 7701 17175 7735
rect 25329 7701 25363 7735
rect 1685 7497 1719 7531
rect 3525 7497 3559 7531
rect 5181 7497 5215 7531
rect 8217 7497 8251 7531
rect 10793 7497 10827 7531
rect 11805 7497 11839 7531
rect 12173 7497 12207 7531
rect 12725 7497 12759 7531
rect 13645 7497 13679 7531
rect 15209 7497 15243 7531
rect 15853 7497 15887 7531
rect 17417 7497 17451 7531
rect 18061 7497 18095 7531
rect 19349 7497 19383 7531
rect 22201 7497 22235 7531
rect 23673 7497 23707 7531
rect 24685 7497 24719 7531
rect 25145 7497 25179 7531
rect 25421 7497 25455 7531
rect 9689 7429 9723 7463
rect 16313 7429 16347 7463
rect 17785 7429 17819 7463
rect 20729 7429 20763 7463
rect 4445 7361 4479 7395
rect 5089 7361 5123 7395
rect 5825 7361 5859 7395
rect 10241 7361 10275 7395
rect 11345 7361 11379 7395
rect 13829 7361 13863 7395
rect 16865 7361 16899 7395
rect 18521 7361 18555 7395
rect 18705 7361 18739 7395
rect 21281 7361 21315 7395
rect 24133 7361 24167 7395
rect 24317 7361 24351 7395
rect 2053 7293 2087 7327
rect 2145 7293 2179 7327
rect 6193 7293 6227 7327
rect 6653 7293 6687 7327
rect 6837 7293 6871 7327
rect 10609 7293 10643 7327
rect 18429 7293 18463 7327
rect 19625 7293 19659 7327
rect 22293 7293 22327 7327
rect 23121 7293 23155 7327
rect 25237 7293 25271 7327
rect 25789 7293 25823 7327
rect 2390 7225 2424 7259
rect 5549 7225 5583 7259
rect 7104 7225 7138 7259
rect 9137 7225 9171 7259
rect 9781 7225 9815 7259
rect 11253 7225 11287 7259
rect 13369 7225 13403 7259
rect 14074 7225 14108 7259
rect 20177 7225 20211 7259
rect 21189 7225 21223 7259
rect 23489 7225 23523 7259
rect 24041 7225 24075 7259
rect 5641 7157 5675 7191
rect 8861 7157 8895 7191
rect 11161 7157 11195 7191
rect 12817 7157 12851 7191
rect 16129 7157 16163 7191
rect 16681 7157 16715 7191
rect 16773 7157 16807 7191
rect 19809 7157 19843 7191
rect 20637 7157 20671 7191
rect 21097 7157 21131 7191
rect 21741 7157 21775 7191
rect 22477 7157 22511 7191
rect 2421 6953 2455 6987
rect 2789 6953 2823 6987
rect 5641 6953 5675 6987
rect 5917 6953 5951 6987
rect 8309 6953 8343 6987
rect 12173 6953 12207 6987
rect 13185 6953 13219 6987
rect 13737 6953 13771 6987
rect 14749 6953 14783 6987
rect 15577 6953 15611 6987
rect 15945 6953 15979 6987
rect 18153 6953 18187 6987
rect 19993 6953 20027 6987
rect 20361 6953 20395 6987
rect 20729 6953 20763 6987
rect 22293 6953 22327 6987
rect 23673 6953 23707 6987
rect 3525 6885 3559 6919
rect 4721 6885 4755 6919
rect 8217 6885 8251 6919
rect 14381 6885 14415 6919
rect 24032 6885 24066 6919
rect 1409 6817 1443 6851
rect 6285 6817 6319 6851
rect 10241 6817 10275 6851
rect 10793 6817 10827 6851
rect 11049 6817 11083 6851
rect 16304 6817 16338 6851
rect 18889 6817 18923 6851
rect 21169 6817 21203 6851
rect 23765 6817 23799 6851
rect 2881 6749 2915 6783
rect 3065 6749 3099 6783
rect 4813 6749 4847 6783
rect 4905 6749 4939 6783
rect 6377 6749 6411 6783
rect 6561 6749 6595 6783
rect 8493 6749 8527 6783
rect 9781 6749 9815 6783
rect 13829 6749 13863 6783
rect 13921 6749 13955 6783
rect 16037 6749 16071 6783
rect 18981 6749 19015 6783
rect 19073 6749 19107 6783
rect 20913 6749 20947 6783
rect 1593 6681 1627 6715
rect 4353 6681 4387 6715
rect 7021 6681 7055 6715
rect 7389 6681 7423 6715
rect 7757 6681 7791 6715
rect 12909 6681 12943 6715
rect 2237 6613 2271 6647
rect 3801 6613 3835 6647
rect 7849 6613 7883 6647
rect 8861 6613 8895 6647
rect 9229 6613 9263 6647
rect 10701 6613 10735 6647
rect 13369 6613 13403 6647
rect 17417 6613 17451 6647
rect 18521 6613 18555 6647
rect 19625 6613 19659 6647
rect 22845 6613 22879 6647
rect 25145 6613 25179 6647
rect 2513 6409 2547 6443
rect 2789 6409 2823 6443
rect 3801 6409 3835 6443
rect 4077 6409 4111 6443
rect 6009 6409 6043 6443
rect 6285 6409 6319 6443
rect 9505 6409 9539 6443
rect 13369 6409 13403 6443
rect 15117 6409 15151 6443
rect 17509 6409 17543 6443
rect 17877 6409 17911 6443
rect 23121 6409 23155 6443
rect 23489 6409 23523 6443
rect 23949 6409 23983 6443
rect 2145 6341 2179 6375
rect 3249 6273 3283 6307
rect 3433 6273 3467 6307
rect 3157 6205 3191 6239
rect 4353 6341 4387 6375
rect 5365 6341 5399 6375
rect 10333 6341 10367 6375
rect 10425 6341 10459 6375
rect 11621 6341 11655 6375
rect 18705 6341 18739 6375
rect 4905 6273 4939 6307
rect 6837 6273 6871 6307
rect 11161 6273 11195 6307
rect 13737 6273 13771 6307
rect 16865 6273 16899 6307
rect 17049 6273 17083 6307
rect 22661 6273 22695 6307
rect 24133 6273 24167 6307
rect 4261 6205 4295 6239
rect 4721 6205 4755 6239
rect 8125 6205 8159 6239
rect 10333 6205 10367 6239
rect 11069 6205 11103 6239
rect 12265 6205 12299 6239
rect 12633 6205 12667 6239
rect 15853 6205 15887 6239
rect 18153 6205 18187 6239
rect 19257 6205 19291 6239
rect 22385 6205 22419 6239
rect 22477 6205 22511 6239
rect 24400 6205 24434 6239
rect 4077 6137 4111 6171
rect 4813 6137 4847 6171
rect 7665 6137 7699 6171
rect 8392 6137 8426 6171
rect 14004 6137 14038 6171
rect 16313 6137 16347 6171
rect 19073 6137 19107 6171
rect 19524 6137 19558 6171
rect 21557 6137 21591 6171
rect 1409 6069 1443 6103
rect 8033 6069 8067 6103
rect 10057 6069 10091 6103
rect 10609 6069 10643 6103
rect 10977 6069 11011 6103
rect 12817 6069 12851 6103
rect 16405 6069 16439 6103
rect 16773 6069 16807 6103
rect 18337 6069 18371 6103
rect 20637 6069 20671 6103
rect 21833 6069 21867 6103
rect 22017 6069 22051 6103
rect 25513 6069 25547 6103
rect 1593 5865 1627 5899
rect 2329 5865 2363 5899
rect 3433 5865 3467 5899
rect 4077 5865 4111 5899
rect 4537 5865 4571 5899
rect 5641 5865 5675 5899
rect 8033 5865 8067 5899
rect 9689 5865 9723 5899
rect 10885 5865 10919 5899
rect 11345 5865 11379 5899
rect 12541 5865 12575 5899
rect 14105 5865 14139 5899
rect 14657 5865 14691 5899
rect 15025 5865 15059 5899
rect 16129 5865 16163 5899
rect 16497 5865 16531 5899
rect 18797 5865 18831 5899
rect 19073 5865 19107 5899
rect 19717 5865 19751 5899
rect 21557 5865 21591 5899
rect 22017 5865 22051 5899
rect 24133 5865 24167 5899
rect 24409 5865 24443 5899
rect 24961 5865 24995 5899
rect 3801 5797 3835 5831
rect 6009 5797 6043 5831
rect 8401 5797 8435 5831
rect 12992 5797 13026 5831
rect 17040 5797 17074 5831
rect 19625 5797 19659 5831
rect 2697 5729 2731 5763
rect 4445 5729 4479 5763
rect 5181 5729 5215 5763
rect 10057 5729 10091 5763
rect 11621 5729 11655 5763
rect 15301 5729 15335 5763
rect 16773 5729 16807 5763
rect 20269 5729 20303 5763
rect 21005 5729 21039 5763
rect 22109 5729 22143 5763
rect 22376 5729 22410 5763
rect 2789 5661 2823 5695
rect 2881 5661 2915 5695
rect 4721 5661 4755 5695
rect 6101 5661 6135 5695
rect 6285 5661 6319 5695
rect 6929 5661 6963 5695
rect 8493 5661 8527 5695
rect 8677 5661 8711 5695
rect 10149 5661 10183 5695
rect 10333 5661 10367 5695
rect 12725 5661 12759 5695
rect 19901 5661 19935 5695
rect 25053 5661 25087 5695
rect 25145 5661 25179 5695
rect 1961 5593 1995 5627
rect 5549 5593 5583 5627
rect 7941 5593 7975 5627
rect 24593 5593 24627 5627
rect 7205 5525 7239 5559
rect 9413 5525 9447 5559
rect 11805 5525 11839 5559
rect 15485 5525 15519 5559
rect 18153 5525 18187 5559
rect 19257 5525 19291 5559
rect 20637 5525 20671 5559
rect 21189 5525 21223 5559
rect 23489 5525 23523 5559
rect 1409 5321 1443 5355
rect 3801 5321 3835 5355
rect 4169 5321 4203 5355
rect 5641 5321 5675 5355
rect 11253 5321 11287 5355
rect 13461 5321 13495 5355
rect 17049 5321 17083 5355
rect 17785 5321 17819 5355
rect 19993 5321 20027 5355
rect 23029 5321 23063 5355
rect 23949 5321 23983 5355
rect 24409 5321 24443 5355
rect 25421 5321 25455 5355
rect 8769 5253 8803 5287
rect 10701 5253 10735 5287
rect 12173 5253 12207 5287
rect 13553 5253 13587 5287
rect 19441 5253 19475 5287
rect 24225 5253 24259 5287
rect 1961 5185 1995 5219
rect 3249 5185 3283 5219
rect 13001 5185 13035 5219
rect 14013 5185 14047 5219
rect 14105 5185 14139 5219
rect 18061 5185 18095 5219
rect 21189 5185 21223 5219
rect 21557 5185 21591 5219
rect 24961 5185 24995 5219
rect 1777 5117 1811 5151
rect 4261 5117 4295 5151
rect 6561 5117 6595 5151
rect 6837 5117 6871 5151
rect 7104 5117 7138 5151
rect 9321 5117 9355 5151
rect 12449 5117 12483 5151
rect 14933 5117 14967 5151
rect 15117 5117 15151 5151
rect 18317 5117 18351 5151
rect 20913 5117 20947 5151
rect 22477 5117 22511 5151
rect 24869 5117 24903 5151
rect 2421 5049 2455 5083
rect 4528 5049 4562 5083
rect 9566 5049 9600 5083
rect 13921 5049 13955 5083
rect 14657 5049 14691 5083
rect 15362 5049 15396 5083
rect 17509 5049 17543 5083
rect 21005 5049 21039 5083
rect 24777 5049 24811 5083
rect 1869 4981 1903 5015
rect 2881 4981 2915 5015
rect 6193 4981 6227 5015
rect 8217 4981 8251 5015
rect 9137 4981 9171 5015
rect 11897 4981 11931 5015
rect 12633 4981 12667 5015
rect 16497 4981 16531 5015
rect 20361 4981 20395 5015
rect 20545 4981 20579 5015
rect 22109 4981 22143 5015
rect 22661 4981 22695 5015
rect 1593 4777 1627 4811
rect 2053 4777 2087 4811
rect 2421 4777 2455 4811
rect 5181 4777 5215 4811
rect 5273 4777 5307 4811
rect 6377 4777 6411 4811
rect 6745 4777 6779 4811
rect 7941 4777 7975 4811
rect 9321 4777 9355 4811
rect 10701 4777 10735 4811
rect 12541 4777 12575 4811
rect 13645 4777 13679 4811
rect 15025 4777 15059 4811
rect 15761 4777 15795 4811
rect 16313 4777 16347 4811
rect 16773 4777 16807 4811
rect 17233 4777 17267 4811
rect 17969 4777 18003 4811
rect 19165 4777 19199 4811
rect 19533 4777 19567 4811
rect 20177 4777 20211 4811
rect 20637 4777 20671 4811
rect 20913 4777 20947 4811
rect 21281 4777 21315 4811
rect 22201 4777 22235 4811
rect 24501 4777 24535 4811
rect 2513 4709 2547 4743
rect 6837 4709 6871 4743
rect 8401 4709 8435 4743
rect 11406 4709 11440 4743
rect 14105 4709 14139 4743
rect 17325 4709 17359 4743
rect 19073 4709 19107 4743
rect 19625 4709 19659 4743
rect 21373 4709 21407 4743
rect 24869 4709 24903 4743
rect 3893 4641 3927 4675
rect 4721 4641 4755 4675
rect 8309 4641 8343 4675
rect 10057 4641 10091 4675
rect 11161 4641 11195 4675
rect 14013 4641 14047 4675
rect 15669 4641 15703 4675
rect 22477 4641 22511 4675
rect 22744 4641 22778 4675
rect 24961 4641 24995 4675
rect 2697 4573 2731 4607
rect 3433 4573 3467 4607
rect 5365 4573 5399 4607
rect 6929 4573 6963 4607
rect 8493 4573 8527 4607
rect 14197 4573 14231 4607
rect 15853 4573 15887 4607
rect 17509 4573 17543 4607
rect 19717 4573 19751 4607
rect 21557 4573 21591 4607
rect 4813 4505 4847 4539
rect 6285 4505 6319 4539
rect 7481 4505 7515 4539
rect 7849 4505 7883 4539
rect 10241 4505 10275 4539
rect 16865 4505 16899 4539
rect 3065 4437 3099 4471
rect 4261 4437 4295 4471
rect 5825 4437 5859 4471
rect 9045 4437 9079 4471
rect 9965 4437 9999 4471
rect 11069 4437 11103 4471
rect 13185 4437 13219 4471
rect 13553 4437 13587 4471
rect 14749 4437 14783 4471
rect 15301 4437 15335 4471
rect 18337 4437 18371 4471
rect 18705 4437 18739 4471
rect 23857 4437 23891 4471
rect 25145 4437 25179 4471
rect 5181 4233 5215 4267
rect 9965 4233 9999 4267
rect 13093 4233 13127 4267
rect 14105 4233 14139 4267
rect 16221 4233 16255 4267
rect 17325 4233 17359 4267
rect 19349 4233 19383 4267
rect 21741 4233 21775 4267
rect 23397 4233 23431 4267
rect 25881 4233 25915 4267
rect 4537 4165 4571 4199
rect 4905 4165 4939 4199
rect 11161 4165 11195 4199
rect 11529 4165 11563 4199
rect 1961 4097 1995 4131
rect 2053 4097 2087 4131
rect 5733 4097 5767 4131
rect 7389 4097 7423 4131
rect 8861 4097 8895 4131
rect 9045 4097 9079 4131
rect 9873 4097 9907 4131
rect 10517 4097 10551 4131
rect 13553 4097 13587 4131
rect 13645 4097 13679 4131
rect 14565 4097 14599 4131
rect 15209 4097 15243 4131
rect 16773 4097 16807 4131
rect 17877 4097 17911 4131
rect 18705 4097 18739 4131
rect 18889 4097 18923 4131
rect 19901 4097 19935 4131
rect 21281 4097 21315 4131
rect 23029 4097 23063 4131
rect 24777 4097 24811 4131
rect 5641 4029 5675 4063
rect 7297 4029 7331 4063
rect 9413 4029 9447 4063
rect 10425 4029 10459 4063
rect 12173 4029 12207 4063
rect 13001 4029 13035 4063
rect 15117 4029 15151 4063
rect 15945 4029 15979 4063
rect 16589 4029 16623 4063
rect 18613 4029 18647 4063
rect 21097 4029 21131 4063
rect 22477 4029 22511 4063
rect 24501 4029 24535 4063
rect 2320 3961 2354 3995
rect 5549 3961 5583 3995
rect 8769 3961 8803 3995
rect 13461 3961 13495 3995
rect 15025 3961 15059 3995
rect 16037 3961 16071 3995
rect 16681 3961 16715 3995
rect 20269 3961 20303 3995
rect 22201 3961 22235 3995
rect 24593 3961 24627 3995
rect 25513 3961 25547 3995
rect 3433 3893 3467 3927
rect 4077 3893 4111 3927
rect 6193 3893 6227 3927
rect 6561 3893 6595 3927
rect 6837 3893 6871 3927
rect 7205 3893 7239 3927
rect 8033 3893 8067 3927
rect 8401 3893 8435 3927
rect 10333 3893 10367 3927
rect 14657 3893 14691 3927
rect 15669 3893 15703 3927
rect 15945 3893 15979 3927
rect 18245 3893 18279 3927
rect 20545 3893 20579 3927
rect 20729 3893 20763 3927
rect 21189 3893 21223 3927
rect 22661 3893 22695 3927
rect 23949 3893 23983 3927
rect 24133 3893 24167 3927
rect 25145 3893 25179 3927
rect 2513 3689 2547 3723
rect 3157 3689 3191 3723
rect 3433 3689 3467 3723
rect 5457 3689 5491 3723
rect 6561 3689 6595 3723
rect 8033 3689 8067 3723
rect 9505 3689 9539 3723
rect 10701 3689 10735 3723
rect 12173 3689 12207 3723
rect 12725 3689 12759 3723
rect 13277 3689 13311 3723
rect 14289 3689 14323 3723
rect 15025 3689 15059 3723
rect 15301 3689 15335 3723
rect 15761 3689 15795 3723
rect 16681 3689 16715 3723
rect 17049 3689 17083 3723
rect 17417 3689 17451 3723
rect 18061 3689 18095 3723
rect 18521 3689 18555 3723
rect 19073 3689 19107 3723
rect 19533 3689 19567 3723
rect 21373 3689 21407 3723
rect 21925 3689 21959 3723
rect 22293 3689 22327 3723
rect 23029 3689 23063 3723
rect 2421 3621 2455 3655
rect 4322 3621 4356 3655
rect 10241 3621 10275 3655
rect 11060 3621 11094 3655
rect 18429 3621 18463 3655
rect 21281 3621 21315 3655
rect 23848 3621 23882 3655
rect 6929 3553 6963 3587
rect 9689 3553 9723 3587
rect 10793 3553 10827 3587
rect 13185 3553 13219 3587
rect 13645 3553 13679 3587
rect 15669 3553 15703 3587
rect 16405 3553 16439 3587
rect 16865 3553 16899 3587
rect 19717 3553 19751 3587
rect 20269 3553 20303 3587
rect 20729 3553 20763 3587
rect 22477 3553 22511 3587
rect 23581 3553 23615 3587
rect 2697 3485 2731 3519
rect 4077 3485 4111 3519
rect 7021 3485 7055 3519
rect 7113 3485 7147 3519
rect 7665 3485 7699 3519
rect 8585 3485 8619 3519
rect 13737 3485 13771 3519
rect 13829 3485 13863 3519
rect 15853 3485 15887 3519
rect 18613 3485 18647 3519
rect 21465 3485 21499 3519
rect 2053 3417 2087 3451
rect 17969 3417 18003 3451
rect 20913 3417 20947 3451
rect 1685 3349 1719 3383
rect 3893 3349 3927 3383
rect 6009 3349 6043 3383
rect 6377 3349 6411 3383
rect 8401 3349 8435 3383
rect 9137 3349 9171 3383
rect 9873 3349 9907 3383
rect 14657 3349 14691 3383
rect 19901 3349 19935 3383
rect 22661 3349 22695 3383
rect 23489 3349 23523 3383
rect 24961 3349 24995 3383
rect 2973 3145 3007 3179
rect 6193 3145 6227 3179
rect 6837 3145 6871 3179
rect 7941 3145 7975 3179
rect 8585 3145 8619 3179
rect 10149 3145 10183 3179
rect 10885 3145 10919 3179
rect 11805 3145 11839 3179
rect 14197 3145 14231 3179
rect 16129 3145 16163 3179
rect 17049 3145 17083 3179
rect 17509 3145 17543 3179
rect 17785 3145 17819 3179
rect 19441 3145 19475 3179
rect 20085 3145 20119 3179
rect 22477 3145 22511 3179
rect 23489 3145 23523 3179
rect 23949 3145 23983 3179
rect 25513 3145 25547 3179
rect 26065 3145 26099 3179
rect 12173 3077 12207 3111
rect 12449 3077 12483 3111
rect 13921 3077 13955 3111
rect 16681 3077 16715 3111
rect 21925 3077 21959 3111
rect 23121 3077 23155 3111
rect 1593 3009 1627 3043
rect 7389 3009 7423 3043
rect 8309 3009 8343 3043
rect 13001 3009 13035 3043
rect 18061 3009 18095 3043
rect 24133 3009 24167 3043
rect 1860 2941 1894 2975
rect 4261 2941 4295 2975
rect 4517 2941 4551 2975
rect 7297 2941 7331 2975
rect 8769 2941 8803 2975
rect 9036 2941 9070 2975
rect 11253 2941 11287 2975
rect 12909 2941 12943 2975
rect 14749 2941 14783 2975
rect 18317 2941 18351 2975
rect 20545 2941 20579 2975
rect 24400 2941 24434 2975
rect 3709 2873 3743 2907
rect 4077 2873 4111 2907
rect 6561 2873 6595 2907
rect 12817 2873 12851 2907
rect 14994 2873 15028 2907
rect 20790 2873 20824 2907
rect 5641 2805 5675 2839
rect 7205 2805 7239 2839
rect 11437 2805 11471 2839
rect 13461 2805 13495 2839
rect 14565 2805 14599 2839
rect 20453 2805 20487 2839
rect 1685 2601 1719 2635
rect 1869 2601 1903 2635
rect 2881 2601 2915 2635
rect 3893 2601 3927 2635
rect 5733 2601 5767 2635
rect 6745 2601 6779 2635
rect 9137 2601 9171 2635
rect 9781 2601 9815 2635
rect 10149 2601 10183 2635
rect 10885 2601 10919 2635
rect 14013 2601 14047 2635
rect 16865 2601 16899 2635
rect 18061 2601 18095 2635
rect 19717 2601 19751 2635
rect 20637 2601 20671 2635
rect 20913 2601 20947 2635
rect 22569 2601 22603 2635
rect 23765 2601 23799 2635
rect 24225 2601 24259 2635
rect 2329 2533 2363 2567
rect 2237 2465 2271 2499
rect 4353 2465 4387 2499
rect 4620 2465 4654 2499
rect 6653 2465 6687 2499
rect 2513 2397 2547 2431
rect 3525 2397 3559 2431
rect 7472 2533 7506 2567
rect 10241 2533 10275 2567
rect 12081 2533 12115 2567
rect 12878 2533 12912 2567
rect 18604 2533 18638 2567
rect 21456 2533 21490 2567
rect 24593 2533 24627 2567
rect 7205 2465 7239 2499
rect 11253 2465 11287 2499
rect 11437 2465 11471 2499
rect 15209 2465 15243 2499
rect 15485 2465 15519 2499
rect 15741 2465 15775 2499
rect 17693 2465 17727 2499
rect 18337 2465 18371 2499
rect 21189 2465 21223 2499
rect 10333 2397 10367 2431
rect 12357 2397 12391 2431
rect 12633 2397 12667 2431
rect 14933 2397 14967 2431
rect 23489 2397 23523 2431
rect 24685 2397 24719 2431
rect 24777 2397 24811 2431
rect 25237 2397 25271 2431
rect 8585 2329 8619 2363
rect 6745 2261 6779 2295
rect 9505 2261 9539 2295
rect 11621 2261 11655 2295
<< metal1 >>
rect 17218 26800 17224 26852
rect 17276 26840 17282 26852
rect 23474 26840 23480 26852
rect 17276 26812 23480 26840
rect 17276 26800 17282 26812
rect 23474 26800 23480 26812
rect 23532 26800 23538 26852
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 24762 23304 24768 23316
rect 24723 23276 24768 23304
rect 24762 23264 24768 23276
rect 24820 23264 24826 23316
rect 24581 23171 24639 23177
rect 24581 23137 24593 23171
rect 24627 23168 24639 23171
rect 24670 23168 24676 23180
rect 24627 23140 24676 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1578 22760 1584 22772
rect 1539 22732 1584 22760
rect 1578 22720 1584 22732
rect 1636 22720 1642 22772
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22556 1455 22559
rect 1762 22556 1768 22568
rect 1443 22528 1768 22556
rect 1443 22525 1455 22528
rect 1397 22519 1455 22525
rect 1762 22516 1768 22528
rect 1820 22556 1826 22568
rect 1949 22559 2007 22565
rect 1949 22556 1961 22559
rect 1820 22528 1961 22556
rect 1820 22516 1826 22528
rect 1949 22525 1961 22528
rect 1995 22525 2007 22559
rect 1949 22519 2007 22525
rect 24578 22420 24584 22432
rect 24539 22392 24584 22420
rect 24578 22380 24584 22392
rect 24636 22380 24642 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 23753 22219 23811 22225
rect 23753 22185 23765 22219
rect 23799 22216 23811 22219
rect 24578 22216 24584 22228
rect 23799 22188 24584 22216
rect 23799 22185 23811 22188
rect 23753 22179 23811 22185
rect 24578 22176 24584 22188
rect 24636 22176 24642 22228
rect 23569 22083 23627 22089
rect 23569 22049 23581 22083
rect 23615 22080 23627 22083
rect 23842 22080 23848 22092
rect 23615 22052 23848 22080
rect 23615 22049 23627 22052
rect 23569 22043 23627 22049
rect 23842 22040 23848 22052
rect 23900 22040 23906 22092
rect 24118 22040 24124 22092
rect 24176 22080 24182 22092
rect 24581 22083 24639 22089
rect 24581 22080 24593 22083
rect 24176 22052 24593 22080
rect 24176 22040 24182 22052
rect 24581 22049 24593 22052
rect 24627 22049 24639 22083
rect 24581 22043 24639 22049
rect 24762 21944 24768 21956
rect 24723 21916 24768 21944
rect 24762 21904 24768 21916
rect 24820 21904 24826 21956
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 24670 21632 24676 21684
rect 24728 21672 24734 21684
rect 24765 21675 24823 21681
rect 24765 21672 24777 21675
rect 24728 21644 24777 21672
rect 24728 21632 24734 21644
rect 24765 21641 24777 21644
rect 24811 21641 24823 21675
rect 24765 21635 24823 21641
rect 23842 21468 23848 21480
rect 23803 21440 23848 21468
rect 23842 21428 23848 21440
rect 23900 21428 23906 21480
rect 23934 21428 23940 21480
rect 23992 21468 23998 21480
rect 24581 21471 24639 21477
rect 24581 21468 24593 21471
rect 23992 21440 24593 21468
rect 23992 21428 23998 21440
rect 24581 21437 24593 21440
rect 24627 21468 24639 21471
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24627 21440 25145 21468
rect 24627 21437 24639 21440
rect 24581 21431 24639 21437
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 24118 21292 24124 21344
rect 24176 21332 24182 21344
rect 24397 21335 24455 21341
rect 24397 21332 24409 21335
rect 24176 21304 24409 21332
rect 24176 21292 24182 21304
rect 24397 21301 24409 21304
rect 24443 21301 24455 21335
rect 24397 21295 24455 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1762 21128 1768 21140
rect 1723 21100 1768 21128
rect 1762 21088 1768 21100
rect 1820 21088 1826 21140
rect 1581 20995 1639 21001
rect 1581 20961 1593 20995
rect 1627 20992 1639 20995
rect 2498 20992 2504 21004
rect 1627 20964 2504 20992
rect 1627 20961 1639 20964
rect 1581 20955 1639 20961
rect 2498 20952 2504 20964
rect 2556 20952 2562 21004
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1578 20584 1584 20596
rect 1539 20556 1584 20584
rect 1578 20544 1584 20556
rect 1636 20544 1642 20596
rect 13262 20408 13268 20460
rect 13320 20448 13326 20460
rect 13357 20451 13415 20457
rect 13357 20448 13369 20451
rect 13320 20420 13369 20448
rect 13320 20408 13326 20420
rect 13357 20417 13369 20420
rect 13403 20417 13415 20451
rect 13357 20411 13415 20417
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 1443 20352 1808 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 1780 20256 1808 20352
rect 13265 20315 13323 20321
rect 13265 20281 13277 20315
rect 13311 20312 13323 20315
rect 13624 20315 13682 20321
rect 13624 20312 13636 20315
rect 13311 20284 13636 20312
rect 13311 20281 13323 20284
rect 13265 20275 13323 20281
rect 13624 20281 13636 20284
rect 13670 20312 13682 20315
rect 13722 20312 13728 20324
rect 13670 20284 13728 20312
rect 13670 20281 13682 20284
rect 13624 20275 13682 20281
rect 13722 20272 13728 20284
rect 13780 20272 13786 20324
rect 1762 20204 1768 20256
rect 1820 20244 1826 20256
rect 1949 20247 2007 20253
rect 1949 20244 1961 20247
rect 1820 20216 1961 20244
rect 1820 20204 1826 20216
rect 1949 20213 1961 20216
rect 1995 20213 2007 20247
rect 1949 20207 2007 20213
rect 2409 20247 2467 20253
rect 2409 20213 2421 20247
rect 2455 20244 2467 20247
rect 2498 20244 2504 20256
rect 2455 20216 2504 20244
rect 2455 20213 2467 20216
rect 2409 20207 2467 20213
rect 2498 20204 2504 20216
rect 2556 20204 2562 20256
rect 14734 20244 14740 20256
rect 14695 20216 14740 20244
rect 14734 20204 14740 20216
rect 14792 20204 14798 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1486 20000 1492 20052
rect 1544 20040 1550 20052
rect 1581 20043 1639 20049
rect 1581 20040 1593 20043
rect 1544 20012 1593 20040
rect 1544 20000 1550 20012
rect 1581 20009 1593 20012
rect 1627 20009 1639 20043
rect 1581 20003 1639 20009
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 2130 19904 2136 19916
rect 1443 19876 2136 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 2130 19864 2136 19876
rect 2188 19864 2194 19916
rect 13262 19660 13268 19712
rect 13320 19700 13326 19712
rect 13357 19703 13415 19709
rect 13357 19700 13369 19703
rect 13320 19672 13369 19700
rect 13320 19660 13326 19672
rect 13357 19669 13369 19672
rect 13403 19669 13415 19703
rect 13357 19663 13415 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19261 1455 19295
rect 13541 19295 13599 19301
rect 13541 19292 13553 19295
rect 1397 19255 1455 19261
rect 13372 19264 13553 19292
rect 1412 19224 1440 19255
rect 2406 19224 2412 19236
rect 1412 19196 2412 19224
rect 2406 19184 2412 19196
rect 2464 19184 2470 19236
rect 1394 19116 1400 19168
rect 1452 19156 1458 19168
rect 1581 19159 1639 19165
rect 1581 19156 1593 19159
rect 1452 19128 1593 19156
rect 1452 19116 1458 19128
rect 1581 19125 1593 19128
rect 1627 19125 1639 19159
rect 1581 19119 1639 19125
rect 2041 19159 2099 19165
rect 2041 19125 2053 19159
rect 2087 19156 2099 19159
rect 2130 19156 2136 19168
rect 2087 19128 2136 19156
rect 2087 19125 2099 19128
rect 2041 19119 2099 19125
rect 2130 19116 2136 19128
rect 2188 19116 2194 19168
rect 13262 19116 13268 19168
rect 13320 19156 13326 19168
rect 13372 19165 13400 19264
rect 13541 19261 13553 19264
rect 13587 19261 13599 19295
rect 13541 19255 13599 19261
rect 13808 19227 13866 19233
rect 13808 19193 13820 19227
rect 13854 19224 13866 19227
rect 14090 19224 14096 19236
rect 13854 19196 14096 19224
rect 13854 19193 13866 19196
rect 13808 19187 13866 19193
rect 14090 19184 14096 19196
rect 14148 19184 14154 19236
rect 13357 19159 13415 19165
rect 13357 19156 13369 19159
rect 13320 19128 13369 19156
rect 13320 19116 13326 19128
rect 13357 19125 13369 19128
rect 13403 19125 13415 19159
rect 14918 19156 14924 19168
rect 14879 19128 14924 19156
rect 13357 19119 13415 19125
rect 14918 19116 14924 19128
rect 14976 19116 14982 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1762 18952 1768 18964
rect 1723 18924 1768 18952
rect 1762 18912 1768 18924
rect 1820 18912 1826 18964
rect 1581 18819 1639 18825
rect 1581 18785 1593 18819
rect 1627 18816 1639 18819
rect 2406 18816 2412 18828
rect 1627 18788 2412 18816
rect 1627 18785 1639 18788
rect 1581 18779 1639 18785
rect 2406 18776 2412 18788
rect 2464 18776 2470 18828
rect 12802 18816 12808 18828
rect 12763 18788 12808 18816
rect 12802 18776 12808 18788
rect 12860 18776 12866 18828
rect 14918 18816 14924 18828
rect 13096 18788 14924 18816
rect 13096 18760 13124 18788
rect 14918 18776 14924 18788
rect 14976 18776 14982 18828
rect 12897 18751 12955 18757
rect 12897 18717 12909 18751
rect 12943 18717 12955 18751
rect 13078 18748 13084 18760
rect 12991 18720 13084 18748
rect 12897 18711 12955 18717
rect 12434 18640 12440 18692
rect 12492 18680 12498 18692
rect 12492 18652 12537 18680
rect 12492 18640 12498 18652
rect 12342 18612 12348 18624
rect 12255 18584 12348 18612
rect 12342 18572 12348 18584
rect 12400 18612 12406 18624
rect 12912 18612 12940 18711
rect 13078 18708 13084 18720
rect 13136 18708 13142 18760
rect 13998 18748 14004 18760
rect 13959 18720 14004 18748
rect 13998 18708 14004 18720
rect 14056 18708 14062 18760
rect 12400 18584 12940 18612
rect 13633 18615 13691 18621
rect 12400 18572 12406 18584
rect 13633 18581 13645 18615
rect 13679 18612 13691 18615
rect 14090 18612 14096 18624
rect 13679 18584 14096 18612
rect 13679 18581 13691 18584
rect 13633 18575 13691 18581
rect 14090 18572 14096 18584
rect 14148 18572 14154 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1578 18408 1584 18420
rect 1539 18380 1584 18408
rect 1578 18368 1584 18380
rect 1636 18368 1642 18420
rect 2406 18408 2412 18420
rect 2367 18380 2412 18408
rect 2406 18368 2412 18380
rect 2464 18368 2470 18420
rect 11517 18411 11575 18417
rect 11517 18377 11529 18411
rect 11563 18408 11575 18411
rect 12802 18408 12808 18420
rect 11563 18380 12808 18408
rect 11563 18377 11575 18380
rect 11517 18371 11575 18377
rect 12802 18368 12808 18380
rect 12860 18368 12866 18420
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 1443 18176 2084 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 2056 18080 2084 18176
rect 11808 18176 12449 18204
rect 2038 18068 2044 18080
rect 1999 18040 2044 18068
rect 2038 18028 2044 18040
rect 2096 18028 2102 18080
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11808 18077 11836 18176
rect 12437 18173 12449 18176
rect 12483 18204 12495 18207
rect 13262 18204 13268 18216
rect 12483 18176 13268 18204
rect 12483 18173 12495 18176
rect 12437 18167 12495 18173
rect 13262 18164 13268 18176
rect 13320 18164 13326 18216
rect 12710 18145 12716 18148
rect 12704 18136 12716 18145
rect 12671 18108 12716 18136
rect 12704 18099 12716 18108
rect 12710 18096 12716 18099
rect 12768 18096 12774 18148
rect 11793 18071 11851 18077
rect 11793 18068 11805 18071
rect 11112 18040 11805 18068
rect 11112 18028 11118 18040
rect 11793 18037 11805 18040
rect 11839 18037 11851 18071
rect 11793 18031 11851 18037
rect 12253 18071 12311 18077
rect 12253 18037 12265 18071
rect 12299 18068 12311 18071
rect 13078 18068 13084 18080
rect 12299 18040 13084 18068
rect 12299 18037 12311 18040
rect 12253 18031 12311 18037
rect 13078 18028 13084 18040
rect 13136 18028 13142 18080
rect 13817 18071 13875 18077
rect 13817 18037 13829 18071
rect 13863 18068 13875 18071
rect 14090 18068 14096 18080
rect 13863 18040 14096 18068
rect 13863 18037 13875 18040
rect 13817 18031 13875 18037
rect 14090 18028 14096 18040
rect 14148 18028 14154 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1581 17867 1639 17873
rect 1581 17833 1593 17867
rect 1627 17864 1639 17867
rect 1670 17864 1676 17876
rect 1627 17836 1676 17864
rect 1627 17833 1639 17836
rect 1581 17827 1639 17833
rect 1670 17824 1676 17836
rect 1728 17824 1734 17876
rect 12802 17824 12808 17876
rect 12860 17864 12866 17876
rect 13541 17867 13599 17873
rect 13541 17864 13553 17867
rect 12860 17836 13553 17864
rect 12860 17824 12866 17836
rect 13541 17833 13553 17836
rect 13587 17833 13599 17867
rect 13541 17827 13599 17833
rect 13909 17867 13967 17873
rect 13909 17833 13921 17867
rect 13955 17864 13967 17867
rect 13998 17864 14004 17876
rect 13955 17836 14004 17864
rect 13955 17833 13967 17836
rect 13909 17827 13967 17833
rect 13998 17824 14004 17836
rect 14056 17824 14062 17876
rect 14645 17867 14703 17873
rect 14645 17833 14657 17867
rect 14691 17864 14703 17867
rect 14734 17864 14740 17876
rect 14691 17836 14740 17864
rect 14691 17833 14703 17836
rect 14645 17827 14703 17833
rect 14734 17824 14740 17836
rect 14792 17824 14798 17876
rect 24762 17864 24768 17876
rect 24723 17836 24768 17864
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 2314 17728 2320 17740
rect 1443 17700 2320 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 2314 17688 2320 17700
rect 2372 17688 2378 17740
rect 10778 17688 10784 17740
rect 10836 17728 10842 17740
rect 11313 17731 11371 17737
rect 11313 17728 11325 17731
rect 10836 17700 11325 17728
rect 10836 17688 10842 17700
rect 11313 17697 11325 17700
rect 11359 17697 11371 17731
rect 11313 17691 11371 17697
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 24670 17728 24676 17740
rect 24627 17700 24676 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 24670 17688 24676 17700
rect 24728 17688 24734 17740
rect 11054 17660 11060 17672
rect 11015 17632 11060 17660
rect 11054 17620 11060 17632
rect 11112 17620 11118 17672
rect 13538 17620 13544 17672
rect 13596 17660 13602 17672
rect 14001 17663 14059 17669
rect 14001 17660 14013 17663
rect 13596 17632 14013 17660
rect 13596 17620 13602 17632
rect 14001 17629 14013 17632
rect 14047 17629 14059 17663
rect 14001 17623 14059 17629
rect 14090 17620 14096 17672
rect 14148 17660 14154 17672
rect 15289 17663 15347 17669
rect 14148 17632 14193 17660
rect 14148 17620 14154 17632
rect 15289 17629 15301 17663
rect 15335 17660 15347 17663
rect 15654 17660 15660 17672
rect 15335 17632 15660 17660
rect 15335 17629 15347 17632
rect 15289 17623 15347 17629
rect 15654 17620 15660 17632
rect 15712 17620 15718 17672
rect 12437 17595 12495 17601
rect 12437 17561 12449 17595
rect 12483 17592 12495 17595
rect 12710 17592 12716 17604
rect 12483 17564 12716 17592
rect 12483 17561 12495 17564
rect 12437 17555 12495 17561
rect 12710 17552 12716 17564
rect 12768 17592 12774 17604
rect 13081 17595 13139 17601
rect 13081 17592 13093 17595
rect 12768 17564 13093 17592
rect 12768 17552 12774 17564
rect 13081 17561 13093 17564
rect 13127 17592 13139 17595
rect 13630 17592 13636 17604
rect 13127 17564 13636 17592
rect 13127 17561 13139 17564
rect 13081 17555 13139 17561
rect 13630 17552 13636 17564
rect 13688 17552 13694 17604
rect 10781 17527 10839 17533
rect 10781 17493 10793 17527
rect 10827 17524 10839 17527
rect 11330 17524 11336 17536
rect 10827 17496 11336 17524
rect 10827 17493 10839 17496
rect 10781 17487 10839 17493
rect 11330 17484 11336 17496
rect 11388 17484 11394 17536
rect 13354 17524 13360 17536
rect 13315 17496 13360 17524
rect 13354 17484 13360 17496
rect 13412 17484 13418 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1486 17280 1492 17332
rect 1544 17320 1550 17332
rect 1581 17323 1639 17329
rect 1581 17320 1593 17323
rect 1544 17292 1593 17320
rect 1544 17280 1550 17292
rect 1581 17289 1593 17292
rect 1627 17289 1639 17323
rect 2314 17320 2320 17332
rect 2275 17292 2320 17320
rect 1581 17283 1639 17289
rect 2314 17280 2320 17292
rect 2372 17280 2378 17332
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 12492 17292 12537 17320
rect 12492 17280 12498 17292
rect 24210 17280 24216 17332
rect 24268 17320 24274 17332
rect 24765 17323 24823 17329
rect 24765 17320 24777 17323
rect 24268 17292 24777 17320
rect 24268 17280 24274 17292
rect 24765 17289 24777 17292
rect 24811 17289 24823 17323
rect 24765 17283 24823 17289
rect 14185 17255 14243 17261
rect 14185 17252 14197 17255
rect 12176 17224 14197 17252
rect 10134 17144 10140 17196
rect 10192 17184 10198 17196
rect 11149 17187 11207 17193
rect 11149 17184 11161 17187
rect 10192 17156 11161 17184
rect 10192 17144 10198 17156
rect 11149 17153 11161 17156
rect 11195 17153 11207 17187
rect 11330 17184 11336 17196
rect 11243 17156 11336 17184
rect 11149 17147 11207 17153
rect 11330 17144 11336 17156
rect 11388 17184 11394 17196
rect 11790 17184 11796 17196
rect 11388 17156 11796 17184
rect 11388 17144 11394 17156
rect 11790 17144 11796 17156
rect 11848 17144 11854 17196
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 10597 17119 10655 17125
rect 1443 17088 2084 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 2056 16989 2084 17088
rect 10597 17085 10609 17119
rect 10643 17116 10655 17119
rect 10778 17116 10784 17128
rect 10643 17088 10784 17116
rect 10643 17085 10655 17088
rect 10597 17079 10655 17085
rect 10778 17076 10784 17088
rect 10836 17076 10842 17128
rect 9861 17051 9919 17057
rect 9861 17017 9873 17051
rect 9907 17048 9919 17051
rect 9907 17020 11100 17048
rect 9907 17017 9919 17020
rect 9861 17011 9919 17017
rect 11072 16992 11100 17020
rect 2041 16983 2099 16989
rect 2041 16949 2053 16983
rect 2087 16980 2099 16983
rect 3326 16980 3332 16992
rect 2087 16952 3332 16980
rect 2087 16949 2099 16952
rect 2041 16943 2099 16949
rect 3326 16940 3332 16952
rect 3384 16940 3390 16992
rect 10134 16980 10140 16992
rect 10095 16952 10140 16980
rect 10134 16940 10140 16952
rect 10192 16940 10198 16992
rect 10686 16980 10692 16992
rect 10647 16952 10692 16980
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 11054 16980 11060 16992
rect 11015 16952 11060 16980
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 11238 16940 11244 16992
rect 11296 16980 11302 16992
rect 11701 16983 11759 16989
rect 11701 16980 11713 16983
rect 11296 16952 11713 16980
rect 11296 16940 11302 16952
rect 11701 16949 11713 16952
rect 11747 16980 11759 16983
rect 12176 16980 12204 17224
rect 14185 17221 14197 17224
rect 14231 17252 14243 17255
rect 14231 17224 14412 17252
rect 14231 17221 14243 17224
rect 14185 17215 14243 17221
rect 14384 17196 14412 17224
rect 12526 17144 12532 17196
rect 12584 17184 12590 17196
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 12584 17156 13001 17184
rect 12584 17144 12590 17156
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 14366 17184 14372 17196
rect 14279 17156 14372 17184
rect 12989 17147 13047 17153
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 12897 17119 12955 17125
rect 12897 17085 12909 17119
rect 12943 17116 12955 17119
rect 13354 17116 13360 17128
rect 12943 17088 13360 17116
rect 12943 17085 12955 17088
rect 12897 17079 12955 17085
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 23658 17076 23664 17128
rect 23716 17116 23722 17128
rect 24581 17119 24639 17125
rect 24581 17116 24593 17119
rect 23716 17088 24593 17116
rect 23716 17076 23722 17088
rect 24581 17085 24593 17088
rect 24627 17116 24639 17119
rect 25133 17119 25191 17125
rect 25133 17116 25145 17119
rect 24627 17088 25145 17116
rect 24627 17085 24639 17088
rect 24581 17079 24639 17085
rect 25133 17085 25145 17088
rect 25179 17085 25191 17119
rect 25133 17079 25191 17085
rect 13906 17008 13912 17060
rect 13964 17048 13970 17060
rect 14636 17051 14694 17057
rect 14636 17048 14648 17051
rect 13964 17020 14648 17048
rect 13964 17008 13970 17020
rect 14636 17017 14648 17020
rect 14682 17048 14694 17051
rect 14734 17048 14740 17060
rect 14682 17020 14740 17048
rect 14682 17017 14694 17020
rect 14636 17011 14694 17017
rect 14734 17008 14740 17020
rect 14792 17008 14798 17060
rect 11747 16952 12204 16980
rect 11747 16949 11759 16952
rect 11701 16943 11759 16949
rect 12250 16940 12256 16992
rect 12308 16980 12314 16992
rect 12805 16983 12863 16989
rect 12805 16980 12817 16983
rect 12308 16952 12817 16980
rect 12308 16940 12314 16952
rect 12805 16949 12817 16952
rect 12851 16949 12863 16983
rect 13538 16980 13544 16992
rect 13499 16952 13544 16980
rect 12805 16943 12863 16949
rect 13538 16940 13544 16952
rect 13596 16940 13602 16992
rect 15378 16940 15384 16992
rect 15436 16980 15442 16992
rect 15749 16983 15807 16989
rect 15749 16980 15761 16983
rect 15436 16952 15761 16980
rect 15436 16940 15442 16952
rect 15749 16949 15761 16952
rect 15795 16949 15807 16983
rect 24394 16980 24400 16992
rect 24355 16952 24400 16980
rect 15749 16943 15807 16949
rect 24394 16940 24400 16952
rect 24452 16940 24458 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1578 16776 1584 16788
rect 1539 16748 1584 16776
rect 1578 16736 1584 16748
rect 1636 16736 1642 16788
rect 10778 16736 10784 16788
rect 10836 16776 10842 16788
rect 11885 16779 11943 16785
rect 11885 16776 11897 16779
rect 10836 16748 11897 16776
rect 10836 16736 10842 16748
rect 11885 16745 11897 16748
rect 11931 16745 11943 16779
rect 12526 16776 12532 16788
rect 12487 16748 12532 16776
rect 11885 16739 11943 16745
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 12989 16779 13047 16785
rect 12989 16745 13001 16779
rect 13035 16776 13047 16779
rect 13354 16776 13360 16788
rect 13035 16748 13360 16776
rect 13035 16745 13047 16748
rect 12989 16739 13047 16745
rect 13354 16736 13360 16748
rect 13412 16736 13418 16788
rect 13998 16776 14004 16788
rect 13959 16748 14004 16776
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 14734 16736 14740 16788
rect 14792 16776 14798 16788
rect 15013 16779 15071 16785
rect 15013 16776 15025 16779
rect 14792 16748 15025 16776
rect 14792 16736 14798 16748
rect 15013 16745 15025 16748
rect 15059 16745 15071 16779
rect 17034 16776 17040 16788
rect 16995 16748 17040 16776
rect 15013 16739 15071 16745
rect 12544 16708 12572 16736
rect 14090 16708 14096 16720
rect 12544 16680 14096 16708
rect 14090 16668 14096 16680
rect 14148 16708 14154 16720
rect 14369 16711 14427 16717
rect 14369 16708 14381 16711
rect 14148 16680 14381 16708
rect 14148 16668 14154 16680
rect 14369 16677 14381 16680
rect 14415 16677 14427 16711
rect 15028 16708 15056 16739
rect 17034 16736 17040 16748
rect 17092 16736 17098 16788
rect 23753 16779 23811 16785
rect 23753 16745 23765 16779
rect 23799 16776 23811 16779
rect 24394 16776 24400 16788
rect 23799 16748 24400 16776
rect 23799 16745 23811 16748
rect 23753 16739 23811 16745
rect 24394 16736 24400 16748
rect 24452 16736 24458 16788
rect 24762 16776 24768 16788
rect 24723 16748 24768 16776
rect 24762 16736 24768 16748
rect 24820 16736 24826 16788
rect 15028 16680 15884 16708
rect 14369 16671 14427 16677
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 2406 16640 2412 16652
rect 1443 16612 2412 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 2406 16600 2412 16612
rect 2464 16600 2470 16652
rect 9766 16600 9772 16652
rect 9824 16640 9830 16652
rect 10761 16643 10819 16649
rect 10761 16640 10773 16643
rect 9824 16612 10773 16640
rect 9824 16600 9830 16612
rect 10761 16609 10773 16612
rect 10807 16609 10819 16643
rect 13357 16643 13415 16649
rect 13357 16640 13369 16643
rect 10761 16603 10819 16609
rect 12360 16612 13369 16640
rect 10505 16575 10563 16581
rect 10505 16541 10517 16575
rect 10551 16541 10563 16575
rect 10505 16535 10563 16541
rect 8757 16439 8815 16445
rect 8757 16405 8769 16439
rect 8803 16436 8815 16439
rect 9214 16436 9220 16448
rect 8803 16408 9220 16436
rect 8803 16405 8815 16408
rect 8757 16399 8815 16405
rect 9214 16396 9220 16408
rect 9272 16396 9278 16448
rect 10318 16436 10324 16448
rect 10279 16408 10324 16436
rect 10318 16396 10324 16408
rect 10376 16396 10382 16448
rect 10520 16436 10548 16535
rect 12158 16532 12164 16584
rect 12216 16572 12222 16584
rect 12360 16572 12388 16612
rect 13357 16609 13369 16612
rect 13403 16640 13415 16643
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 13403 16612 13768 16640
rect 13403 16609 13415 16612
rect 13357 16603 13415 16609
rect 12216 16544 12388 16572
rect 12216 16532 12222 16544
rect 13262 16532 13268 16584
rect 13320 16572 13326 16584
rect 13449 16575 13507 16581
rect 13449 16572 13461 16575
rect 13320 16544 13461 16572
rect 13320 16532 13326 16544
rect 13449 16541 13461 16544
rect 13495 16541 13507 16575
rect 13630 16572 13636 16584
rect 13591 16544 13636 16572
rect 13449 16535 13507 16541
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 13740 16572 13768 16612
rect 15120 16612 15669 16640
rect 14734 16572 14740 16584
rect 13740 16544 14740 16572
rect 14734 16532 14740 16544
rect 14792 16572 14798 16584
rect 15120 16572 15148 16612
rect 15657 16609 15669 16612
rect 15703 16609 15715 16643
rect 15657 16603 15715 16609
rect 15856 16584 15884 16680
rect 16853 16643 16911 16649
rect 16853 16609 16865 16643
rect 16899 16640 16911 16643
rect 17126 16640 17132 16652
rect 16899 16612 17132 16640
rect 16899 16609 16911 16612
rect 16853 16603 16911 16609
rect 17126 16600 17132 16612
rect 17184 16600 17190 16652
rect 23569 16643 23627 16649
rect 23569 16609 23581 16643
rect 23615 16640 23627 16643
rect 23842 16640 23848 16652
rect 23615 16612 23848 16640
rect 23615 16609 23627 16612
rect 23569 16603 23627 16609
rect 23842 16600 23848 16612
rect 23900 16600 23906 16652
rect 24118 16600 24124 16652
rect 24176 16640 24182 16652
rect 24581 16643 24639 16649
rect 24581 16640 24593 16643
rect 24176 16612 24593 16640
rect 24176 16600 24182 16612
rect 24581 16609 24593 16612
rect 24627 16609 24639 16643
rect 24581 16603 24639 16609
rect 14792 16544 15148 16572
rect 15749 16575 15807 16581
rect 14792 16532 14798 16544
rect 15749 16541 15761 16575
rect 15795 16541 15807 16575
rect 15749 16535 15807 16541
rect 12897 16507 12955 16513
rect 12897 16473 12909 16507
rect 12943 16504 12955 16507
rect 13722 16504 13728 16516
rect 12943 16476 13728 16504
rect 12943 16473 12955 16476
rect 12897 16467 12955 16473
rect 13722 16464 13728 16476
rect 13780 16464 13786 16516
rect 14090 16464 14096 16516
rect 14148 16504 14154 16516
rect 15289 16507 15347 16513
rect 15289 16504 15301 16507
rect 14148 16476 15301 16504
rect 14148 16464 14154 16476
rect 15289 16473 15301 16476
rect 15335 16473 15347 16507
rect 15289 16467 15347 16473
rect 11238 16436 11244 16448
rect 10520 16408 11244 16436
rect 11238 16396 11244 16408
rect 11296 16396 11302 16448
rect 13078 16396 13084 16448
rect 13136 16436 13142 16448
rect 15764 16436 15792 16535
rect 15838 16532 15844 16584
rect 15896 16572 15902 16584
rect 15896 16544 15989 16572
rect 15896 16532 15902 16544
rect 16758 16436 16764 16448
rect 13136 16408 16764 16436
rect 13136 16396 13142 16408
rect 16758 16396 16764 16408
rect 16816 16436 16822 16448
rect 17218 16436 17224 16448
rect 16816 16408 17224 16436
rect 16816 16396 16822 16408
rect 17218 16396 17224 16408
rect 17276 16396 17282 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2314 16192 2320 16244
rect 2372 16232 2378 16244
rect 2685 16235 2743 16241
rect 2685 16232 2697 16235
rect 2372 16204 2697 16232
rect 2372 16192 2378 16204
rect 2685 16201 2697 16204
rect 2731 16201 2743 16235
rect 2685 16195 2743 16201
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 10229 16235 10287 16241
rect 10229 16232 10241 16235
rect 9732 16204 10241 16232
rect 9732 16192 9738 16204
rect 10229 16201 10241 16204
rect 10275 16201 10287 16235
rect 10229 16195 10287 16201
rect 13630 16192 13636 16244
rect 13688 16232 13694 16244
rect 14277 16235 14335 16241
rect 14277 16232 14289 16235
rect 13688 16204 14289 16232
rect 13688 16192 13694 16204
rect 14277 16201 14289 16204
rect 14323 16201 14335 16235
rect 14734 16232 14740 16244
rect 14695 16204 14740 16232
rect 14277 16195 14335 16201
rect 14734 16192 14740 16204
rect 14792 16192 14798 16244
rect 16758 16232 16764 16244
rect 16719 16204 16764 16232
rect 16758 16192 16764 16204
rect 16816 16192 16822 16244
rect 24118 16192 24124 16244
rect 24176 16232 24182 16244
rect 24673 16235 24731 16241
rect 24673 16232 24685 16235
rect 24176 16204 24685 16232
rect 24176 16192 24182 16204
rect 24673 16201 24685 16204
rect 24719 16201 24731 16235
rect 24673 16195 24731 16201
rect 1581 16167 1639 16173
rect 1581 16133 1593 16167
rect 1627 16164 1639 16167
rect 3050 16164 3056 16176
rect 1627 16136 3056 16164
rect 1627 16133 1639 16136
rect 1581 16127 1639 16133
rect 3050 16124 3056 16136
rect 3108 16124 3114 16176
rect 9766 16164 9772 16176
rect 9727 16136 9772 16164
rect 9766 16124 9772 16136
rect 9824 16164 9830 16176
rect 11330 16164 11336 16176
rect 9824 16136 11336 16164
rect 9824 16124 9830 16136
rect 11330 16124 11336 16136
rect 11388 16124 11394 16176
rect 13265 16167 13323 16173
rect 13265 16133 13277 16167
rect 13311 16164 13323 16167
rect 13998 16164 14004 16176
rect 13311 16136 14004 16164
rect 13311 16133 13323 16136
rect 13265 16127 13323 16133
rect 13998 16124 14004 16136
rect 14056 16124 14062 16176
rect 18230 16164 18236 16176
rect 18191 16136 18236 16164
rect 18230 16124 18236 16136
rect 18288 16124 18294 16176
rect 2424 16068 3096 16096
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 2424 16028 2452 16068
rect 2493 16031 2551 16037
rect 2493 16028 2505 16031
rect 1443 16000 2084 16028
rect 2424 16000 2505 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 2056 15904 2084 16000
rect 2493 15997 2505 16000
rect 2539 15997 2551 16031
rect 2493 15991 2551 15997
rect 3068 15969 3096 16068
rect 8386 16056 8392 16108
rect 8444 16096 8450 16108
rect 9217 16099 9275 16105
rect 9217 16096 9229 16099
rect 8444 16068 9229 16096
rect 8444 16056 8450 16068
rect 9217 16065 9229 16068
rect 9263 16065 9275 16099
rect 9217 16059 9275 16065
rect 10318 16056 10324 16108
rect 10376 16096 10382 16108
rect 10686 16096 10692 16108
rect 10376 16068 10692 16096
rect 10376 16056 10382 16068
rect 10686 16056 10692 16068
rect 10744 16056 10750 16108
rect 10778 16056 10784 16108
rect 10836 16096 10842 16108
rect 13906 16096 13912 16108
rect 10836 16068 10929 16096
rect 13867 16068 13912 16096
rect 10836 16056 10842 16068
rect 13906 16056 13912 16068
rect 13964 16056 13970 16108
rect 14366 16056 14372 16108
rect 14424 16096 14430 16108
rect 14829 16099 14887 16105
rect 14829 16096 14841 16099
rect 14424 16068 14841 16096
rect 14424 16056 14430 16068
rect 14829 16065 14841 16068
rect 14875 16065 14887 16099
rect 14829 16059 14887 16065
rect 10137 16031 10195 16037
rect 10137 15997 10149 16031
rect 10183 16028 10195 16031
rect 10796 16028 10824 16056
rect 10183 16000 10824 16028
rect 15096 16031 15154 16037
rect 10183 15997 10195 16000
rect 10137 15991 10195 15997
rect 15096 15997 15108 16031
rect 15142 16028 15154 16031
rect 15378 16028 15384 16040
rect 15142 16000 15384 16028
rect 15142 15997 15154 16000
rect 15096 15991 15154 15997
rect 15378 15988 15384 16000
rect 15436 15988 15442 16040
rect 17678 15988 17684 16040
rect 17736 16028 17742 16040
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 17736 16000 18061 16028
rect 17736 15988 17742 16000
rect 18049 15997 18061 16000
rect 18095 16028 18107 16031
rect 18509 16031 18567 16037
rect 18509 16028 18521 16031
rect 18095 16000 18521 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 18509 15997 18521 16000
rect 18555 15997 18567 16031
rect 23842 16028 23848 16040
rect 23803 16000 23848 16028
rect 18509 15991 18567 15997
rect 23842 15988 23848 16000
rect 23900 15988 23906 16040
rect 3053 15963 3111 15969
rect 3053 15929 3065 15963
rect 3099 15960 3111 15963
rect 7558 15960 7564 15972
rect 3099 15932 7564 15960
rect 3099 15929 3111 15932
rect 3053 15923 3111 15929
rect 7558 15920 7564 15932
rect 7616 15920 7622 15972
rect 8573 15963 8631 15969
rect 8573 15929 8585 15963
rect 8619 15960 8631 15963
rect 10597 15963 10655 15969
rect 8619 15932 9076 15960
rect 8619 15929 8631 15932
rect 8573 15923 8631 15929
rect 9048 15904 9076 15932
rect 10597 15929 10609 15963
rect 10643 15960 10655 15963
rect 10778 15960 10784 15972
rect 10643 15932 10784 15960
rect 10643 15929 10655 15932
rect 10597 15923 10655 15929
rect 10778 15920 10784 15932
rect 10836 15960 10842 15972
rect 11609 15963 11667 15969
rect 11609 15960 11621 15963
rect 10836 15932 11621 15960
rect 10836 15920 10842 15932
rect 11609 15929 11621 15932
rect 11655 15929 11667 15963
rect 11609 15923 11667 15929
rect 12713 15963 12771 15969
rect 12713 15929 12725 15963
rect 12759 15960 12771 15963
rect 13538 15960 13544 15972
rect 12759 15932 13544 15960
rect 12759 15929 12771 15932
rect 12713 15923 12771 15929
rect 13538 15920 13544 15932
rect 13596 15960 13602 15972
rect 13633 15963 13691 15969
rect 13633 15960 13645 15963
rect 13596 15932 13645 15960
rect 13596 15920 13602 15932
rect 13633 15929 13645 15932
rect 13679 15960 13691 15963
rect 15562 15960 15568 15972
rect 13679 15932 15568 15960
rect 13679 15929 13691 15932
rect 13633 15923 13691 15929
rect 15562 15920 15568 15932
rect 15620 15920 15626 15972
rect 2038 15892 2044 15904
rect 1999 15864 2044 15892
rect 2038 15852 2044 15864
rect 2096 15852 2102 15904
rect 2406 15892 2412 15904
rect 2367 15864 2412 15892
rect 2406 15852 2412 15864
rect 2464 15852 2470 15904
rect 8205 15895 8263 15901
rect 8205 15861 8217 15895
rect 8251 15892 8263 15895
rect 8386 15892 8392 15904
rect 8251 15864 8392 15892
rect 8251 15861 8263 15864
rect 8205 15855 8263 15861
rect 8386 15852 8392 15864
rect 8444 15852 8450 15904
rect 8662 15892 8668 15904
rect 8623 15864 8668 15892
rect 8662 15852 8668 15864
rect 8720 15852 8726 15904
rect 9030 15892 9036 15904
rect 8991 15864 9036 15892
rect 9030 15852 9036 15864
rect 9088 15852 9094 15904
rect 9125 15895 9183 15901
rect 9125 15861 9137 15895
rect 9171 15892 9183 15895
rect 9214 15892 9220 15904
rect 9171 15864 9220 15892
rect 9171 15861 9183 15864
rect 9125 15855 9183 15861
rect 9214 15852 9220 15864
rect 9272 15852 9278 15904
rect 11238 15892 11244 15904
rect 11199 15864 11244 15892
rect 11238 15852 11244 15864
rect 11296 15852 11302 15904
rect 12158 15892 12164 15904
rect 12119 15864 12164 15892
rect 12158 15852 12164 15864
rect 12216 15852 12222 15904
rect 13081 15895 13139 15901
rect 13081 15861 13093 15895
rect 13127 15892 13139 15895
rect 13262 15892 13268 15904
rect 13127 15864 13268 15892
rect 13127 15861 13139 15864
rect 13081 15855 13139 15861
rect 13262 15852 13268 15864
rect 13320 15852 13326 15904
rect 13354 15852 13360 15904
rect 13412 15892 13418 15904
rect 13725 15895 13783 15901
rect 13725 15892 13737 15895
rect 13412 15864 13737 15892
rect 13412 15852 13418 15864
rect 13725 15861 13737 15864
rect 13771 15861 13783 15895
rect 13725 15855 13783 15861
rect 16209 15895 16267 15901
rect 16209 15861 16221 15895
rect 16255 15892 16267 15895
rect 16574 15892 16580 15904
rect 16255 15864 16580 15892
rect 16255 15861 16267 15864
rect 16209 15855 16267 15861
rect 16574 15852 16580 15864
rect 16632 15852 16638 15904
rect 17126 15892 17132 15904
rect 17087 15864 17132 15892
rect 17126 15852 17132 15864
rect 17184 15852 17190 15904
rect 23842 15852 23848 15904
rect 23900 15892 23906 15904
rect 24213 15895 24271 15901
rect 24213 15892 24225 15895
rect 23900 15864 24225 15892
rect 23900 15852 23906 15864
rect 24213 15861 24225 15864
rect 24259 15861 24271 15895
rect 24213 15855 24271 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1394 15648 1400 15700
rect 1452 15688 1458 15700
rect 1581 15691 1639 15697
rect 1581 15688 1593 15691
rect 1452 15660 1593 15688
rect 1452 15648 1458 15660
rect 1581 15657 1593 15660
rect 1627 15657 1639 15691
rect 1581 15651 1639 15657
rect 7929 15691 7987 15697
rect 7929 15657 7941 15691
rect 7975 15688 7987 15691
rect 8389 15691 8447 15697
rect 8389 15688 8401 15691
rect 7975 15660 8401 15688
rect 7975 15657 7987 15660
rect 7929 15651 7987 15657
rect 8389 15657 8401 15660
rect 8435 15688 8447 15691
rect 8662 15688 8668 15700
rect 8435 15660 8668 15688
rect 8435 15657 8447 15660
rect 8389 15651 8447 15657
rect 8662 15648 8668 15660
rect 8720 15648 8726 15700
rect 13814 15648 13820 15700
rect 13872 15688 13878 15700
rect 14090 15688 14096 15700
rect 13872 15660 14096 15688
rect 13872 15648 13878 15660
rect 14090 15648 14096 15660
rect 14148 15648 14154 15700
rect 14366 15648 14372 15700
rect 14424 15688 14430 15700
rect 14829 15691 14887 15697
rect 14829 15688 14841 15691
rect 14424 15660 14841 15688
rect 14424 15648 14430 15660
rect 14829 15657 14841 15660
rect 14875 15657 14887 15691
rect 14829 15651 14887 15657
rect 15378 15648 15384 15700
rect 15436 15688 15442 15700
rect 16301 15691 16359 15697
rect 16301 15688 16313 15691
rect 15436 15660 16313 15688
rect 15436 15648 15442 15660
rect 16301 15657 16313 15660
rect 16347 15657 16359 15691
rect 16301 15651 16359 15657
rect 19426 15648 19432 15700
rect 19484 15688 19490 15700
rect 19613 15691 19671 15697
rect 19613 15688 19625 15691
rect 19484 15660 19625 15688
rect 19484 15648 19490 15660
rect 19613 15657 19625 15660
rect 19659 15657 19671 15691
rect 19613 15651 19671 15657
rect 24670 15648 24676 15700
rect 24728 15688 24734 15700
rect 24765 15691 24823 15697
rect 24765 15688 24777 15691
rect 24728 15660 24777 15688
rect 24728 15648 24734 15660
rect 24765 15657 24777 15660
rect 24811 15657 24823 15691
rect 24765 15651 24823 15657
rect 10597 15623 10655 15629
rect 10597 15589 10609 15623
rect 10643 15620 10655 15623
rect 10934 15623 10992 15629
rect 10934 15620 10946 15623
rect 10643 15592 10946 15620
rect 10643 15589 10655 15592
rect 10597 15583 10655 15589
rect 10934 15589 10946 15592
rect 10980 15620 10992 15623
rect 11054 15620 11060 15632
rect 10980 15592 11060 15620
rect 10980 15589 10992 15592
rect 10934 15583 10992 15589
rect 11054 15580 11060 15592
rect 11112 15620 11118 15632
rect 12621 15623 12679 15629
rect 12621 15620 12633 15623
rect 11112 15592 12633 15620
rect 11112 15580 11118 15592
rect 12621 15589 12633 15592
rect 12667 15589 12679 15623
rect 12621 15583 12679 15589
rect 15657 15623 15715 15629
rect 15657 15589 15669 15623
rect 15703 15620 15715 15623
rect 16022 15620 16028 15632
rect 15703 15592 16028 15620
rect 15703 15589 15715 15592
rect 15657 15583 15715 15589
rect 16022 15580 16028 15592
rect 16080 15580 16086 15632
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 1854 15552 1860 15564
rect 1443 15524 1860 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 1854 15512 1860 15524
rect 1912 15512 1918 15564
rect 8481 15555 8539 15561
rect 8481 15521 8493 15555
rect 8527 15552 8539 15555
rect 8662 15552 8668 15564
rect 8527 15524 8668 15552
rect 8527 15521 8539 15524
rect 8481 15515 8539 15521
rect 8662 15512 8668 15524
rect 8720 15512 8726 15564
rect 11238 15552 11244 15564
rect 10704 15524 11244 15552
rect 8294 15444 8300 15496
rect 8352 15484 8358 15496
rect 8573 15487 8631 15493
rect 8573 15484 8585 15487
rect 8352 15456 8585 15484
rect 8352 15444 8358 15456
rect 8573 15453 8585 15456
rect 8619 15453 8631 15487
rect 9674 15484 9680 15496
rect 9635 15456 9680 15484
rect 8573 15447 8631 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 10226 15444 10232 15496
rect 10284 15484 10290 15496
rect 10704 15493 10732 15524
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 13998 15552 14004 15564
rect 13959 15524 14004 15552
rect 13998 15512 14004 15524
rect 14056 15512 14062 15564
rect 15749 15555 15807 15561
rect 15749 15521 15761 15555
rect 15795 15552 15807 15555
rect 16390 15552 16396 15564
rect 15795 15524 16396 15552
rect 15795 15521 15807 15524
rect 15749 15515 15807 15521
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 17221 15555 17279 15561
rect 17221 15521 17233 15555
rect 17267 15552 17279 15555
rect 17586 15552 17592 15564
rect 17267 15524 17592 15552
rect 17267 15521 17279 15524
rect 17221 15515 17279 15521
rect 17586 15512 17592 15524
rect 17644 15512 17650 15564
rect 18414 15552 18420 15564
rect 18375 15524 18420 15552
rect 18414 15512 18420 15524
rect 18472 15512 18478 15564
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 19429 15555 19487 15561
rect 19429 15552 19441 15555
rect 19392 15524 19441 15552
rect 19392 15512 19398 15524
rect 19429 15521 19441 15524
rect 19475 15521 19487 15555
rect 19429 15515 19487 15521
rect 23569 15555 23627 15561
rect 23569 15521 23581 15555
rect 23615 15552 23627 15555
rect 23934 15552 23940 15564
rect 23615 15524 23940 15552
rect 23615 15521 23627 15524
rect 23569 15515 23627 15521
rect 23934 15512 23940 15524
rect 23992 15512 23998 15564
rect 24581 15555 24639 15561
rect 24581 15521 24593 15555
rect 24627 15552 24639 15555
rect 24854 15552 24860 15564
rect 24627 15524 24860 15552
rect 24627 15521 24639 15524
rect 24581 15515 24639 15521
rect 24854 15512 24860 15524
rect 24912 15512 24918 15564
rect 10689 15487 10747 15493
rect 10689 15484 10701 15487
rect 10284 15456 10701 15484
rect 10284 15444 10290 15456
rect 10689 15453 10701 15456
rect 10735 15453 10747 15487
rect 10689 15447 10747 15453
rect 11882 15444 11888 15496
rect 11940 15484 11946 15496
rect 12250 15484 12256 15496
rect 11940 15456 12256 15484
rect 11940 15444 11946 15456
rect 12250 15444 12256 15456
rect 12308 15484 12314 15496
rect 13265 15487 13323 15493
rect 13265 15484 13277 15487
rect 12308 15456 13277 15484
rect 12308 15444 12314 15456
rect 13265 15453 13277 15456
rect 13311 15484 13323 15487
rect 13354 15484 13360 15496
rect 13311 15456 13360 15484
rect 13311 15453 13323 15456
rect 13265 15447 13323 15453
rect 13354 15444 13360 15456
rect 13412 15444 13418 15496
rect 13538 15444 13544 15496
rect 13596 15484 13602 15496
rect 14277 15487 14335 15493
rect 14277 15484 14289 15487
rect 13596 15456 14289 15484
rect 13596 15444 13602 15456
rect 14277 15453 14289 15456
rect 14323 15484 14335 15487
rect 15378 15484 15384 15496
rect 14323 15456 15384 15484
rect 14323 15453 14335 15456
rect 14277 15447 14335 15453
rect 15378 15444 15384 15456
rect 15436 15444 15442 15496
rect 15838 15444 15844 15496
rect 15896 15484 15902 15496
rect 17310 15484 17316 15496
rect 15896 15456 15941 15484
rect 17271 15456 17316 15484
rect 15896 15444 15902 15456
rect 17310 15444 17316 15456
rect 17368 15444 17374 15496
rect 17405 15487 17463 15493
rect 17405 15453 17417 15487
rect 17451 15453 17463 15487
rect 17405 15447 17463 15453
rect 8018 15416 8024 15428
rect 7979 15388 8024 15416
rect 8018 15376 8024 15388
rect 8076 15376 8082 15428
rect 13630 15416 13636 15428
rect 13591 15388 13636 15416
rect 13630 15376 13636 15388
rect 13688 15376 13694 15428
rect 16574 15376 16580 15428
rect 16632 15416 16638 15428
rect 17420 15416 17448 15447
rect 22278 15444 22284 15496
rect 22336 15484 22342 15496
rect 22557 15487 22615 15493
rect 22557 15484 22569 15487
rect 22336 15456 22569 15484
rect 22336 15444 22342 15456
rect 22557 15453 22569 15456
rect 22603 15453 22615 15487
rect 22557 15447 22615 15453
rect 16632 15388 17448 15416
rect 16632 15376 16638 15388
rect 4246 15348 4252 15360
rect 4207 15320 4252 15348
rect 4246 15308 4252 15320
rect 4304 15308 4310 15360
rect 11330 15308 11336 15360
rect 11388 15348 11394 15360
rect 12069 15351 12127 15357
rect 12069 15348 12081 15351
rect 11388 15320 12081 15348
rect 11388 15308 11394 15320
rect 12069 15317 12081 15320
rect 12115 15317 12127 15351
rect 15286 15348 15292 15360
rect 15247 15320 15292 15348
rect 12069 15311 12127 15317
rect 15286 15308 15292 15320
rect 15344 15308 15350 15360
rect 16482 15308 16488 15360
rect 16540 15348 16546 15360
rect 16761 15351 16819 15357
rect 16761 15348 16773 15351
rect 16540 15320 16773 15348
rect 16540 15308 16546 15320
rect 16761 15317 16773 15320
rect 16807 15348 16819 15351
rect 16853 15351 16911 15357
rect 16853 15348 16865 15351
rect 16807 15320 16865 15348
rect 16807 15317 16819 15320
rect 16761 15311 16819 15317
rect 16853 15317 16865 15320
rect 16899 15317 16911 15351
rect 16853 15311 16911 15317
rect 18230 15308 18236 15360
rect 18288 15348 18294 15360
rect 18601 15351 18659 15357
rect 18601 15348 18613 15351
rect 18288 15320 18613 15348
rect 18288 15308 18294 15320
rect 18601 15317 18613 15320
rect 18647 15317 18659 15351
rect 18601 15311 18659 15317
rect 22462 15308 22468 15360
rect 22520 15348 22526 15360
rect 23753 15351 23811 15357
rect 23753 15348 23765 15351
rect 22520 15320 23765 15348
rect 22520 15308 22526 15320
rect 23753 15317 23765 15320
rect 23799 15317 23811 15351
rect 23753 15311 23811 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1946 15104 1952 15156
rect 2004 15144 2010 15156
rect 2041 15147 2099 15153
rect 2041 15144 2053 15147
rect 2004 15116 2053 15144
rect 2004 15104 2010 15116
rect 2041 15113 2053 15116
rect 2087 15113 2099 15147
rect 2041 15107 2099 15113
rect 7469 15147 7527 15153
rect 7469 15113 7481 15147
rect 7515 15144 7527 15147
rect 8294 15144 8300 15156
rect 7515 15116 8300 15144
rect 7515 15113 7527 15116
rect 7469 15107 7527 15113
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 9674 15104 9680 15156
rect 9732 15144 9738 15156
rect 9861 15147 9919 15153
rect 9861 15144 9873 15147
rect 9732 15116 9873 15144
rect 9732 15104 9738 15116
rect 9861 15113 9873 15116
rect 9907 15144 9919 15147
rect 13538 15144 13544 15156
rect 9907 15116 11192 15144
rect 13499 15116 13544 15144
rect 9907 15113 9919 15116
rect 9861 15107 9919 15113
rect 10778 15076 10784 15088
rect 10739 15048 10784 15076
rect 10778 15036 10784 15048
rect 10836 15036 10842 15088
rect 3789 15011 3847 15017
rect 3789 14977 3801 15011
rect 3835 15008 3847 15011
rect 4433 15011 4491 15017
rect 4433 15008 4445 15011
rect 3835 14980 4445 15008
rect 3835 14977 3847 14980
rect 3789 14971 3847 14977
rect 4433 14977 4445 14980
rect 4479 15008 4491 15011
rect 5718 15008 5724 15020
rect 4479 14980 5724 15008
rect 4479 14977 4491 14980
rect 4433 14971 4491 14977
rect 5718 14968 5724 14980
rect 5776 14968 5782 15020
rect 1857 14943 1915 14949
rect 1857 14909 1869 14943
rect 1903 14940 1915 14943
rect 4246 14940 4252 14952
rect 1903 14912 2544 14940
rect 4207 14912 4252 14940
rect 1903 14909 1915 14912
rect 1857 14903 1915 14909
rect 2516 14816 2544 14912
rect 4246 14900 4252 14912
rect 4304 14900 4310 14952
rect 11164 14949 11192 15116
rect 13538 15104 13544 15116
rect 13596 15104 13602 15156
rect 13909 15147 13967 15153
rect 13909 15113 13921 15147
rect 13955 15144 13967 15147
rect 14366 15144 14372 15156
rect 13955 15116 14372 15144
rect 13955 15113 13967 15116
rect 13909 15107 13967 15113
rect 12802 15036 12808 15088
rect 12860 15076 12866 15088
rect 14016 15076 14044 15116
rect 14366 15104 14372 15116
rect 14424 15104 14430 15156
rect 16022 15144 16028 15156
rect 15983 15116 16028 15144
rect 16022 15104 16028 15116
rect 16080 15104 16086 15156
rect 16114 15104 16120 15156
rect 16172 15144 16178 15156
rect 16390 15144 16396 15156
rect 16172 15116 16396 15144
rect 16172 15104 16178 15116
rect 16390 15104 16396 15116
rect 16448 15104 16454 15156
rect 17310 15144 17316 15156
rect 17271 15116 17316 15144
rect 17310 15104 17316 15116
rect 17368 15104 17374 15156
rect 24762 15144 24768 15156
rect 24723 15116 24768 15144
rect 24762 15104 24768 15116
rect 24820 15104 24826 15156
rect 12860 15048 14044 15076
rect 12860 15036 12866 15048
rect 11330 15008 11336 15020
rect 11291 14980 11336 15008
rect 11330 14968 11336 14980
rect 11388 14968 11394 15020
rect 11698 14968 11704 15020
rect 11756 15008 11762 15020
rect 11885 15011 11943 15017
rect 11885 15008 11897 15011
rect 11756 14980 11897 15008
rect 11756 14968 11762 14980
rect 11885 14977 11897 14980
rect 11931 15008 11943 15011
rect 12618 15008 12624 15020
rect 11931 14980 12624 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 12618 14968 12624 14980
rect 12676 14968 12682 15020
rect 12986 15008 12992 15020
rect 12947 14980 12992 15008
rect 12986 14968 12992 14980
rect 13044 14968 13050 15020
rect 14016 15017 14044 15048
rect 19337 15079 19395 15085
rect 19337 15045 19349 15079
rect 19383 15076 19395 15079
rect 20438 15076 20444 15088
rect 19383 15048 20444 15076
rect 19383 15045 19395 15048
rect 19337 15039 19395 15045
rect 20438 15036 20444 15048
rect 20496 15036 20502 15088
rect 14001 15011 14059 15017
rect 14001 14977 14013 15011
rect 14047 14977 14059 15011
rect 14001 14971 14059 14977
rect 7929 14943 7987 14949
rect 7929 14940 7941 14943
rect 7760 14912 7941 14940
rect 4341 14875 4399 14881
rect 4341 14872 4353 14875
rect 3344 14844 4353 14872
rect 1673 14807 1731 14813
rect 1673 14773 1685 14807
rect 1719 14804 1731 14807
rect 1854 14804 1860 14816
rect 1719 14776 1860 14804
rect 1719 14773 1731 14776
rect 1673 14767 1731 14773
rect 1854 14764 1860 14776
rect 1912 14764 1918 14816
rect 2498 14804 2504 14816
rect 2459 14776 2504 14804
rect 2498 14764 2504 14776
rect 2556 14764 2562 14816
rect 3050 14764 3056 14816
rect 3108 14804 3114 14816
rect 3344 14813 3372 14844
rect 4341 14841 4353 14844
rect 4387 14841 4399 14875
rect 4341 14835 4399 14841
rect 3329 14807 3387 14813
rect 3329 14804 3341 14807
rect 3108 14776 3341 14804
rect 3108 14764 3114 14776
rect 3329 14773 3341 14776
rect 3375 14773 3387 14807
rect 3878 14804 3884 14816
rect 3839 14776 3884 14804
rect 3329 14767 3387 14773
rect 3878 14764 3884 14776
rect 3936 14764 3942 14816
rect 6914 14804 6920 14816
rect 6875 14776 6920 14804
rect 6914 14764 6920 14776
rect 6972 14764 6978 14816
rect 7098 14764 7104 14816
rect 7156 14804 7162 14816
rect 7760 14813 7788 14912
rect 7929 14909 7941 14912
rect 7975 14909 7987 14943
rect 7929 14903 7987 14909
rect 11149 14943 11207 14949
rect 11149 14909 11161 14943
rect 11195 14909 11207 14943
rect 16298 14940 16304 14952
rect 11149 14903 11207 14909
rect 13004 14912 16304 14940
rect 8196 14875 8254 14881
rect 8196 14841 8208 14875
rect 8242 14872 8254 14875
rect 8570 14872 8576 14884
rect 8242 14844 8576 14872
rect 8242 14841 8254 14844
rect 8196 14835 8254 14841
rect 8570 14832 8576 14844
rect 8628 14832 8634 14884
rect 9674 14832 9680 14884
rect 9732 14872 9738 14884
rect 10226 14872 10232 14884
rect 9732 14844 10232 14872
rect 9732 14832 9738 14844
rect 10226 14832 10232 14844
rect 10284 14832 10290 14884
rect 12253 14875 12311 14881
rect 12253 14841 12265 14875
rect 12299 14872 12311 14875
rect 12342 14872 12348 14884
rect 12299 14844 12348 14872
rect 12299 14841 12311 14844
rect 12253 14835 12311 14841
rect 12342 14832 12348 14844
rect 12400 14872 12406 14884
rect 12805 14875 12863 14881
rect 12805 14872 12817 14875
rect 12400 14844 12817 14872
rect 12400 14832 12406 14844
rect 12805 14841 12817 14844
rect 12851 14841 12863 14875
rect 12805 14835 12863 14841
rect 12897 14875 12955 14881
rect 12897 14841 12909 14875
rect 12943 14872 12955 14875
rect 13004 14872 13032 14912
rect 16298 14900 16304 14912
rect 16356 14900 16362 14952
rect 16482 14940 16488 14952
rect 16443 14912 16488 14940
rect 16482 14900 16488 14912
rect 16540 14900 16546 14952
rect 18874 14900 18880 14952
rect 18932 14940 18938 14952
rect 19153 14943 19211 14949
rect 19153 14940 19165 14943
rect 18932 14912 19165 14940
rect 18932 14900 18938 14912
rect 19153 14909 19165 14912
rect 19199 14909 19211 14943
rect 19153 14903 19211 14909
rect 12943 14844 13032 14872
rect 12943 14841 12955 14844
rect 12897 14835 12955 14841
rect 7745 14807 7803 14813
rect 7745 14804 7757 14807
rect 7156 14776 7757 14804
rect 7156 14764 7162 14776
rect 7745 14773 7757 14776
rect 7791 14773 7803 14807
rect 7745 14767 7803 14773
rect 9309 14807 9367 14813
rect 9309 14773 9321 14807
rect 9355 14804 9367 14807
rect 9950 14804 9956 14816
rect 9355 14776 9956 14804
rect 9355 14773 9367 14776
rect 9309 14767 9367 14773
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 10689 14807 10747 14813
rect 10689 14773 10701 14807
rect 10735 14804 10747 14807
rect 11238 14804 11244 14816
rect 10735 14776 11244 14804
rect 10735 14773 10747 14776
rect 10689 14767 10747 14773
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 12434 14764 12440 14816
rect 12492 14804 12498 14816
rect 12492 14776 12537 14804
rect 12492 14764 12498 14776
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 12912 14804 12940 14835
rect 14090 14832 14096 14884
rect 14148 14872 14154 14884
rect 14246 14875 14304 14881
rect 14246 14872 14258 14875
rect 14148 14844 14258 14872
rect 14148 14832 14154 14844
rect 14246 14841 14258 14844
rect 14292 14872 14304 14875
rect 16574 14872 16580 14884
rect 14292 14844 16580 14872
rect 14292 14841 14304 14844
rect 14246 14835 14304 14841
rect 16574 14832 16580 14844
rect 16632 14872 16638 14884
rect 16945 14875 17003 14881
rect 16945 14872 16957 14875
rect 16632 14844 16957 14872
rect 16632 14832 16638 14844
rect 16945 14841 16957 14844
rect 16991 14841 17003 14875
rect 16945 14835 17003 14841
rect 17954 14832 17960 14884
rect 18012 14872 18018 14884
rect 18414 14872 18420 14884
rect 18012 14844 18420 14872
rect 18012 14832 18018 14844
rect 18414 14832 18420 14844
rect 18472 14872 18478 14884
rect 18509 14875 18567 14881
rect 18509 14872 18521 14875
rect 18472 14844 18521 14872
rect 18472 14832 18478 14844
rect 18509 14841 18521 14844
rect 18555 14841 18567 14875
rect 19168 14872 19196 14903
rect 19334 14900 19340 14952
rect 19392 14940 19398 14952
rect 19613 14943 19671 14949
rect 19613 14940 19625 14943
rect 19392 14912 19625 14940
rect 19392 14900 19398 14912
rect 19613 14909 19625 14912
rect 19659 14909 19671 14943
rect 20346 14940 20352 14952
rect 20307 14912 20352 14940
rect 19613 14903 19671 14909
rect 20346 14900 20352 14912
rect 20404 14940 20410 14952
rect 20809 14943 20867 14949
rect 20809 14940 20821 14943
rect 20404 14912 20821 14940
rect 20404 14900 20410 14912
rect 20809 14909 20821 14912
rect 20855 14909 20867 14943
rect 20809 14903 20867 14909
rect 22557 14943 22615 14949
rect 22557 14909 22569 14943
rect 22603 14940 22615 14943
rect 22603 14912 23152 14940
rect 22603 14909 22615 14912
rect 22557 14903 22615 14909
rect 19981 14875 20039 14881
rect 19981 14872 19993 14875
rect 19168 14844 19993 14872
rect 18509 14835 18567 14841
rect 19981 14841 19993 14844
rect 20027 14841 20039 14875
rect 19981 14835 20039 14841
rect 12676 14776 12940 14804
rect 12676 14764 12682 14776
rect 15194 14764 15200 14816
rect 15252 14804 15258 14816
rect 15381 14807 15439 14813
rect 15381 14804 15393 14807
rect 15252 14776 15393 14804
rect 15252 14764 15258 14776
rect 15381 14773 15393 14776
rect 15427 14773 15439 14807
rect 15381 14767 15439 14773
rect 16669 14807 16727 14813
rect 16669 14773 16681 14807
rect 16715 14804 16727 14807
rect 16850 14804 16856 14816
rect 16715 14776 16856 14804
rect 16715 14773 16727 14776
rect 16669 14767 16727 14773
rect 16850 14764 16856 14776
rect 16908 14764 16914 14816
rect 17586 14764 17592 14816
rect 17644 14804 17650 14816
rect 17681 14807 17739 14813
rect 17681 14804 17693 14807
rect 17644 14776 17693 14804
rect 17644 14764 17650 14776
rect 17681 14773 17693 14776
rect 17727 14773 17739 14807
rect 17681 14767 17739 14773
rect 18049 14807 18107 14813
rect 18049 14773 18061 14807
rect 18095 14804 18107 14807
rect 18690 14804 18696 14816
rect 18095 14776 18696 14804
rect 18095 14773 18107 14776
rect 18049 14767 18107 14773
rect 18690 14764 18696 14776
rect 18748 14764 18754 14816
rect 20530 14804 20536 14816
rect 20491 14776 20536 14804
rect 20530 14764 20536 14776
rect 20588 14764 20594 14816
rect 21542 14804 21548 14816
rect 21503 14776 21548 14804
rect 21542 14764 21548 14776
rect 21600 14764 21606 14816
rect 22738 14804 22744 14816
rect 22699 14776 22744 14804
rect 22738 14764 22744 14776
rect 22796 14764 22802 14816
rect 23124 14813 23152 14912
rect 24118 14900 24124 14952
rect 24176 14940 24182 14952
rect 24581 14943 24639 14949
rect 24581 14940 24593 14943
rect 24176 14912 24593 14940
rect 24176 14900 24182 14912
rect 24581 14909 24593 14912
rect 24627 14940 24639 14943
rect 25133 14943 25191 14949
rect 25133 14940 25145 14943
rect 24627 14912 25145 14940
rect 24627 14909 24639 14912
rect 24581 14903 24639 14909
rect 25133 14909 25145 14912
rect 25179 14909 25191 14943
rect 25133 14903 25191 14909
rect 23566 14832 23572 14884
rect 23624 14872 23630 14884
rect 24946 14872 24952 14884
rect 23624 14844 24952 14872
rect 23624 14832 23630 14844
rect 24946 14832 24952 14844
rect 25004 14832 25010 14884
rect 23109 14807 23167 14813
rect 23109 14773 23121 14807
rect 23155 14804 23167 14807
rect 23198 14804 23204 14816
rect 23155 14776 23204 14804
rect 23155 14773 23167 14776
rect 23109 14767 23167 14773
rect 23198 14764 23204 14776
rect 23256 14764 23262 14816
rect 23934 14804 23940 14816
rect 23895 14776 23940 14804
rect 23934 14764 23940 14776
rect 23992 14764 23998 14816
rect 24118 14764 24124 14816
rect 24176 14804 24182 14816
rect 24397 14807 24455 14813
rect 24397 14804 24409 14807
rect 24176 14776 24409 14804
rect 24176 14764 24182 14776
rect 24397 14773 24409 14776
rect 24443 14804 24455 14807
rect 24854 14804 24860 14816
rect 24443 14776 24860 14804
rect 24443 14773 24455 14776
rect 24397 14767 24455 14773
rect 24854 14764 24860 14776
rect 24912 14764 24918 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1578 14600 1584 14612
rect 1539 14572 1584 14600
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 2498 14560 2504 14612
rect 2556 14600 2562 14612
rect 2685 14603 2743 14609
rect 2685 14600 2697 14603
rect 2556 14572 2697 14600
rect 2556 14560 2562 14572
rect 2685 14569 2697 14572
rect 2731 14569 2743 14603
rect 2685 14563 2743 14569
rect 4065 14603 4123 14609
rect 4065 14569 4077 14603
rect 4111 14600 4123 14603
rect 4246 14600 4252 14612
rect 4111 14572 4252 14600
rect 4111 14569 4123 14572
rect 4065 14563 4123 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 11054 14600 11060 14612
rect 11015 14572 11060 14600
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 11330 14560 11336 14612
rect 11388 14600 11394 14612
rect 11609 14603 11667 14609
rect 11609 14600 11621 14603
rect 11388 14572 11621 14600
rect 11388 14560 11394 14572
rect 11609 14569 11621 14572
rect 11655 14569 11667 14603
rect 13722 14600 13728 14612
rect 13683 14572 13728 14600
rect 11609 14563 11667 14569
rect 13722 14560 13728 14572
rect 13780 14560 13786 14612
rect 13998 14560 14004 14612
rect 14056 14600 14062 14612
rect 14645 14603 14703 14609
rect 14645 14600 14657 14603
rect 14056 14572 14657 14600
rect 14056 14560 14062 14572
rect 14645 14569 14657 14572
rect 14691 14569 14703 14603
rect 14645 14563 14703 14569
rect 14826 14560 14832 14612
rect 14884 14600 14890 14612
rect 15013 14603 15071 14609
rect 15013 14600 15025 14603
rect 14884 14572 15025 14600
rect 14884 14560 14890 14572
rect 15013 14569 15025 14572
rect 15059 14569 15071 14603
rect 15013 14563 15071 14569
rect 15286 14560 15292 14612
rect 15344 14600 15350 14612
rect 15749 14603 15807 14609
rect 15749 14600 15761 14603
rect 15344 14572 15761 14600
rect 15344 14560 15350 14572
rect 15749 14569 15761 14572
rect 15795 14600 15807 14603
rect 15838 14600 15844 14612
rect 15795 14572 15844 14600
rect 15795 14569 15807 14572
rect 15749 14563 15807 14569
rect 15838 14560 15844 14572
rect 15896 14560 15902 14612
rect 17310 14600 17316 14612
rect 17223 14572 17316 14600
rect 17310 14560 17316 14572
rect 17368 14600 17374 14612
rect 17770 14600 17776 14612
rect 17368 14572 17776 14600
rect 17368 14560 17374 14572
rect 17770 14560 17776 14572
rect 17828 14560 17834 14612
rect 18598 14600 18604 14612
rect 18559 14572 18604 14600
rect 18598 14560 18604 14572
rect 18656 14560 18662 14612
rect 24210 14560 24216 14612
rect 24268 14600 24274 14612
rect 24765 14603 24823 14609
rect 24765 14600 24777 14603
rect 24268 14572 24777 14600
rect 24268 14560 24274 14572
rect 24765 14569 24777 14572
rect 24811 14569 24823 14603
rect 24765 14563 24823 14569
rect 3878 14532 3884 14544
rect 2516 14504 3884 14532
rect 1394 14464 1400 14476
rect 1355 14436 1400 14464
rect 1394 14424 1400 14436
rect 1452 14424 1458 14476
rect 2516 14473 2544 14504
rect 3878 14492 3884 14504
rect 3936 14492 3942 14544
rect 4154 14492 4160 14544
rect 4212 14532 4218 14544
rect 4212 14504 5672 14532
rect 4212 14492 4218 14504
rect 2409 14467 2467 14473
rect 2409 14433 2421 14467
rect 2455 14464 2467 14467
rect 2501 14467 2559 14473
rect 2501 14464 2513 14467
rect 2455 14436 2513 14464
rect 2455 14433 2467 14436
rect 2409 14427 2467 14433
rect 2501 14433 2513 14436
rect 2547 14433 2559 14467
rect 2501 14427 2559 14433
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 3510 14464 3516 14476
rect 2832 14436 3516 14464
rect 2832 14424 2838 14436
rect 3510 14424 3516 14436
rect 3568 14424 3574 14476
rect 4430 14464 4436 14476
rect 4391 14436 4436 14464
rect 4430 14424 4436 14436
rect 4488 14424 4494 14476
rect 5644 14473 5672 14504
rect 5718 14492 5724 14544
rect 5776 14532 5782 14544
rect 5874 14535 5932 14541
rect 5874 14532 5886 14535
rect 5776 14504 5886 14532
rect 5776 14492 5782 14504
rect 5874 14501 5886 14504
rect 5920 14501 5932 14535
rect 14090 14532 14096 14544
rect 14051 14504 14096 14532
rect 5874 14495 5932 14501
rect 14090 14492 14096 14504
rect 14148 14492 14154 14544
rect 15654 14532 15660 14544
rect 15615 14504 15660 14532
rect 15654 14492 15660 14504
rect 15712 14492 15718 14544
rect 16574 14492 16580 14544
rect 16632 14532 16638 14544
rect 16632 14504 17356 14532
rect 16632 14492 16638 14504
rect 9950 14473 9956 14476
rect 4525 14467 4583 14473
rect 4525 14433 4537 14467
rect 4571 14433 4583 14467
rect 4525 14427 4583 14433
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14433 5687 14467
rect 9944 14464 9956 14473
rect 9911 14436 9956 14464
rect 5629 14427 5687 14433
rect 9944 14427 9956 14436
rect 4540 14396 4568 14427
rect 9950 14424 9956 14427
rect 10008 14424 10014 14476
rect 12250 14424 12256 14476
rect 12308 14464 12314 14476
rect 12529 14467 12587 14473
rect 12529 14464 12541 14467
rect 12308 14436 12541 14464
rect 12308 14424 12314 14436
rect 12529 14433 12541 14436
rect 12575 14433 12587 14467
rect 14182 14464 14188 14476
rect 14143 14436 14188 14464
rect 12529 14427 12587 14433
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 17218 14464 17224 14476
rect 17179 14436 17224 14464
rect 17218 14424 17224 14436
rect 17276 14424 17282 14476
rect 17328 14464 17356 14504
rect 17328 14436 17448 14464
rect 3804 14368 4568 14396
rect 4709 14399 4767 14405
rect 2774 14288 2780 14340
rect 2832 14328 2838 14340
rect 3804 14337 3832 14368
rect 4709 14365 4721 14399
rect 4755 14365 4767 14399
rect 8202 14396 8208 14408
rect 8163 14368 8208 14396
rect 4709 14359 4767 14365
rect 3789 14331 3847 14337
rect 3789 14328 3801 14331
rect 2832 14300 3801 14328
rect 2832 14288 2838 14300
rect 3789 14297 3801 14300
rect 3835 14297 3847 14331
rect 3789 14291 3847 14297
rect 4522 14288 4528 14340
rect 4580 14328 4586 14340
rect 4724 14328 4752 14359
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 9674 14396 9680 14408
rect 9635 14368 9680 14396
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 12618 14396 12624 14408
rect 12579 14368 12624 14396
rect 12618 14356 12624 14368
rect 12676 14356 12682 14408
rect 12713 14399 12771 14405
rect 12713 14365 12725 14399
rect 12759 14396 12771 14399
rect 12986 14396 12992 14408
rect 12759 14368 12992 14396
rect 12759 14365 12771 14368
rect 12713 14359 12771 14365
rect 5077 14331 5135 14337
rect 5077 14328 5089 14331
rect 4580 14300 5089 14328
rect 4580 14288 4586 14300
rect 5077 14297 5089 14300
rect 5123 14297 5135 14331
rect 5077 14291 5135 14297
rect 8021 14331 8079 14337
rect 8021 14297 8033 14331
rect 8067 14328 8079 14331
rect 8570 14328 8576 14340
rect 8067 14300 8576 14328
rect 8067 14297 8079 14300
rect 8021 14291 8079 14297
rect 8570 14288 8576 14300
rect 8628 14288 8634 14340
rect 11054 14288 11060 14340
rect 11112 14328 11118 14340
rect 12728 14328 12756 14359
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 13265 14399 13323 14405
rect 13265 14365 13277 14399
rect 13311 14396 13323 14399
rect 13354 14396 13360 14408
rect 13311 14368 13360 14396
rect 13311 14365 13323 14368
rect 13265 14359 13323 14365
rect 13354 14356 13360 14368
rect 13412 14396 13418 14408
rect 15194 14396 15200 14408
rect 13412 14368 15200 14396
rect 13412 14356 13418 14368
rect 15194 14356 15200 14368
rect 15252 14356 15258 14408
rect 15378 14356 15384 14408
rect 15436 14396 15442 14408
rect 15746 14396 15752 14408
rect 15436 14368 15752 14396
rect 15436 14356 15442 14368
rect 15746 14356 15752 14368
rect 15804 14396 15810 14408
rect 17420 14405 17448 14436
rect 17770 14424 17776 14476
rect 17828 14464 17834 14476
rect 18417 14467 18475 14473
rect 18417 14464 18429 14467
rect 17828 14436 18429 14464
rect 17828 14424 17834 14436
rect 18417 14433 18429 14436
rect 18463 14464 18475 14467
rect 19426 14464 19432 14476
rect 18463 14436 19432 14464
rect 18463 14433 18475 14436
rect 18417 14427 18475 14433
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 19521 14467 19579 14473
rect 19521 14433 19533 14467
rect 19567 14464 19579 14467
rect 20162 14464 20168 14476
rect 19567 14436 20168 14464
rect 19567 14433 19579 14436
rect 19521 14427 19579 14433
rect 20162 14424 20168 14436
rect 20220 14424 20226 14476
rect 20622 14424 20628 14476
rect 20680 14464 20686 14476
rect 20901 14467 20959 14473
rect 20901 14464 20913 14467
rect 20680 14436 20913 14464
rect 20680 14424 20686 14436
rect 20901 14433 20913 14436
rect 20947 14433 20959 14467
rect 22554 14464 22560 14476
rect 22515 14436 22560 14464
rect 20901 14427 20959 14433
rect 22554 14424 22560 14436
rect 22612 14424 22618 14476
rect 23566 14464 23572 14476
rect 23527 14436 23572 14464
rect 23566 14424 23572 14436
rect 23624 14424 23630 14476
rect 24581 14467 24639 14473
rect 24581 14433 24593 14467
rect 24627 14464 24639 14467
rect 24670 14464 24676 14476
rect 24627 14436 24676 14464
rect 24627 14433 24639 14436
rect 24581 14427 24639 14433
rect 24670 14424 24676 14436
rect 24728 14424 24734 14476
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 15804 14368 15853 14396
rect 15804 14356 15810 14368
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 17405 14399 17463 14405
rect 17405 14365 17417 14399
rect 17451 14365 17463 14399
rect 17405 14359 17463 14365
rect 11112 14300 12756 14328
rect 15289 14331 15347 14337
rect 11112 14288 11118 14300
rect 15289 14297 15301 14331
rect 15335 14328 15347 14331
rect 17586 14328 17592 14340
rect 15335 14300 17592 14328
rect 15335 14297 15347 14300
rect 15289 14291 15347 14297
rect 17586 14288 17592 14300
rect 17644 14288 17650 14340
rect 1946 14260 1952 14272
rect 1907 14232 1952 14260
rect 1946 14220 1952 14232
rect 2004 14220 2010 14272
rect 3142 14260 3148 14272
rect 3103 14232 3148 14260
rect 3142 14220 3148 14232
rect 3200 14220 3206 14272
rect 3418 14260 3424 14272
rect 3379 14232 3424 14260
rect 3418 14220 3424 14232
rect 3476 14220 3482 14272
rect 7009 14263 7067 14269
rect 7009 14229 7021 14263
rect 7055 14260 7067 14263
rect 7282 14260 7288 14272
rect 7055 14232 7288 14260
rect 7055 14229 7067 14232
rect 7009 14223 7067 14229
rect 7282 14220 7288 14232
rect 7340 14220 7346 14272
rect 8662 14260 8668 14272
rect 8623 14232 8668 14260
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 11974 14260 11980 14272
rect 11935 14232 11980 14260
rect 11974 14220 11980 14232
rect 12032 14260 12038 14272
rect 12161 14263 12219 14269
rect 12161 14260 12173 14263
rect 12032 14232 12173 14260
rect 12032 14220 12038 14232
rect 12161 14229 12173 14232
rect 12207 14229 12219 14263
rect 14366 14260 14372 14272
rect 14327 14232 14372 14260
rect 12161 14223 12219 14229
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 16390 14260 16396 14272
rect 16351 14232 16396 14260
rect 16390 14220 16396 14232
rect 16448 14220 16454 14272
rect 16574 14220 16580 14272
rect 16632 14260 16638 14272
rect 16669 14263 16727 14269
rect 16669 14260 16681 14263
rect 16632 14232 16681 14260
rect 16632 14220 16638 14232
rect 16669 14229 16681 14232
rect 16715 14229 16727 14263
rect 16669 14223 16727 14229
rect 16758 14220 16764 14272
rect 16816 14260 16822 14272
rect 16853 14263 16911 14269
rect 16853 14260 16865 14263
rect 16816 14232 16865 14260
rect 16816 14220 16822 14232
rect 16853 14229 16865 14232
rect 16899 14229 16911 14263
rect 16853 14223 16911 14229
rect 18141 14263 18199 14269
rect 18141 14229 18153 14263
rect 18187 14260 18199 14263
rect 18414 14260 18420 14272
rect 18187 14232 18420 14260
rect 18187 14229 18199 14232
rect 18141 14223 18199 14229
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 19061 14263 19119 14269
rect 19061 14229 19073 14263
rect 19107 14260 19119 14263
rect 19242 14260 19248 14272
rect 19107 14232 19248 14260
rect 19107 14229 19119 14232
rect 19061 14223 19119 14229
rect 19242 14220 19248 14232
rect 19300 14220 19306 14272
rect 19705 14263 19763 14269
rect 19705 14229 19717 14263
rect 19751 14260 19763 14263
rect 19978 14260 19984 14272
rect 19751 14232 19984 14260
rect 19751 14229 19763 14232
rect 19705 14223 19763 14229
rect 19978 14220 19984 14232
rect 20036 14220 20042 14272
rect 20254 14220 20260 14272
rect 20312 14260 20318 14272
rect 21085 14263 21143 14269
rect 21085 14260 21097 14263
rect 20312 14232 21097 14260
rect 20312 14220 20318 14232
rect 21085 14229 21097 14232
rect 21131 14229 21143 14263
rect 21085 14223 21143 14229
rect 22741 14263 22799 14269
rect 22741 14229 22753 14263
rect 22787 14260 22799 14263
rect 22922 14260 22928 14272
rect 22787 14232 22928 14260
rect 22787 14229 22799 14232
rect 22741 14223 22799 14229
rect 22922 14220 22928 14232
rect 22980 14220 22986 14272
rect 23750 14260 23756 14272
rect 23711 14232 23756 14260
rect 23750 14220 23756 14232
rect 23808 14220 23814 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1394 14016 1400 14068
rect 1452 14056 1458 14068
rect 2222 14056 2228 14068
rect 1452 14028 2228 14056
rect 1452 14016 1458 14028
rect 2222 14016 2228 14028
rect 2280 14056 2286 14068
rect 2317 14059 2375 14065
rect 2317 14056 2329 14059
rect 2280 14028 2329 14056
rect 2280 14016 2286 14028
rect 2317 14025 2329 14028
rect 2363 14025 2375 14059
rect 2317 14019 2375 14025
rect 3789 14059 3847 14065
rect 3789 14025 3801 14059
rect 3835 14056 3847 14059
rect 4430 14056 4436 14068
rect 3835 14028 4436 14056
rect 3835 14025 3847 14028
rect 3789 14019 3847 14025
rect 4430 14016 4436 14028
rect 4488 14016 4494 14068
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 5629 14059 5687 14065
rect 5629 14056 5641 14059
rect 5592 14028 5641 14056
rect 5592 14016 5598 14028
rect 5629 14025 5641 14028
rect 5675 14056 5687 14059
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 5675 14028 6561 14056
rect 5675 14025 5687 14028
rect 5629 14019 5687 14025
rect 6549 14025 6561 14028
rect 6595 14025 6607 14059
rect 9674 14056 9680 14068
rect 9635 14028 9680 14056
rect 6549 14019 6607 14025
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 10505 14059 10563 14065
rect 10505 14025 10517 14059
rect 10551 14056 10563 14059
rect 10686 14056 10692 14068
rect 10551 14028 10692 14056
rect 10551 14025 10563 14028
rect 10505 14019 10563 14025
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 11054 14016 11060 14068
rect 11112 14016 11118 14068
rect 12250 14056 12256 14068
rect 12211 14028 12256 14056
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 15381 14059 15439 14065
rect 15381 14025 15393 14059
rect 15427 14056 15439 14059
rect 15654 14056 15660 14068
rect 15427 14028 15660 14056
rect 15427 14025 15439 14028
rect 15381 14019 15439 14025
rect 15654 14016 15660 14028
rect 15712 14016 15718 14068
rect 15746 14016 15752 14068
rect 15804 14056 15810 14068
rect 17221 14059 17279 14065
rect 15804 14028 15849 14056
rect 15804 14016 15810 14028
rect 17221 14025 17233 14059
rect 17267 14056 17279 14059
rect 17310 14056 17316 14068
rect 17267 14028 17316 14056
rect 17267 14025 17279 14028
rect 17221 14019 17279 14025
rect 17310 14016 17316 14028
rect 17368 14016 17374 14068
rect 18046 14056 18052 14068
rect 18007 14028 18052 14056
rect 18046 14016 18052 14028
rect 18104 14016 18110 14068
rect 19426 14056 19432 14068
rect 19387 14028 19432 14056
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 21177 14059 21235 14065
rect 21177 14025 21189 14059
rect 21223 14056 21235 14059
rect 22186 14056 22192 14068
rect 21223 14028 22192 14056
rect 21223 14025 21235 14028
rect 21177 14019 21235 14025
rect 22186 14016 22192 14028
rect 22244 14016 22250 14068
rect 22554 14016 22560 14068
rect 22612 14056 22618 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 22612 14028 23397 14056
rect 22612 14016 22618 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 23385 14019 23443 14025
rect 1581 13991 1639 13997
rect 1581 13957 1593 13991
rect 1627 13988 1639 13991
rect 2130 13988 2136 14000
rect 1627 13960 2136 13988
rect 1627 13957 1639 13960
rect 1581 13951 1639 13957
rect 2130 13948 2136 13960
rect 2188 13948 2194 14000
rect 4154 13988 4160 14000
rect 4115 13960 4160 13988
rect 4154 13948 4160 13960
rect 4212 13988 4218 14000
rect 11072 13988 11100 14016
rect 12618 13988 12624 14000
rect 4212 13960 4292 13988
rect 11072 13960 11744 13988
rect 12579 13960 12624 13988
rect 4212 13948 4218 13960
rect 4264 13929 4292 13960
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13920 9459 13923
rect 10962 13920 10968 13932
rect 9447 13892 10968 13920
rect 9447 13889 9459 13892
rect 9401 13883 9459 13889
rect 10962 13880 10968 13892
rect 11020 13880 11026 13932
rect 11054 13880 11060 13932
rect 11112 13920 11118 13932
rect 11149 13923 11207 13929
rect 11149 13920 11161 13923
rect 11112 13892 11161 13920
rect 11112 13880 11118 13892
rect 11149 13889 11161 13892
rect 11195 13920 11207 13923
rect 11330 13920 11336 13932
rect 11195 13892 11336 13920
rect 11195 13889 11207 13892
rect 11149 13883 11207 13889
rect 11330 13880 11336 13892
rect 11388 13880 11394 13932
rect 11716 13920 11744 13960
rect 12618 13948 12624 13960
rect 12676 13948 12682 14000
rect 16117 13991 16175 13997
rect 16117 13957 16129 13991
rect 16163 13988 16175 13991
rect 16482 13988 16488 14000
rect 16163 13960 16488 13988
rect 16163 13957 16175 13960
rect 16117 13951 16175 13957
rect 16482 13948 16488 13960
rect 16540 13948 16546 14000
rect 24762 13988 24768 14000
rect 24723 13960 24768 13988
rect 24762 13948 24768 13960
rect 24820 13948 24826 14000
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11716 13892 11805 13920
rect 11793 13889 11805 13892
rect 11839 13889 11851 13923
rect 11793 13883 11851 13889
rect 12526 13880 12532 13932
rect 12584 13920 12590 13932
rect 12584 13892 13216 13920
rect 12584 13880 12590 13892
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 2038 13852 2044 13864
rect 1443 13824 2044 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 2130 13812 2136 13864
rect 2188 13852 2194 13864
rect 4522 13861 4528 13864
rect 2501 13855 2559 13861
rect 2501 13852 2513 13855
rect 2188 13824 2513 13852
rect 2188 13812 2194 13824
rect 2501 13821 2513 13824
rect 2547 13852 2559 13855
rect 2961 13855 3019 13861
rect 2961 13852 2973 13855
rect 2547 13824 2973 13852
rect 2547 13821 2559 13824
rect 2501 13815 2559 13821
rect 2961 13821 2973 13824
rect 3007 13821 3019 13855
rect 4505 13855 4528 13861
rect 4505 13852 4517 13855
rect 2961 13815 3019 13821
rect 3620 13824 4517 13852
rect 3620 13728 3648 13824
rect 4505 13821 4517 13824
rect 4580 13852 4586 13864
rect 5534 13852 5540 13864
rect 4580 13824 5540 13852
rect 4505 13815 4528 13821
rect 4522 13812 4528 13815
rect 4580 13812 4586 13824
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 6273 13855 6331 13861
rect 6273 13821 6285 13855
rect 6319 13852 6331 13855
rect 7098 13852 7104 13864
rect 6319 13824 7104 13852
rect 6319 13821 6331 13824
rect 6273 13815 6331 13821
rect 7098 13812 7104 13824
rect 7156 13852 7162 13864
rect 7193 13855 7251 13861
rect 7193 13852 7205 13855
rect 7156 13824 7205 13852
rect 7156 13812 7162 13824
rect 7193 13821 7205 13824
rect 7239 13821 7251 13855
rect 7193 13815 7251 13821
rect 7282 13812 7288 13864
rect 7340 13852 7346 13864
rect 7449 13855 7507 13861
rect 7449 13852 7461 13855
rect 7340 13824 7461 13852
rect 7340 13812 7346 13824
rect 7449 13821 7461 13824
rect 7495 13821 7507 13855
rect 9950 13852 9956 13864
rect 7449 13815 7507 13821
rect 8220 13824 9956 13852
rect 8110 13744 8116 13796
rect 8168 13784 8174 13796
rect 8220 13784 8248 13824
rect 9950 13812 9956 13824
rect 10008 13852 10014 13864
rect 10045 13855 10103 13861
rect 10045 13852 10057 13855
rect 10008 13824 10057 13852
rect 10008 13812 10014 13824
rect 10045 13821 10057 13824
rect 10091 13821 10103 13855
rect 11974 13852 11980 13864
rect 10045 13815 10103 13821
rect 10980 13824 11980 13852
rect 8168 13756 8248 13784
rect 10873 13787 10931 13793
rect 8168 13744 8174 13756
rect 10873 13753 10885 13787
rect 10919 13784 10931 13787
rect 10980 13784 11008 13824
rect 11974 13812 11980 13824
rect 12032 13812 12038 13864
rect 12802 13812 12808 13864
rect 12860 13852 12866 13864
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 12860 13824 13093 13852
rect 12860 13812 12866 13824
rect 13081 13821 13093 13824
rect 13127 13821 13139 13855
rect 13188 13852 13216 13892
rect 16390 13880 16396 13932
rect 16448 13920 16454 13932
rect 16666 13920 16672 13932
rect 16448 13892 16672 13920
rect 16448 13880 16454 13892
rect 16666 13880 16672 13892
rect 16724 13880 16730 13932
rect 18598 13920 18604 13932
rect 18559 13892 18604 13920
rect 18598 13880 18604 13892
rect 18656 13920 18662 13932
rect 19061 13923 19119 13929
rect 19061 13920 19073 13923
rect 18656 13892 19073 13920
rect 18656 13880 18662 13892
rect 19061 13889 19073 13892
rect 19107 13889 19119 13923
rect 19061 13883 19119 13889
rect 13354 13861 13360 13864
rect 13348 13852 13360 13861
rect 13188 13824 13360 13852
rect 13081 13815 13139 13821
rect 13348 13815 13360 13824
rect 13412 13852 13418 13864
rect 13412 13824 13768 13852
rect 13354 13812 13360 13815
rect 13412 13812 13418 13824
rect 10919 13756 11008 13784
rect 13740 13784 13768 13824
rect 15194 13812 15200 13864
rect 15252 13852 15258 13864
rect 16577 13855 16635 13861
rect 16577 13852 16589 13855
rect 15252 13824 16589 13852
rect 15252 13812 15258 13824
rect 16577 13821 16589 13824
rect 16623 13821 16635 13855
rect 16577 13815 16635 13821
rect 17218 13812 17224 13864
rect 17276 13852 17282 13864
rect 17589 13855 17647 13861
rect 17589 13852 17601 13855
rect 17276 13824 17601 13852
rect 17276 13812 17282 13824
rect 17589 13821 17601 13824
rect 17635 13852 17647 13855
rect 18509 13855 18567 13861
rect 17635 13824 17908 13852
rect 17635 13821 17647 13824
rect 17589 13815 17647 13821
rect 14642 13784 14648 13796
rect 13740 13756 14648 13784
rect 10919 13753 10931 13756
rect 10873 13747 10931 13753
rect 14642 13744 14648 13756
rect 14700 13744 14706 13796
rect 15930 13744 15936 13796
rect 15988 13784 15994 13796
rect 16485 13787 16543 13793
rect 16485 13784 16497 13787
rect 15988 13756 16497 13784
rect 15988 13744 15994 13756
rect 16485 13753 16497 13756
rect 16531 13784 16543 13787
rect 16758 13784 16764 13796
rect 16531 13756 16764 13784
rect 16531 13753 16543 13756
rect 16485 13747 16543 13753
rect 16758 13744 16764 13756
rect 16816 13744 16822 13796
rect 17880 13784 17908 13824
rect 18509 13821 18521 13855
rect 18555 13852 18567 13855
rect 19242 13852 19248 13864
rect 18555 13824 19248 13852
rect 18555 13821 18567 13824
rect 18509 13815 18567 13821
rect 19242 13812 19248 13824
rect 19300 13812 19306 13864
rect 20162 13852 20168 13864
rect 20123 13824 20168 13852
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 20993 13855 21051 13861
rect 20993 13821 21005 13855
rect 21039 13852 21051 13855
rect 21634 13852 21640 13864
rect 21039 13824 21640 13852
rect 21039 13821 21051 13824
rect 20993 13815 21051 13821
rect 21634 13812 21640 13824
rect 21692 13852 21698 13864
rect 21821 13855 21879 13861
rect 21821 13852 21833 13855
rect 21692 13824 21833 13852
rect 21692 13812 21698 13824
rect 21821 13821 21833 13824
rect 21867 13821 21879 13855
rect 21821 13815 21879 13821
rect 22557 13855 22615 13861
rect 22557 13821 22569 13855
rect 22603 13852 22615 13855
rect 23014 13852 23020 13864
rect 22603 13824 23020 13852
rect 22603 13821 22615 13824
rect 22557 13815 22615 13821
rect 23014 13812 23020 13824
rect 23072 13812 23078 13864
rect 23566 13812 23572 13864
rect 23624 13852 23630 13864
rect 23845 13855 23903 13861
rect 23845 13852 23857 13855
rect 23624 13824 23857 13852
rect 23624 13812 23630 13824
rect 23845 13821 23857 13824
rect 23891 13821 23903 13855
rect 24578 13852 24584 13864
rect 24539 13824 24584 13852
rect 23845 13815 23903 13821
rect 24578 13812 24584 13824
rect 24636 13852 24642 13864
rect 25133 13855 25191 13861
rect 25133 13852 25145 13855
rect 24636 13824 25145 13852
rect 24636 13812 24642 13824
rect 25133 13821 25145 13824
rect 25179 13821 25191 13855
rect 25133 13815 25191 13821
rect 19613 13787 19671 13793
rect 19613 13784 19625 13787
rect 17880 13756 19625 13784
rect 19613 13753 19625 13756
rect 19659 13753 19671 13787
rect 19613 13747 19671 13753
rect 2682 13716 2688 13728
rect 2643 13688 2688 13716
rect 2682 13676 2688 13688
rect 2740 13676 2746 13728
rect 3421 13719 3479 13725
rect 3421 13685 3433 13719
rect 3467 13716 3479 13719
rect 3602 13716 3608 13728
rect 3467 13688 3608 13716
rect 3467 13685 3479 13688
rect 3421 13679 3479 13685
rect 3602 13676 3608 13688
rect 3660 13676 3666 13728
rect 8570 13716 8576 13728
rect 8531 13688 8576 13716
rect 8570 13676 8576 13688
rect 8628 13676 8634 13728
rect 14274 13676 14280 13728
rect 14332 13716 14338 13728
rect 14461 13719 14519 13725
rect 14461 13716 14473 13719
rect 14332 13688 14473 13716
rect 14332 13676 14338 13688
rect 14461 13685 14473 13688
rect 14507 13685 14519 13719
rect 18414 13716 18420 13728
rect 18375 13688 18420 13716
rect 14461 13679 14519 13685
rect 18414 13676 18420 13688
rect 18472 13676 18478 13728
rect 20622 13676 20628 13728
rect 20680 13716 20686 13728
rect 21453 13719 21511 13725
rect 21453 13716 21465 13719
rect 20680 13688 21465 13716
rect 20680 13676 20686 13688
rect 21453 13685 21465 13688
rect 21499 13685 21511 13719
rect 21453 13679 21511 13685
rect 22646 13676 22652 13728
rect 22704 13716 22710 13728
rect 22741 13719 22799 13725
rect 22741 13716 22753 13719
rect 22704 13688 22753 13716
rect 22704 13676 22710 13688
rect 22741 13685 22753 13688
rect 22787 13685 22799 13719
rect 24394 13716 24400 13728
rect 24355 13688 24400 13716
rect 22741 13679 22799 13685
rect 24394 13676 24400 13688
rect 24452 13716 24458 13728
rect 24670 13716 24676 13728
rect 24452 13688 24676 13716
rect 24452 13676 24458 13688
rect 24670 13676 24676 13688
rect 24728 13676 24734 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1394 13472 1400 13524
rect 1452 13512 1458 13524
rect 2041 13515 2099 13521
rect 2041 13512 2053 13515
rect 1452 13484 2053 13512
rect 1452 13472 1458 13484
rect 2041 13481 2053 13484
rect 2087 13512 2099 13515
rect 2682 13512 2688 13524
rect 2087 13484 2688 13512
rect 2087 13481 2099 13484
rect 2041 13475 2099 13481
rect 2682 13472 2688 13484
rect 2740 13472 2746 13524
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 5629 13515 5687 13521
rect 5629 13512 5641 13515
rect 5592 13484 5641 13512
rect 5592 13472 5598 13484
rect 5629 13481 5641 13484
rect 5675 13481 5687 13515
rect 7282 13512 7288 13524
rect 7243 13484 7288 13512
rect 5629 13475 5687 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 7558 13512 7564 13524
rect 7519 13484 7564 13512
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 9122 13472 9128 13524
rect 9180 13512 9186 13524
rect 10137 13515 10195 13521
rect 10137 13512 10149 13515
rect 9180 13484 10149 13512
rect 9180 13472 9186 13484
rect 10137 13481 10149 13484
rect 10183 13481 10195 13515
rect 10137 13475 10195 13481
rect 10781 13515 10839 13521
rect 10781 13481 10793 13515
rect 10827 13512 10839 13515
rect 10962 13512 10968 13524
rect 10827 13484 10968 13512
rect 10827 13481 10839 13484
rect 10781 13475 10839 13481
rect 6638 13404 6644 13456
rect 6696 13444 6702 13456
rect 7742 13444 7748 13456
rect 6696 13416 7748 13444
rect 6696 13404 6702 13416
rect 7742 13404 7748 13416
rect 7800 13444 7806 13456
rect 8021 13447 8079 13453
rect 8021 13444 8033 13447
rect 7800 13416 8033 13444
rect 7800 13404 7806 13416
rect 8021 13413 8033 13416
rect 8067 13413 8079 13447
rect 10152 13444 10180 13475
rect 10962 13472 10968 13484
rect 11020 13472 11026 13524
rect 12250 13512 12256 13524
rect 12211 13484 12256 13512
rect 12250 13472 12256 13484
rect 12308 13472 12314 13524
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 13081 13515 13139 13521
rect 13081 13512 13093 13515
rect 12860 13484 13093 13512
rect 12860 13472 12866 13484
rect 13081 13481 13093 13484
rect 13127 13481 13139 13515
rect 13081 13475 13139 13481
rect 13541 13515 13599 13521
rect 13541 13481 13553 13515
rect 13587 13481 13599 13515
rect 13541 13475 13599 13481
rect 10152 13416 11008 13444
rect 8021 13407 8079 13413
rect 10980 13388 11008 13416
rect 11146 13404 11152 13456
rect 11204 13444 11210 13456
rect 12345 13447 12403 13453
rect 12345 13444 12357 13447
rect 11204 13416 12357 13444
rect 11204 13404 11210 13416
rect 12345 13413 12357 13416
rect 12391 13413 12403 13447
rect 12345 13407 12403 13413
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 2038 13376 2044 13388
rect 1443 13348 2044 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 2038 13336 2044 13348
rect 2096 13336 2102 13388
rect 2498 13376 2504 13388
rect 2411 13348 2504 13376
rect 2498 13336 2504 13348
rect 2556 13376 2562 13388
rect 3421 13379 3479 13385
rect 3421 13376 3433 13379
rect 2556 13348 3433 13376
rect 2556 13336 2562 13348
rect 3421 13345 3433 13348
rect 3467 13345 3479 13379
rect 3421 13339 3479 13345
rect 4154 13336 4160 13388
rect 4212 13376 4218 13388
rect 4249 13379 4307 13385
rect 4249 13376 4261 13379
rect 4212 13348 4261 13376
rect 4212 13336 4218 13348
rect 4249 13345 4261 13348
rect 4295 13345 4307 13379
rect 4249 13339 4307 13345
rect 4516 13379 4574 13385
rect 4516 13345 4528 13379
rect 4562 13376 4574 13379
rect 5074 13376 5080 13388
rect 4562 13348 5080 13376
rect 4562 13345 4574 13348
rect 4516 13339 4574 13345
rect 5074 13336 5080 13348
rect 5132 13336 5138 13388
rect 6917 13379 6975 13385
rect 6917 13345 6929 13379
rect 6963 13376 6975 13379
rect 7558 13376 7564 13388
rect 6963 13348 7564 13376
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 7558 13336 7564 13348
rect 7616 13376 7622 13388
rect 7929 13379 7987 13385
rect 7929 13376 7941 13379
rect 7616 13348 7941 13376
rect 7616 13336 7622 13348
rect 7929 13345 7941 13348
rect 7975 13345 7987 13379
rect 7929 13339 7987 13345
rect 9306 13336 9312 13388
rect 9364 13376 9370 13388
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 9364 13348 10057 13376
rect 9364 13336 9370 13348
rect 10045 13345 10057 13348
rect 10091 13376 10103 13379
rect 10686 13376 10692 13388
rect 10091 13348 10692 13376
rect 10091 13345 10103 13348
rect 10045 13339 10103 13345
rect 10686 13336 10692 13348
rect 10744 13336 10750 13388
rect 10962 13336 10968 13388
rect 11020 13336 11026 13388
rect 12360 13376 12388 13407
rect 12618 13376 12624 13388
rect 12360 13348 12624 13376
rect 12618 13336 12624 13348
rect 12676 13336 12682 13388
rect 13096 13376 13124 13475
rect 13556 13444 13584 13475
rect 14182 13472 14188 13524
rect 14240 13512 14246 13524
rect 14366 13512 14372 13524
rect 14240 13484 14372 13512
rect 14240 13472 14246 13484
rect 14366 13472 14372 13484
rect 14424 13512 14430 13524
rect 14553 13515 14611 13521
rect 14553 13512 14565 13515
rect 14424 13484 14565 13512
rect 14424 13472 14430 13484
rect 14553 13481 14565 13484
rect 14599 13481 14611 13515
rect 15102 13512 15108 13524
rect 15063 13484 15108 13512
rect 14553 13475 14611 13481
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 15838 13512 15844 13524
rect 15799 13484 15844 13512
rect 15838 13472 15844 13484
rect 15896 13472 15902 13524
rect 16666 13472 16672 13524
rect 16724 13512 16730 13524
rect 17310 13512 17316 13524
rect 16724 13484 17316 13512
rect 16724 13472 16730 13484
rect 17310 13472 17316 13484
rect 17368 13512 17374 13524
rect 17405 13515 17463 13521
rect 17405 13512 17417 13515
rect 17368 13484 17417 13512
rect 17368 13472 17374 13484
rect 17405 13481 17417 13484
rect 17451 13481 17463 13515
rect 17405 13475 17463 13481
rect 23753 13515 23811 13521
rect 23753 13481 23765 13515
rect 23799 13512 23811 13515
rect 24394 13512 24400 13524
rect 23799 13484 24400 13512
rect 23799 13481 23811 13484
rect 23753 13475 23811 13481
rect 24394 13472 24400 13484
rect 24452 13472 24458 13524
rect 24762 13512 24768 13524
rect 24723 13484 24768 13512
rect 24762 13472 24768 13484
rect 24820 13472 24826 13524
rect 15120 13444 15148 13472
rect 13556 13416 15148 13444
rect 19426 13404 19432 13456
rect 19484 13444 19490 13456
rect 19794 13444 19800 13456
rect 19484 13416 19800 13444
rect 19484 13404 19490 13416
rect 19794 13404 19800 13416
rect 19852 13404 19858 13456
rect 13630 13376 13636 13388
rect 13096 13348 13636 13376
rect 13630 13336 13636 13348
rect 13688 13336 13694 13388
rect 13906 13376 13912 13388
rect 13867 13348 13912 13376
rect 13906 13336 13912 13348
rect 13964 13336 13970 13388
rect 14001 13379 14059 13385
rect 14001 13345 14013 13379
rect 14047 13376 14059 13379
rect 14458 13376 14464 13388
rect 14047 13348 14464 13376
rect 14047 13345 14059 13348
rect 14001 13339 14059 13345
rect 2866 13308 2872 13320
rect 1504 13280 2872 13308
rect 1504 13172 1532 13280
rect 2866 13268 2872 13280
rect 2924 13268 2930 13320
rect 8110 13308 8116 13320
rect 8071 13280 8116 13308
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 12526 13308 12532 13320
rect 10284 13280 10329 13308
rect 12487 13280 12532 13308
rect 10284 13268 10290 13280
rect 12526 13268 12532 13280
rect 12584 13268 12590 13320
rect 2409 13243 2467 13249
rect 2409 13209 2421 13243
rect 2455 13240 2467 13243
rect 2590 13240 2596 13252
rect 2455 13212 2596 13240
rect 2455 13209 2467 13212
rect 2409 13203 2467 13209
rect 2590 13200 2596 13212
rect 2648 13200 2654 13252
rect 11885 13243 11943 13249
rect 11885 13209 11897 13243
rect 11931 13240 11943 13243
rect 14016 13240 14044 13339
rect 14458 13336 14464 13348
rect 14516 13336 14522 13388
rect 16281 13379 16339 13385
rect 16281 13376 16293 13379
rect 15672 13348 16293 13376
rect 14182 13308 14188 13320
rect 14143 13280 14188 13308
rect 14182 13268 14188 13280
rect 14240 13308 14246 13320
rect 15672 13308 15700 13348
rect 16281 13345 16293 13348
rect 16327 13376 16339 13379
rect 16574 13376 16580 13388
rect 16327 13348 16580 13376
rect 16327 13345 16339 13348
rect 16281 13339 16339 13345
rect 16574 13336 16580 13348
rect 16632 13336 16638 13388
rect 18782 13336 18788 13388
rect 18840 13376 18846 13388
rect 18877 13379 18935 13385
rect 18877 13376 18889 13379
rect 18840 13348 18889 13376
rect 18840 13336 18846 13348
rect 18877 13345 18889 13348
rect 18923 13345 18935 13379
rect 18877 13339 18935 13345
rect 23474 13336 23480 13388
rect 23532 13376 23538 13388
rect 23569 13379 23627 13385
rect 23569 13376 23581 13379
rect 23532 13348 23581 13376
rect 23532 13336 23538 13348
rect 23569 13345 23581 13348
rect 23615 13345 23627 13379
rect 23569 13339 23627 13345
rect 24210 13336 24216 13388
rect 24268 13376 24274 13388
rect 24581 13379 24639 13385
rect 24581 13376 24593 13379
rect 24268 13348 24593 13376
rect 24268 13336 24274 13348
rect 24581 13345 24593 13348
rect 24627 13345 24639 13379
rect 24581 13339 24639 13345
rect 16022 13308 16028 13320
rect 14240 13280 15700 13308
rect 15983 13280 16028 13308
rect 14240 13268 14246 13280
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 18966 13308 18972 13320
rect 18927 13280 18972 13308
rect 18966 13268 18972 13280
rect 19024 13268 19030 13320
rect 19058 13268 19064 13320
rect 19116 13308 19122 13320
rect 19116 13280 19161 13308
rect 19116 13268 19122 13280
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 20070 13308 20076 13320
rect 19484 13280 20076 13308
rect 19484 13268 19490 13280
rect 20070 13268 20076 13280
rect 20128 13268 20134 13320
rect 20901 13311 20959 13317
rect 20901 13277 20913 13311
rect 20947 13308 20959 13311
rect 21082 13308 21088 13320
rect 20947 13280 21088 13308
rect 20947 13277 20959 13280
rect 20901 13271 20959 13277
rect 21082 13268 21088 13280
rect 21140 13268 21146 13320
rect 22557 13311 22615 13317
rect 22557 13277 22569 13311
rect 22603 13308 22615 13311
rect 23106 13308 23112 13320
rect 22603 13280 23112 13308
rect 22603 13277 22615 13280
rect 22557 13271 22615 13277
rect 23106 13268 23112 13280
rect 23164 13268 23170 13320
rect 23842 13268 23848 13320
rect 23900 13308 23906 13320
rect 24762 13308 24768 13320
rect 23900 13280 24768 13308
rect 23900 13268 23906 13280
rect 24762 13268 24768 13280
rect 24820 13268 24826 13320
rect 11931 13212 14044 13240
rect 11931 13209 11943 13212
rect 11885 13203 11943 13209
rect 14274 13200 14280 13252
rect 14332 13240 14338 13252
rect 14550 13240 14556 13252
rect 14332 13212 14556 13240
rect 14332 13200 14338 13212
rect 14550 13200 14556 13212
rect 14608 13200 14614 13252
rect 20346 13240 20352 13252
rect 19628 13212 20352 13240
rect 19628 13184 19656 13212
rect 20346 13200 20352 13212
rect 20404 13200 20410 13252
rect 1581 13175 1639 13181
rect 1581 13172 1593 13175
rect 1504 13144 1593 13172
rect 1581 13141 1593 13144
rect 1627 13141 1639 13175
rect 1581 13135 1639 13141
rect 1670 13132 1676 13184
rect 1728 13172 1734 13184
rect 2685 13175 2743 13181
rect 2685 13172 2697 13175
rect 1728 13144 2697 13172
rect 1728 13132 1734 13144
rect 2685 13141 2697 13144
rect 2731 13141 2743 13175
rect 2685 13135 2743 13141
rect 2774 13132 2780 13184
rect 2832 13172 2838 13184
rect 3053 13175 3111 13181
rect 3053 13172 3065 13175
rect 2832 13144 3065 13172
rect 2832 13132 2838 13144
rect 3053 13141 3065 13144
rect 3099 13141 3111 13175
rect 3878 13172 3884 13184
rect 3839 13144 3884 13172
rect 3053 13135 3111 13141
rect 3878 13132 3884 13144
rect 3936 13132 3942 13184
rect 8570 13172 8576 13184
rect 8531 13144 8576 13172
rect 8570 13132 8576 13144
rect 8628 13132 8634 13184
rect 9398 13172 9404 13184
rect 9359 13144 9404 13172
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 9677 13175 9735 13181
rect 9677 13141 9689 13175
rect 9723 13172 9735 13175
rect 9766 13172 9772 13184
rect 9723 13144 9772 13172
rect 9723 13141 9735 13144
rect 9677 13135 9735 13141
rect 9766 13132 9772 13144
rect 9824 13132 9830 13184
rect 11330 13172 11336 13184
rect 11291 13144 11336 13172
rect 11330 13132 11336 13144
rect 11388 13132 11394 13184
rect 11793 13175 11851 13181
rect 11793 13141 11805 13175
rect 11839 13172 11851 13175
rect 12802 13172 12808 13184
rect 11839 13144 12808 13172
rect 11839 13141 11851 13144
rect 11793 13135 11851 13141
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 15562 13172 15568 13184
rect 15523 13144 15568 13172
rect 15562 13132 15568 13144
rect 15620 13132 15626 13184
rect 18141 13175 18199 13181
rect 18141 13141 18153 13175
rect 18187 13172 18199 13175
rect 18322 13172 18328 13184
rect 18187 13144 18328 13172
rect 18187 13141 18199 13144
rect 18141 13135 18199 13141
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 18506 13172 18512 13184
rect 18467 13144 18512 13172
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 19610 13172 19616 13184
rect 19571 13144 19616 13172
rect 19610 13132 19616 13144
rect 19668 13132 19674 13184
rect 20070 13172 20076 13184
rect 20031 13144 20076 13172
rect 20070 13132 20076 13144
rect 20128 13132 20134 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1486 12928 1492 12980
rect 1544 12968 1550 12980
rect 1581 12971 1639 12977
rect 1581 12968 1593 12971
rect 1544 12940 1593 12968
rect 1544 12928 1550 12940
rect 1581 12937 1593 12940
rect 1627 12937 1639 12971
rect 1581 12931 1639 12937
rect 1670 12928 1676 12980
rect 1728 12968 1734 12980
rect 1854 12968 1860 12980
rect 1728 12940 1860 12968
rect 1728 12928 1734 12940
rect 1854 12928 1860 12940
rect 1912 12928 1918 12980
rect 3050 12968 3056 12980
rect 3011 12940 3056 12968
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 6638 12968 6644 12980
rect 6599 12940 6644 12968
rect 6638 12928 6644 12940
rect 6696 12928 6702 12980
rect 7558 12928 7564 12980
rect 7616 12968 7622 12980
rect 8113 12971 8171 12977
rect 8113 12968 8125 12971
rect 7616 12940 8125 12968
rect 7616 12928 7622 12940
rect 8113 12937 8125 12940
rect 8159 12937 8171 12971
rect 9122 12968 9128 12980
rect 9083 12940 9128 12968
rect 8113 12931 8171 12937
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 9306 12928 9312 12980
rect 9364 12968 9370 12980
rect 9493 12971 9551 12977
rect 9493 12968 9505 12971
rect 9364 12940 9505 12968
rect 9364 12928 9370 12940
rect 9493 12937 9505 12940
rect 9539 12937 9551 12971
rect 11146 12968 11152 12980
rect 11107 12940 11152 12968
rect 9493 12931 9551 12937
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 11977 12971 12035 12977
rect 11977 12937 11989 12971
rect 12023 12968 12035 12971
rect 12250 12968 12256 12980
rect 12023 12940 12256 12968
rect 12023 12937 12035 12940
rect 11977 12931 12035 12937
rect 12250 12928 12256 12940
rect 12308 12928 12314 12980
rect 13633 12971 13691 12977
rect 13633 12937 13645 12971
rect 13679 12968 13691 12971
rect 13906 12968 13912 12980
rect 13679 12940 13912 12968
rect 13679 12937 13691 12940
rect 13633 12931 13691 12937
rect 13906 12928 13912 12940
rect 13964 12928 13970 12980
rect 14642 12968 14648 12980
rect 14603 12940 14648 12968
rect 14642 12928 14648 12940
rect 14700 12928 14706 12980
rect 15197 12971 15255 12977
rect 15197 12937 15209 12971
rect 15243 12968 15255 12971
rect 15930 12968 15936 12980
rect 15243 12940 15936 12968
rect 15243 12937 15255 12940
rect 15197 12931 15255 12937
rect 15930 12928 15936 12940
rect 15988 12928 15994 12980
rect 16022 12928 16028 12980
rect 16080 12968 16086 12980
rect 16209 12971 16267 12977
rect 16209 12968 16221 12971
rect 16080 12940 16221 12968
rect 16080 12928 16086 12940
rect 16209 12937 16221 12940
rect 16255 12937 16267 12971
rect 16574 12968 16580 12980
rect 16535 12940 16580 12968
rect 16209 12931 16267 12937
rect 16574 12928 16580 12940
rect 16632 12928 16638 12980
rect 16945 12971 17003 12977
rect 16945 12937 16957 12971
rect 16991 12968 17003 12971
rect 17770 12968 17776 12980
rect 16991 12940 17776 12968
rect 16991 12937 17003 12940
rect 16945 12931 17003 12937
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 19334 12928 19340 12980
rect 19392 12968 19398 12980
rect 19613 12971 19671 12977
rect 19613 12968 19625 12971
rect 19392 12940 19625 12968
rect 19392 12928 19398 12940
rect 19613 12937 19625 12940
rect 19659 12937 19671 12971
rect 20714 12968 20720 12980
rect 20675 12940 20720 12968
rect 19613 12931 19671 12937
rect 20714 12928 20720 12940
rect 20772 12928 20778 12980
rect 20898 12928 20904 12980
rect 20956 12968 20962 12980
rect 20993 12971 21051 12977
rect 20993 12968 21005 12971
rect 20956 12940 21005 12968
rect 20956 12928 20962 12940
rect 20993 12937 21005 12940
rect 21039 12937 21051 12971
rect 20993 12931 21051 12937
rect 23474 12928 23480 12980
rect 23532 12968 23538 12980
rect 23845 12971 23903 12977
rect 23845 12968 23857 12971
rect 23532 12940 23857 12968
rect 23532 12928 23538 12940
rect 23845 12937 23857 12940
rect 23891 12937 23903 12971
rect 23845 12931 23903 12937
rect 24765 12971 24823 12977
rect 24765 12937 24777 12971
rect 24811 12968 24823 12971
rect 24946 12968 24952 12980
rect 24811 12940 24952 12968
rect 24811 12937 24823 12940
rect 24765 12931 24823 12937
rect 24946 12928 24952 12940
rect 25004 12928 25010 12980
rect 4617 12903 4675 12909
rect 4617 12900 4629 12903
rect 3528 12872 4629 12900
rect 2314 12792 2320 12844
rect 2372 12832 2378 12844
rect 2590 12832 2596 12844
rect 2372 12804 2596 12832
rect 2372 12792 2378 12804
rect 2590 12792 2596 12804
rect 2648 12792 2654 12844
rect 3142 12792 3148 12844
rect 3200 12832 3206 12844
rect 3528 12841 3556 12872
rect 4617 12869 4629 12872
rect 4663 12869 4675 12903
rect 4617 12863 4675 12869
rect 3513 12835 3571 12841
rect 3513 12832 3525 12835
rect 3200 12804 3525 12832
rect 3200 12792 3206 12804
rect 3513 12801 3525 12804
rect 3559 12801 3571 12835
rect 3513 12795 3571 12801
rect 3602 12792 3608 12844
rect 3660 12832 3666 12844
rect 3660 12804 3705 12832
rect 3660 12792 3666 12804
rect 5074 12792 5080 12844
rect 5132 12832 5138 12844
rect 5169 12835 5227 12841
rect 5169 12832 5181 12835
rect 5132 12804 5181 12832
rect 5132 12792 5138 12804
rect 5169 12801 5181 12804
rect 5215 12832 5227 12835
rect 5629 12835 5687 12841
rect 5629 12832 5641 12835
rect 5215 12804 5641 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 5629 12801 5641 12804
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 8570 12792 8576 12844
rect 8628 12832 8634 12844
rect 8665 12835 8723 12841
rect 8665 12832 8677 12835
rect 8628 12804 8677 12832
rect 8628 12792 8634 12804
rect 8665 12801 8677 12804
rect 8711 12801 8723 12835
rect 10226 12832 10232 12844
rect 10187 12804 10232 12832
rect 8665 12795 8723 12801
rect 10226 12792 10232 12804
rect 10284 12792 10290 12844
rect 14277 12835 14335 12841
rect 14277 12801 14289 12835
rect 14323 12832 14335 12835
rect 14660 12832 14688 12928
rect 17954 12900 17960 12912
rect 16776 12872 17960 12900
rect 14323 12804 14688 12832
rect 14323 12801 14335 12804
rect 14277 12795 14335 12801
rect 15562 12792 15568 12844
rect 15620 12832 15626 12844
rect 15749 12835 15807 12841
rect 15749 12832 15761 12835
rect 15620 12804 15761 12832
rect 15620 12792 15626 12804
rect 15749 12801 15761 12804
rect 15795 12832 15807 12835
rect 15930 12832 15936 12844
rect 15795 12804 15936 12832
rect 15795 12801 15807 12804
rect 15749 12795 15807 12801
rect 15930 12792 15936 12804
rect 15988 12792 15994 12844
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 2038 12764 2044 12776
rect 1999 12736 2044 12764
rect 2038 12724 2044 12736
rect 2096 12724 2102 12776
rect 3418 12764 3424 12776
rect 3379 12736 3424 12764
rect 3418 12724 3424 12736
rect 3476 12764 3482 12776
rect 4154 12764 4160 12776
rect 3476 12736 4160 12764
rect 3476 12724 3482 12736
rect 4154 12724 4160 12736
rect 4212 12724 4218 12776
rect 7101 12767 7159 12773
rect 7101 12733 7113 12767
rect 7147 12764 7159 12767
rect 7374 12764 7380 12776
rect 7147 12736 7380 12764
rect 7147 12733 7159 12736
rect 7101 12727 7159 12733
rect 7374 12724 7380 12736
rect 7432 12724 7438 12776
rect 7653 12767 7711 12773
rect 7653 12733 7665 12767
rect 7699 12764 7711 12767
rect 8202 12764 8208 12776
rect 7699 12736 8208 12764
rect 7699 12733 7711 12736
rect 7653 12727 7711 12733
rect 8202 12724 8208 12736
rect 8260 12764 8266 12776
rect 8481 12767 8539 12773
rect 8481 12764 8493 12767
rect 8260 12736 8493 12764
rect 8260 12724 8266 12736
rect 8481 12733 8493 12736
rect 8527 12733 8539 12767
rect 11330 12764 11336 12776
rect 11291 12736 11336 12764
rect 8481 12727 8539 12733
rect 11330 12724 11336 12736
rect 11388 12724 11394 12776
rect 12621 12767 12679 12773
rect 12621 12733 12633 12767
rect 12667 12764 12679 12767
rect 12802 12764 12808 12776
rect 12667 12736 12808 12764
rect 12667 12733 12679 12736
rect 12621 12727 12679 12733
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 13354 12724 13360 12776
rect 13412 12764 13418 12776
rect 13541 12767 13599 12773
rect 13541 12764 13553 12767
rect 13412 12736 13553 12764
rect 13412 12724 13418 12736
rect 13541 12733 13553 12736
rect 13587 12764 13599 12767
rect 13998 12764 14004 12776
rect 13587 12736 14004 12764
rect 13587 12733 13599 12736
rect 13541 12727 13599 12733
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 16574 12724 16580 12776
rect 16632 12764 16638 12776
rect 16776 12773 16804 12872
rect 17954 12860 17960 12872
rect 18012 12860 18018 12912
rect 22741 12903 22799 12909
rect 22741 12869 22753 12903
rect 22787 12900 22799 12903
rect 24210 12900 24216 12912
rect 22787 12872 24216 12900
rect 22787 12869 22799 12872
rect 22741 12863 22799 12869
rect 24210 12860 24216 12872
rect 24268 12900 24274 12912
rect 24397 12903 24455 12909
rect 24397 12900 24409 12903
rect 24268 12872 24409 12900
rect 24268 12860 24274 12872
rect 24397 12869 24409 12872
rect 24443 12869 24455 12903
rect 24397 12863 24455 12869
rect 17126 12792 17132 12844
rect 17184 12832 17190 12844
rect 17497 12835 17555 12841
rect 17497 12832 17509 12835
rect 17184 12804 17509 12832
rect 17184 12792 17190 12804
rect 17497 12801 17509 12804
rect 17543 12832 17555 12835
rect 18601 12835 18659 12841
rect 18601 12832 18613 12835
rect 17543 12804 18613 12832
rect 17543 12801 17555 12804
rect 17497 12795 17555 12801
rect 18601 12801 18613 12804
rect 18647 12801 18659 12835
rect 18601 12795 18659 12801
rect 20070 12792 20076 12844
rect 20128 12832 20134 12844
rect 20165 12835 20223 12841
rect 20165 12832 20177 12835
rect 20128 12804 20177 12832
rect 20128 12792 20134 12804
rect 20165 12801 20177 12804
rect 20211 12801 20223 12835
rect 20165 12795 20223 12801
rect 16761 12767 16819 12773
rect 16761 12764 16773 12767
rect 16632 12736 16773 12764
rect 16632 12724 16638 12736
rect 16761 12733 16773 12736
rect 16807 12733 16819 12767
rect 18509 12767 18567 12773
rect 18509 12764 18521 12767
rect 16761 12727 16819 12733
rect 17788 12736 18521 12764
rect 2317 12699 2375 12705
rect 2317 12696 2329 12699
rect 1412 12668 2329 12696
rect 1412 12640 1440 12668
rect 2317 12665 2329 12668
rect 2363 12665 2375 12699
rect 2317 12659 2375 12665
rect 2961 12699 3019 12705
rect 2961 12665 2973 12699
rect 3007 12696 3019 12699
rect 3602 12696 3608 12708
rect 3007 12668 3608 12696
rect 3007 12665 3019 12668
rect 2961 12659 3019 12665
rect 3602 12656 3608 12668
rect 3660 12656 3666 12708
rect 4525 12699 4583 12705
rect 4525 12665 4537 12699
rect 4571 12696 4583 12699
rect 4982 12696 4988 12708
rect 4571 12668 4988 12696
rect 4571 12665 4583 12668
rect 4525 12659 4583 12665
rect 4982 12656 4988 12668
rect 5040 12656 5046 12708
rect 5077 12699 5135 12705
rect 5077 12665 5089 12699
rect 5123 12696 5135 12699
rect 7466 12696 7472 12708
rect 5123 12668 7472 12696
rect 5123 12665 5135 12668
rect 5077 12659 5135 12665
rect 1394 12588 1400 12640
rect 1452 12588 1458 12640
rect 2038 12588 2044 12640
rect 2096 12628 2102 12640
rect 2222 12628 2228 12640
rect 2096 12600 2228 12628
rect 2096 12588 2102 12600
rect 2222 12588 2228 12600
rect 2280 12588 2286 12640
rect 3326 12588 3332 12640
rect 3384 12628 3390 12640
rect 4157 12631 4215 12637
rect 4157 12628 4169 12631
rect 3384 12600 4169 12628
rect 3384 12588 3390 12600
rect 4157 12597 4169 12600
rect 4203 12628 4215 12631
rect 5092 12628 5120 12659
rect 7466 12656 7472 12668
rect 7524 12656 7530 12708
rect 9858 12656 9864 12708
rect 9916 12696 9922 12708
rect 9916 12668 10180 12696
rect 9916 12656 9922 12668
rect 4203 12600 5120 12628
rect 7285 12631 7343 12637
rect 4203 12597 4215 12600
rect 4157 12591 4215 12597
rect 7285 12597 7297 12631
rect 7331 12628 7343 12631
rect 7926 12628 7932 12640
rect 7331 12600 7932 12628
rect 7331 12597 7343 12600
rect 7285 12591 7343 12597
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 8021 12631 8079 12637
rect 8021 12597 8033 12631
rect 8067 12628 8079 12631
rect 8570 12628 8576 12640
rect 8067 12600 8576 12628
rect 8067 12597 8079 12600
rect 8021 12591 8079 12597
rect 8570 12588 8576 12600
rect 8628 12588 8634 12640
rect 9674 12628 9680 12640
rect 9635 12600 9680 12628
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 10042 12628 10048 12640
rect 10003 12600 10048 12628
rect 10042 12588 10048 12600
rect 10100 12588 10106 12640
rect 10152 12637 10180 12668
rect 11238 12656 11244 12708
rect 11296 12696 11302 12708
rect 15105 12699 15163 12705
rect 11296 12668 13216 12696
rect 11296 12656 11302 12668
rect 10137 12631 10195 12637
rect 10137 12597 10149 12631
rect 10183 12628 10195 12631
rect 10689 12631 10747 12637
rect 10689 12628 10701 12631
rect 10183 12600 10701 12628
rect 10183 12597 10195 12600
rect 10137 12591 10195 12597
rect 10689 12597 10701 12600
rect 10735 12597 10747 12631
rect 10689 12591 10747 12597
rect 11330 12588 11336 12640
rect 11388 12628 11394 12640
rect 11517 12631 11575 12637
rect 11517 12628 11529 12631
rect 11388 12600 11529 12628
rect 11388 12588 11394 12600
rect 11517 12597 11529 12600
rect 11563 12597 11575 12631
rect 11517 12591 11575 12597
rect 12526 12588 12532 12640
rect 12584 12628 12590 12640
rect 13188 12637 13216 12668
rect 15105 12665 15117 12699
rect 15151 12696 15163 12699
rect 15286 12696 15292 12708
rect 15151 12668 15292 12696
rect 15151 12665 15163 12668
rect 15105 12659 15163 12665
rect 15286 12656 15292 12668
rect 15344 12696 15350 12708
rect 15565 12699 15623 12705
rect 15565 12696 15577 12699
rect 15344 12668 15577 12696
rect 15344 12656 15350 12668
rect 15565 12665 15577 12668
rect 15611 12665 15623 12699
rect 15565 12659 15623 12665
rect 16666 12656 16672 12708
rect 16724 12696 16730 12708
rect 17788 12705 17816 12736
rect 18509 12733 18521 12736
rect 18555 12733 18567 12767
rect 19610 12764 19616 12776
rect 18509 12727 18567 12733
rect 19444 12736 19616 12764
rect 17773 12699 17831 12705
rect 17773 12696 17785 12699
rect 16724 12668 17785 12696
rect 16724 12656 16730 12668
rect 17773 12665 17785 12668
rect 17819 12665 17831 12699
rect 17773 12659 17831 12665
rect 18138 12656 18144 12708
rect 18196 12696 18202 12708
rect 19058 12696 19064 12708
rect 18196 12668 19064 12696
rect 18196 12656 18202 12668
rect 19058 12656 19064 12668
rect 19116 12656 19122 12708
rect 12805 12631 12863 12637
rect 12805 12628 12817 12631
rect 12584 12600 12817 12628
rect 12584 12588 12590 12600
rect 12805 12597 12817 12600
rect 12851 12597 12863 12631
rect 12805 12591 12863 12597
rect 13173 12631 13231 12637
rect 13173 12597 13185 12631
rect 13219 12628 13231 12631
rect 14093 12631 14151 12637
rect 14093 12628 14105 12631
rect 13219 12600 14105 12628
rect 13219 12597 13231 12600
rect 13173 12591 13231 12597
rect 14093 12597 14105 12600
rect 14139 12628 14151 12631
rect 15470 12628 15476 12640
rect 14139 12600 15476 12628
rect 14139 12597 14151 12600
rect 14093 12591 14151 12597
rect 15470 12588 15476 12600
rect 15528 12588 15534 12640
rect 15654 12628 15660 12640
rect 15615 12600 15660 12628
rect 15654 12588 15660 12600
rect 15712 12588 15718 12640
rect 18046 12628 18052 12640
rect 18007 12600 18052 12628
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 18322 12588 18328 12640
rect 18380 12628 18386 12640
rect 18417 12631 18475 12637
rect 18417 12628 18429 12631
rect 18380 12600 18429 12628
rect 18380 12588 18386 12600
rect 18417 12597 18429 12600
rect 18463 12628 18475 12631
rect 19242 12628 19248 12640
rect 18463 12600 19248 12628
rect 18463 12597 18475 12600
rect 18417 12591 18475 12597
rect 19242 12588 19248 12600
rect 19300 12588 19306 12640
rect 19444 12628 19472 12736
rect 19610 12724 19616 12736
rect 19668 12724 19674 12776
rect 22554 12764 22560 12776
rect 22515 12736 22560 12764
rect 22554 12724 22560 12736
rect 22612 12764 22618 12776
rect 23017 12767 23075 12773
rect 23017 12764 23029 12767
rect 22612 12736 23029 12764
rect 22612 12724 22618 12736
rect 23017 12733 23029 12736
rect 23063 12733 23075 12767
rect 23017 12727 23075 12733
rect 24118 12724 24124 12776
rect 24176 12764 24182 12776
rect 24581 12767 24639 12773
rect 24581 12764 24593 12767
rect 24176 12736 24593 12764
rect 24176 12724 24182 12736
rect 24581 12733 24593 12736
rect 24627 12764 24639 12767
rect 25133 12767 25191 12773
rect 25133 12764 25145 12767
rect 24627 12736 25145 12764
rect 24627 12733 24639 12736
rect 24581 12727 24639 12733
rect 25133 12733 25145 12736
rect 25179 12733 25191 12767
rect 25133 12727 25191 12733
rect 19521 12699 19579 12705
rect 19521 12665 19533 12699
rect 19567 12696 19579 12699
rect 19981 12699 20039 12705
rect 19981 12696 19993 12699
rect 19567 12668 19993 12696
rect 19567 12665 19579 12668
rect 19521 12659 19579 12665
rect 19981 12665 19993 12668
rect 20027 12696 20039 12699
rect 20346 12696 20352 12708
rect 20027 12668 20352 12696
rect 20027 12665 20039 12668
rect 19981 12659 20039 12665
rect 20346 12656 20352 12668
rect 20404 12656 20410 12708
rect 20073 12631 20131 12637
rect 20073 12628 20085 12631
rect 19444 12600 20085 12628
rect 20073 12597 20085 12600
rect 20119 12597 20131 12631
rect 21174 12628 21180 12640
rect 21135 12600 21180 12628
rect 20073 12591 20131 12597
rect 21174 12588 21180 12600
rect 21232 12588 21238 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1486 12384 1492 12436
rect 1544 12424 1550 12436
rect 1762 12424 1768 12436
rect 1544 12396 1768 12424
rect 1544 12384 1550 12396
rect 1762 12384 1768 12396
rect 1820 12384 1826 12436
rect 2409 12427 2467 12433
rect 2409 12393 2421 12427
rect 2455 12424 2467 12427
rect 2682 12424 2688 12436
rect 2455 12396 2688 12424
rect 2455 12393 2467 12396
rect 2409 12387 2467 12393
rect 2682 12384 2688 12396
rect 2740 12384 2746 12436
rect 2777 12427 2835 12433
rect 2777 12393 2789 12427
rect 2823 12424 2835 12427
rect 3142 12424 3148 12436
rect 2823 12396 3148 12424
rect 2823 12393 2835 12396
rect 2777 12387 2835 12393
rect 3142 12384 3148 12396
rect 3200 12424 3206 12436
rect 3510 12424 3516 12436
rect 3200 12396 3516 12424
rect 3200 12384 3206 12396
rect 3510 12384 3516 12396
rect 3568 12384 3574 12436
rect 4249 12427 4307 12433
rect 4249 12393 4261 12427
rect 4295 12424 4307 12427
rect 4430 12424 4436 12436
rect 4295 12396 4436 12424
rect 4295 12393 4307 12396
rect 4249 12387 4307 12393
rect 4430 12384 4436 12396
rect 4488 12384 4494 12436
rect 7742 12424 7748 12436
rect 7703 12396 7748 12424
rect 7742 12384 7748 12396
rect 7800 12384 7806 12436
rect 8110 12384 8116 12436
rect 8168 12384 8174 12436
rect 8849 12427 8907 12433
rect 8849 12393 8861 12427
rect 8895 12424 8907 12427
rect 9582 12424 9588 12436
rect 8895 12396 9588 12424
rect 8895 12393 8907 12396
rect 8849 12387 8907 12393
rect 4801 12359 4859 12365
rect 4801 12356 4813 12359
rect 4264 12328 4813 12356
rect 4264 12300 4292 12328
rect 4801 12325 4813 12328
rect 4847 12356 4859 12359
rect 7098 12356 7104 12368
rect 4847 12328 7104 12356
rect 4847 12325 4859 12328
rect 4801 12319 4859 12325
rect 7098 12316 7104 12328
rect 7156 12316 7162 12368
rect 7653 12359 7711 12365
rect 7653 12325 7665 12359
rect 7699 12356 7711 12359
rect 8128 12356 8156 12384
rect 7699 12328 8156 12356
rect 7699 12325 7711 12328
rect 7653 12319 7711 12325
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1946 12288 1952 12300
rect 1443 12260 1952 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1946 12248 1952 12260
rect 2004 12248 2010 12300
rect 2038 12248 2044 12300
rect 2096 12248 2102 12300
rect 2869 12291 2927 12297
rect 2869 12257 2881 12291
rect 2915 12288 2927 12291
rect 3326 12288 3332 12300
rect 2915 12260 3332 12288
rect 2915 12257 2927 12260
rect 2869 12251 2927 12257
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 4246 12248 4252 12300
rect 4304 12248 4310 12300
rect 5629 12291 5687 12297
rect 5629 12257 5641 12291
rect 5675 12288 5687 12291
rect 6178 12288 6184 12300
rect 5675 12260 6184 12288
rect 5675 12257 5687 12260
rect 5629 12251 5687 12257
rect 6178 12248 6184 12260
rect 6236 12248 6242 12300
rect 8113 12291 8171 12297
rect 8113 12257 8125 12291
rect 8159 12288 8171 12291
rect 8864 12288 8892 12387
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 11790 12424 11796 12436
rect 11751 12396 11796 12424
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 14182 12424 14188 12436
rect 12492 12396 12537 12424
rect 14143 12396 14188 12424
rect 12492 12384 12498 12396
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 14458 12384 14464 12436
rect 14516 12424 14522 12436
rect 14553 12427 14611 12433
rect 14553 12424 14565 12427
rect 14516 12396 14565 12424
rect 14516 12384 14522 12396
rect 14553 12393 14565 12396
rect 14599 12393 14611 12427
rect 15286 12424 15292 12436
rect 15247 12396 15292 12424
rect 14553 12387 14611 12393
rect 15286 12384 15292 12396
rect 15344 12384 15350 12436
rect 15838 12424 15844 12436
rect 15799 12396 15844 12424
rect 15838 12384 15844 12396
rect 15896 12384 15902 12436
rect 17954 12384 17960 12436
rect 18012 12424 18018 12436
rect 18509 12427 18567 12433
rect 18509 12424 18521 12427
rect 18012 12396 18521 12424
rect 18012 12384 18018 12396
rect 18509 12393 18521 12396
rect 18555 12393 18567 12427
rect 19058 12424 19064 12436
rect 19019 12396 19064 12424
rect 18509 12387 18567 12393
rect 19058 12384 19064 12396
rect 19116 12384 19122 12436
rect 21818 12424 21824 12436
rect 21779 12396 21824 12424
rect 21818 12384 21824 12396
rect 21876 12384 21882 12436
rect 24026 12384 24032 12436
rect 24084 12424 24090 12436
rect 24765 12427 24823 12433
rect 24765 12424 24777 12427
rect 24084 12396 24777 12424
rect 24084 12384 24090 12396
rect 24765 12393 24777 12396
rect 24811 12393 24823 12427
rect 24765 12387 24823 12393
rect 10680 12359 10738 12365
rect 10680 12325 10692 12359
rect 10726 12356 10738 12359
rect 10870 12356 10876 12368
rect 10726 12328 10876 12356
rect 10726 12325 10738 12328
rect 10680 12319 10738 12325
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 12158 12316 12164 12368
rect 12216 12356 12222 12368
rect 12986 12356 12992 12368
rect 12216 12328 12992 12356
rect 12216 12316 12222 12328
rect 12986 12316 12992 12328
rect 13044 12356 13050 12368
rect 13633 12359 13691 12365
rect 13633 12356 13645 12359
rect 13044 12328 13645 12356
rect 13044 12316 13050 12328
rect 13633 12325 13645 12328
rect 13679 12325 13691 12359
rect 13633 12319 13691 12325
rect 13906 12316 13912 12368
rect 13964 12356 13970 12368
rect 14921 12359 14979 12365
rect 14921 12356 14933 12359
rect 13964 12328 14933 12356
rect 13964 12316 13970 12328
rect 14921 12325 14933 12328
rect 14967 12325 14979 12359
rect 22094 12356 22100 12368
rect 14921 12319 14979 12325
rect 22020 12328 22100 12356
rect 8159 12260 8892 12288
rect 8159 12257 8171 12260
rect 8113 12251 8171 12257
rect 9858 12248 9864 12300
rect 9916 12288 9922 12300
rect 10962 12288 10968 12300
rect 9916 12260 10968 12288
rect 9916 12248 9922 12260
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 13170 12248 13176 12300
rect 13228 12288 13234 12300
rect 13541 12291 13599 12297
rect 13541 12288 13553 12291
rect 13228 12260 13553 12288
rect 13228 12248 13234 12260
rect 13541 12257 13553 12260
rect 13587 12257 13599 12291
rect 13541 12251 13599 12257
rect 16844 12291 16902 12297
rect 16844 12257 16856 12291
rect 16890 12288 16902 12291
rect 17310 12288 17316 12300
rect 16890 12260 17316 12288
rect 16890 12257 16902 12260
rect 16844 12251 16902 12257
rect 17310 12248 17316 12260
rect 17368 12248 17374 12300
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 22020 12297 22048 12328
rect 22094 12316 22100 12328
rect 22152 12316 22158 12368
rect 22278 12297 22284 12300
rect 19429 12291 19487 12297
rect 19429 12288 19441 12291
rect 19392 12260 19441 12288
rect 19392 12248 19398 12260
rect 19429 12257 19441 12260
rect 19475 12288 19487 12291
rect 20441 12291 20499 12297
rect 20441 12288 20453 12291
rect 19475 12260 20453 12288
rect 19475 12257 19487 12260
rect 19429 12251 19487 12257
rect 20441 12257 20453 12260
rect 20487 12257 20499 12291
rect 20441 12251 20499 12257
rect 22005 12291 22063 12297
rect 22005 12257 22017 12291
rect 22051 12257 22063 12291
rect 22005 12251 22063 12257
rect 22272 12251 22284 12297
rect 22336 12288 22342 12300
rect 24581 12291 24639 12297
rect 22336 12260 22372 12288
rect 22278 12248 22284 12251
rect 22336 12248 22342 12260
rect 24581 12257 24593 12291
rect 24627 12288 24639 12291
rect 24670 12288 24676 12300
rect 24627 12260 24676 12288
rect 24627 12257 24639 12260
rect 24581 12251 24639 12257
rect 24670 12248 24676 12260
rect 24728 12248 24734 12300
rect 1854 12180 1860 12232
rect 1912 12220 1918 12232
rect 2056 12220 2084 12248
rect 1912 12192 2084 12220
rect 2317 12223 2375 12229
rect 1912 12180 1918 12192
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 3053 12223 3111 12229
rect 3053 12220 3065 12223
rect 2363 12192 3065 12220
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 3053 12189 3065 12192
rect 3099 12220 3111 12223
rect 5166 12220 5172 12232
rect 3099 12192 5172 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 5166 12180 5172 12192
rect 5224 12180 5230 12232
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 5721 12223 5779 12229
rect 5721 12220 5733 12223
rect 5592 12192 5733 12220
rect 5592 12180 5598 12192
rect 5721 12189 5733 12192
rect 5767 12189 5779 12223
rect 5721 12183 5779 12189
rect 5905 12223 5963 12229
rect 5905 12189 5917 12223
rect 5951 12220 5963 12223
rect 6454 12220 6460 12232
rect 5951 12192 6460 12220
rect 5951 12189 5963 12192
rect 5905 12183 5963 12189
rect 6454 12180 6460 12192
rect 6512 12180 6518 12232
rect 7006 12180 7012 12232
rect 7064 12220 7070 12232
rect 7742 12220 7748 12232
rect 7064 12192 7748 12220
rect 7064 12180 7070 12192
rect 7742 12180 7748 12192
rect 7800 12220 7806 12232
rect 8205 12223 8263 12229
rect 8205 12220 8217 12223
rect 7800 12192 8217 12220
rect 7800 12180 7806 12192
rect 8205 12189 8217 12192
rect 8251 12189 8263 12223
rect 8205 12183 8263 12189
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12220 8355 12223
rect 8478 12220 8484 12232
rect 8343 12192 8484 12220
rect 8343 12189 8355 12192
rect 8297 12183 8355 12189
rect 1581 12155 1639 12161
rect 1581 12121 1593 12155
rect 1627 12152 1639 12155
rect 2498 12152 2504 12164
rect 1627 12124 2504 12152
rect 1627 12121 1639 12124
rect 1581 12115 1639 12121
rect 2498 12112 2504 12124
rect 2556 12112 2562 12164
rect 4154 12112 4160 12164
rect 4212 12152 4218 12164
rect 5261 12155 5319 12161
rect 5261 12152 5273 12155
rect 4212 12124 5273 12152
rect 4212 12112 4218 12124
rect 5261 12121 5273 12124
rect 5307 12121 5319 12155
rect 5261 12115 5319 12121
rect 5994 12112 6000 12164
rect 6052 12152 6058 12164
rect 6052 12124 8064 12152
rect 6052 12112 6058 12124
rect 1946 12084 1952 12096
rect 1907 12056 1952 12084
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 3234 12044 3240 12096
rect 3292 12084 3298 12096
rect 3421 12087 3479 12093
rect 3421 12084 3433 12087
rect 3292 12056 3433 12084
rect 3292 12044 3298 12056
rect 3421 12053 3433 12056
rect 3467 12053 3479 12087
rect 3421 12047 3479 12053
rect 3881 12087 3939 12093
rect 3881 12053 3893 12087
rect 3927 12084 3939 12087
rect 3970 12084 3976 12096
rect 3927 12056 3976 12084
rect 3927 12053 3939 12056
rect 3881 12047 3939 12053
rect 3970 12044 3976 12056
rect 4028 12044 4034 12096
rect 5166 12084 5172 12096
rect 5127 12056 5172 12084
rect 5166 12044 5172 12056
rect 5224 12044 5230 12096
rect 6270 12084 6276 12096
rect 6231 12056 6276 12084
rect 6270 12044 6276 12056
rect 6328 12044 6334 12096
rect 6638 12084 6644 12096
rect 6599 12056 6644 12084
rect 6638 12044 6644 12056
rect 6696 12044 6702 12096
rect 7193 12087 7251 12093
rect 7193 12053 7205 12087
rect 7239 12084 7251 12087
rect 7374 12084 7380 12096
rect 7239 12056 7380 12084
rect 7239 12053 7251 12056
rect 7193 12047 7251 12053
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 8036 12084 8064 12124
rect 8110 12112 8116 12164
rect 8168 12152 8174 12164
rect 8312 12152 8340 12183
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 9490 12220 9496 12232
rect 9403 12192 9496 12220
rect 9490 12180 9496 12192
rect 9548 12220 9554 12232
rect 10229 12223 10287 12229
rect 10229 12220 10241 12223
rect 9548 12192 10241 12220
rect 9548 12180 9554 12192
rect 10229 12189 10241 12192
rect 10275 12189 10287 12223
rect 10410 12220 10416 12232
rect 10371 12192 10416 12220
rect 10229 12183 10287 12189
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12220 13139 12223
rect 13817 12223 13875 12229
rect 13817 12220 13829 12223
rect 13127 12192 13829 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 13817 12189 13829 12192
rect 13863 12220 13875 12223
rect 13906 12220 13912 12232
rect 13863 12192 13912 12220
rect 13863 12189 13875 12192
rect 13817 12183 13875 12189
rect 13906 12180 13912 12192
rect 13964 12180 13970 12232
rect 16022 12180 16028 12232
rect 16080 12220 16086 12232
rect 16574 12220 16580 12232
rect 16080 12192 16580 12220
rect 16080 12180 16086 12192
rect 16574 12180 16580 12192
rect 16632 12180 16638 12232
rect 19518 12220 19524 12232
rect 19479 12192 19524 12220
rect 19518 12180 19524 12192
rect 19576 12180 19582 12232
rect 19610 12180 19616 12232
rect 19668 12220 19674 12232
rect 20901 12223 20959 12229
rect 19668 12192 19713 12220
rect 19668 12180 19674 12192
rect 20901 12189 20913 12223
rect 20947 12220 20959 12223
rect 21266 12220 21272 12232
rect 20947 12192 21272 12220
rect 20947 12189 20959 12192
rect 20901 12183 20959 12189
rect 21266 12180 21272 12192
rect 21324 12180 21330 12232
rect 8168 12124 8340 12152
rect 13173 12155 13231 12161
rect 8168 12112 8174 12124
rect 13173 12121 13185 12155
rect 13219 12152 13231 12155
rect 13446 12152 13452 12164
rect 13219 12124 13452 12152
rect 13219 12121 13231 12124
rect 13173 12115 13231 12121
rect 13446 12112 13452 12124
rect 13504 12112 13510 12164
rect 19536 12152 19564 12180
rect 20073 12155 20131 12161
rect 20073 12152 20085 12155
rect 19536 12124 20085 12152
rect 20073 12121 20085 12124
rect 20119 12121 20131 12155
rect 20073 12115 20131 12121
rect 8386 12084 8392 12096
rect 8036 12056 8392 12084
rect 8386 12044 8392 12056
rect 8444 12084 8450 12096
rect 9490 12084 9496 12096
rect 8444 12056 9496 12084
rect 8444 12044 8450 12056
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 9953 12087 10011 12093
rect 9953 12053 9965 12087
rect 9999 12084 10011 12087
rect 10042 12084 10048 12096
rect 9999 12056 10048 12084
rect 9999 12053 10011 12056
rect 9953 12047 10011 12053
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 15562 12044 15568 12096
rect 15620 12084 15626 12096
rect 16117 12087 16175 12093
rect 16117 12084 16129 12087
rect 15620 12056 16129 12084
rect 15620 12044 15626 12056
rect 16117 12053 16129 12056
rect 16163 12053 16175 12087
rect 17954 12084 17960 12096
rect 17915 12056 17960 12084
rect 16117 12047 16175 12053
rect 17954 12044 17960 12056
rect 18012 12044 18018 12096
rect 18966 12084 18972 12096
rect 18879 12056 18972 12084
rect 18966 12044 18972 12056
rect 19024 12084 19030 12096
rect 19610 12084 19616 12096
rect 19024 12056 19616 12084
rect 19024 12044 19030 12056
rect 19610 12044 19616 12056
rect 19668 12044 19674 12096
rect 20990 12044 20996 12096
rect 21048 12084 21054 12096
rect 21453 12087 21511 12093
rect 21453 12084 21465 12087
rect 21048 12056 21465 12084
rect 21048 12044 21054 12056
rect 21453 12053 21465 12056
rect 21499 12053 21511 12087
rect 21453 12047 21511 12053
rect 23385 12087 23443 12093
rect 23385 12053 23397 12087
rect 23431 12084 23443 12087
rect 24026 12084 24032 12096
rect 23431 12056 24032 12084
rect 23431 12053 23443 12056
rect 23385 12047 23443 12053
rect 24026 12044 24032 12056
rect 24084 12044 24090 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2222 11880 2228 11892
rect 2183 11852 2228 11880
rect 2222 11840 2228 11852
rect 2280 11840 2286 11892
rect 2314 11840 2320 11892
rect 2372 11880 2378 11892
rect 2498 11880 2504 11892
rect 2372 11852 2504 11880
rect 2372 11840 2378 11852
rect 2498 11840 2504 11852
rect 2556 11840 2562 11892
rect 3326 11880 3332 11892
rect 3239 11852 3332 11880
rect 3326 11840 3332 11852
rect 3384 11880 3390 11892
rect 5166 11880 5172 11892
rect 3384 11852 5028 11880
rect 5079 11852 5172 11880
rect 3384 11840 3390 11852
rect 1765 11815 1823 11821
rect 1765 11781 1777 11815
rect 1811 11812 1823 11815
rect 3142 11812 3148 11824
rect 1811 11784 3148 11812
rect 1811 11781 1823 11784
rect 1765 11775 1823 11781
rect 3142 11772 3148 11784
rect 3200 11772 3206 11824
rect 5000 11812 5028 11852
rect 5166 11840 5172 11852
rect 5224 11880 5230 11892
rect 6454 11880 6460 11892
rect 5224 11852 6460 11880
rect 5224 11840 5230 11852
rect 6454 11840 6460 11852
rect 6512 11840 6518 11892
rect 9030 11880 9036 11892
rect 6656 11852 9036 11880
rect 6656 11812 6684 11852
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 9582 11840 9588 11892
rect 9640 11840 9646 11892
rect 9677 11883 9735 11889
rect 9677 11849 9689 11883
rect 9723 11880 9735 11883
rect 9766 11880 9772 11892
rect 9723 11852 9772 11880
rect 9723 11849 9735 11852
rect 9677 11843 9735 11849
rect 9766 11840 9772 11852
rect 9824 11880 9830 11892
rect 10597 11883 10655 11889
rect 10597 11880 10609 11883
rect 9824 11852 10609 11880
rect 9824 11840 9830 11852
rect 10597 11849 10609 11852
rect 10643 11849 10655 11883
rect 13170 11880 13176 11892
rect 13131 11852 13176 11880
rect 10597 11843 10655 11849
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 15654 11840 15660 11892
rect 15712 11880 15718 11892
rect 16117 11883 16175 11889
rect 16117 11880 16129 11883
rect 15712 11852 16129 11880
rect 15712 11840 15718 11852
rect 16117 11849 16129 11852
rect 16163 11880 16175 11883
rect 17218 11880 17224 11892
rect 16163 11852 17224 11880
rect 16163 11849 16175 11852
rect 16117 11843 16175 11849
rect 17218 11840 17224 11852
rect 17276 11840 17282 11892
rect 17310 11840 17316 11892
rect 17368 11880 17374 11892
rect 17497 11883 17555 11889
rect 17497 11880 17509 11883
rect 17368 11852 17509 11880
rect 17368 11840 17374 11852
rect 17497 11849 17509 11852
rect 17543 11849 17555 11883
rect 17497 11843 17555 11849
rect 22094 11840 22100 11892
rect 22152 11880 22158 11892
rect 22833 11883 22891 11889
rect 22833 11880 22845 11883
rect 22152 11852 22845 11880
rect 22152 11840 22158 11852
rect 22833 11849 22845 11852
rect 22879 11880 22891 11883
rect 23385 11883 23443 11889
rect 23385 11880 23397 11883
rect 22879 11852 23397 11880
rect 22879 11849 22891 11852
rect 22833 11843 22891 11849
rect 23385 11849 23397 11852
rect 23431 11849 23443 11883
rect 23385 11843 23443 11849
rect 9600 11812 9628 11840
rect 5000 11784 6684 11812
rect 8312 11784 9628 11812
rect 1946 11704 1952 11756
rect 2004 11744 2010 11756
rect 2777 11747 2835 11753
rect 2777 11744 2789 11747
rect 2004 11716 2789 11744
rect 2004 11704 2010 11716
rect 2777 11713 2789 11716
rect 2823 11713 2835 11747
rect 2777 11707 2835 11713
rect 2314 11568 2320 11620
rect 2372 11608 2378 11620
rect 2682 11608 2688 11620
rect 2372 11580 2688 11608
rect 2372 11568 2378 11580
rect 2682 11568 2688 11580
rect 2740 11568 2746 11620
rect 2133 11543 2191 11549
rect 2133 11509 2145 11543
rect 2179 11540 2191 11543
rect 2590 11540 2596 11552
rect 2179 11512 2596 11540
rect 2179 11509 2191 11512
rect 2133 11503 2191 11509
rect 2590 11500 2596 11512
rect 2648 11500 2654 11552
rect 2792 11540 2820 11707
rect 3697 11679 3755 11685
rect 3697 11645 3709 11679
rect 3743 11676 3755 11679
rect 3789 11679 3847 11685
rect 3789 11676 3801 11679
rect 3743 11648 3801 11676
rect 3743 11645 3755 11648
rect 3697 11639 3755 11645
rect 3789 11645 3801 11648
rect 3835 11676 3847 11679
rect 3835 11648 4292 11676
rect 3835 11645 3847 11648
rect 3789 11639 3847 11645
rect 4264 11620 4292 11648
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 7193 11679 7251 11685
rect 7193 11676 7205 11679
rect 7156 11648 7205 11676
rect 7156 11636 7162 11648
rect 7193 11645 7205 11648
rect 7239 11676 7251 11679
rect 7282 11676 7288 11688
rect 7239 11648 7288 11676
rect 7239 11645 7251 11648
rect 7193 11639 7251 11645
rect 7282 11636 7288 11648
rect 7340 11636 7346 11688
rect 7558 11685 7564 11688
rect 7552 11676 7564 11685
rect 7471 11648 7564 11676
rect 7552 11639 7564 11648
rect 7616 11676 7622 11688
rect 8312 11676 8340 11784
rect 10042 11772 10048 11824
rect 10100 11812 10106 11824
rect 10962 11812 10968 11824
rect 10100 11784 10968 11812
rect 10100 11772 10106 11784
rect 10962 11772 10968 11784
rect 11020 11772 11026 11824
rect 15013 11815 15071 11821
rect 15013 11781 15025 11815
rect 15059 11812 15071 11815
rect 15102 11812 15108 11824
rect 15059 11784 15108 11812
rect 15059 11781 15071 11784
rect 15013 11775 15071 11781
rect 15102 11772 15108 11784
rect 15160 11812 15166 11824
rect 15930 11812 15936 11824
rect 15160 11784 15936 11812
rect 15160 11772 15166 11784
rect 15930 11772 15936 11784
rect 15988 11772 15994 11824
rect 18966 11772 18972 11824
rect 19024 11812 19030 11824
rect 19242 11812 19248 11824
rect 19024 11784 19248 11812
rect 19024 11772 19030 11784
rect 19242 11772 19248 11784
rect 19300 11772 19306 11824
rect 21450 11772 21456 11824
rect 21508 11812 21514 11824
rect 21634 11812 21640 11824
rect 21508 11784 21640 11812
rect 21508 11772 21514 11784
rect 21634 11772 21640 11784
rect 21692 11772 21698 11824
rect 8386 11704 8392 11756
rect 8444 11744 8450 11756
rect 9582 11744 9588 11756
rect 8444 11716 9588 11744
rect 8444 11704 8450 11716
rect 9582 11704 9588 11716
rect 9640 11704 9646 11756
rect 10321 11747 10379 11753
rect 10321 11713 10333 11747
rect 10367 11713 10379 11747
rect 10321 11707 10379 11713
rect 11333 11747 11391 11753
rect 11333 11713 11345 11747
rect 11379 11744 11391 11747
rect 11422 11744 11428 11756
rect 11379 11716 11428 11744
rect 11379 11713 11391 11716
rect 11333 11707 11391 11713
rect 7616 11648 8340 11676
rect 7558 11636 7564 11639
rect 7616 11636 7622 11648
rect 9030 11636 9036 11688
rect 9088 11676 9094 11688
rect 9493 11679 9551 11685
rect 9493 11676 9505 11679
rect 9088 11648 9505 11676
rect 9088 11636 9094 11648
rect 9493 11645 9505 11648
rect 9539 11645 9551 11679
rect 9493 11639 9551 11645
rect 10042 11636 10048 11688
rect 10100 11676 10106 11688
rect 10336 11676 10364 11707
rect 11422 11704 11428 11716
rect 11480 11704 11486 11756
rect 14642 11704 14648 11756
rect 14700 11744 14706 11756
rect 15657 11747 15715 11753
rect 15657 11744 15669 11747
rect 14700 11716 15669 11744
rect 14700 11704 14706 11716
rect 15657 11713 15669 11716
rect 15703 11744 15715 11747
rect 16761 11747 16819 11753
rect 16761 11744 16773 11747
rect 15703 11716 16773 11744
rect 15703 11713 15715 11716
rect 15657 11707 15715 11713
rect 16761 11713 16773 11716
rect 16807 11744 16819 11747
rect 17954 11744 17960 11756
rect 16807 11716 17960 11744
rect 16807 11713 16819 11716
rect 16761 11707 16819 11713
rect 17954 11704 17960 11716
rect 18012 11704 18018 11756
rect 20990 11704 20996 11756
rect 21048 11744 21054 11756
rect 22373 11747 22431 11753
rect 22373 11744 22385 11747
rect 21048 11716 22385 11744
rect 21048 11704 21054 11716
rect 22373 11713 22385 11716
rect 22419 11713 22431 11747
rect 23400 11744 23428 11843
rect 23661 11747 23719 11753
rect 23661 11744 23673 11747
rect 23400 11716 23673 11744
rect 22373 11707 22431 11713
rect 23661 11713 23673 11716
rect 23707 11713 23719 11747
rect 23661 11707 23719 11713
rect 10100 11648 10364 11676
rect 10597 11679 10655 11685
rect 10100 11636 10106 11648
rect 10597 11645 10609 11679
rect 10643 11676 10655 11679
rect 12618 11676 12624 11688
rect 10643 11648 12624 11676
rect 10643 11645 10655 11648
rect 10597 11639 10655 11645
rect 12618 11636 12624 11648
rect 12676 11636 12682 11688
rect 13630 11676 13636 11688
rect 13543 11648 13636 11676
rect 13630 11636 13636 11648
rect 13688 11636 13694 11688
rect 13906 11685 13912 11688
rect 13900 11676 13912 11685
rect 13819 11648 13912 11676
rect 13900 11639 13912 11648
rect 13964 11676 13970 11688
rect 14660 11676 14688 11704
rect 13964 11648 14688 11676
rect 13906 11636 13912 11639
rect 13964 11636 13970 11648
rect 15562 11636 15568 11688
rect 15620 11676 15626 11688
rect 16577 11679 16635 11685
rect 16577 11676 16589 11679
rect 15620 11648 16589 11676
rect 15620 11636 15626 11648
rect 16577 11645 16589 11648
rect 16623 11645 16635 11679
rect 16577 11639 16635 11645
rect 19242 11636 19248 11688
rect 19300 11676 19306 11688
rect 19337 11679 19395 11685
rect 19337 11676 19349 11679
rect 19300 11648 19349 11676
rect 19300 11636 19306 11648
rect 19337 11645 19349 11648
rect 19383 11645 19395 11679
rect 21358 11676 21364 11688
rect 21271 11648 21364 11676
rect 19337 11639 19395 11645
rect 21358 11636 21364 11648
rect 21416 11676 21422 11688
rect 22278 11676 22284 11688
rect 21416 11648 22284 11676
rect 21416 11636 21422 11648
rect 22278 11636 22284 11648
rect 22336 11636 22342 11688
rect 4062 11617 4068 11620
rect 4056 11608 4068 11617
rect 4023 11580 4068 11608
rect 4056 11571 4068 11580
rect 4062 11568 4068 11571
rect 4120 11568 4126 11620
rect 4246 11568 4252 11620
rect 4304 11568 4310 11620
rect 5534 11568 5540 11620
rect 5592 11608 5598 11620
rect 5813 11611 5871 11617
rect 5813 11608 5825 11611
rect 5592 11580 5825 11608
rect 5592 11568 5598 11580
rect 5813 11577 5825 11580
rect 5859 11608 5871 11611
rect 6546 11608 6552 11620
rect 5859 11580 6552 11608
rect 5859 11577 5871 11580
rect 5813 11571 5871 11577
rect 6546 11568 6552 11580
rect 6604 11568 6610 11620
rect 7926 11568 7932 11620
rect 7984 11608 7990 11620
rect 8846 11608 8852 11620
rect 7984 11580 8852 11608
rect 7984 11568 7990 11580
rect 8846 11568 8852 11580
rect 8904 11568 8910 11620
rect 10137 11611 10195 11617
rect 10137 11608 10149 11611
rect 9324 11580 10149 11608
rect 9324 11552 9352 11580
rect 10137 11577 10149 11580
rect 10183 11577 10195 11611
rect 10137 11571 10195 11577
rect 10410 11568 10416 11620
rect 10468 11608 10474 11620
rect 10781 11611 10839 11617
rect 10781 11608 10793 11611
rect 10468 11580 10793 11608
rect 10468 11568 10474 11580
rect 10781 11577 10793 11580
rect 10827 11608 10839 11611
rect 11146 11608 11152 11620
rect 10827 11580 11152 11608
rect 10827 11577 10839 11580
rect 10781 11571 10839 11577
rect 11146 11568 11152 11580
rect 11204 11568 11210 11620
rect 13648 11608 13676 11636
rect 13998 11608 14004 11620
rect 13648 11580 14004 11608
rect 13998 11568 14004 11580
rect 14056 11568 14062 11620
rect 19582 11611 19640 11617
rect 19582 11608 19594 11611
rect 18800 11580 19594 11608
rect 18800 11552 18828 11580
rect 19582 11577 19594 11580
rect 19628 11577 19640 11611
rect 19582 11571 19640 11577
rect 21082 11568 21088 11620
rect 21140 11608 21146 11620
rect 21637 11611 21695 11617
rect 21637 11608 21649 11611
rect 21140 11580 21649 11608
rect 21140 11568 21146 11580
rect 21637 11577 21649 11580
rect 21683 11608 21695 11611
rect 22189 11611 22247 11617
rect 22189 11608 22201 11611
rect 21683 11580 22201 11608
rect 21683 11577 21695 11580
rect 21637 11571 21695 11577
rect 22189 11577 22201 11580
rect 22235 11577 22247 11611
rect 22189 11571 22247 11577
rect 23928 11611 23986 11617
rect 23928 11577 23940 11611
rect 23974 11608 23986 11611
rect 24026 11608 24032 11620
rect 23974 11580 24032 11608
rect 23974 11577 23986 11580
rect 23928 11571 23986 11577
rect 24026 11568 24032 11580
rect 24084 11568 24090 11620
rect 5994 11540 6000 11552
rect 2792 11512 6000 11540
rect 5994 11500 6000 11512
rect 6052 11500 6058 11552
rect 6178 11540 6184 11552
rect 6139 11512 6184 11540
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 8665 11543 8723 11549
rect 8665 11540 8677 11543
rect 8352 11512 8677 11540
rect 8352 11500 8358 11512
rect 8665 11509 8677 11512
rect 8711 11509 8723 11543
rect 9306 11540 9312 11552
rect 9267 11512 9312 11540
rect 8665 11503 8723 11509
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 9490 11540 9496 11552
rect 9451 11512 9496 11540
rect 9490 11500 9496 11512
rect 9548 11500 9554 11552
rect 9766 11540 9772 11552
rect 9727 11512 9772 11540
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 10229 11543 10287 11549
rect 10229 11509 10241 11543
rect 10275 11540 10287 11543
rect 10597 11543 10655 11549
rect 10597 11540 10609 11543
rect 10275 11512 10609 11540
rect 10275 11509 10287 11512
rect 10229 11503 10287 11509
rect 10597 11509 10609 11512
rect 10643 11509 10655 11543
rect 10597 11503 10655 11509
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11238 11540 11244 11552
rect 10928 11512 11244 11540
rect 10928 11500 10934 11512
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 11790 11540 11796 11552
rect 11751 11512 11796 11540
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 12066 11500 12072 11552
rect 12124 11540 12130 11552
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 12124 11512 12173 11540
rect 12124 11500 12130 11512
rect 12161 11509 12173 11512
rect 12207 11509 12219 11543
rect 12161 11503 12219 11509
rect 12621 11543 12679 11549
rect 12621 11509 12633 11543
rect 12667 11540 12679 11543
rect 13446 11540 13452 11552
rect 12667 11512 13452 11540
rect 12667 11509 12679 11512
rect 12621 11503 12679 11509
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 15930 11540 15936 11552
rect 15891 11512 15936 11540
rect 15930 11500 15936 11512
rect 15988 11540 15994 11552
rect 16485 11543 16543 11549
rect 16485 11540 16497 11543
rect 15988 11512 16497 11540
rect 15988 11500 15994 11512
rect 16485 11509 16497 11512
rect 16531 11509 16543 11543
rect 16485 11503 16543 11509
rect 16574 11500 16580 11552
rect 16632 11540 16638 11552
rect 17221 11543 17279 11549
rect 17221 11540 17233 11543
rect 16632 11512 17233 11540
rect 16632 11500 16638 11512
rect 17221 11509 17233 11512
rect 17267 11540 17279 11543
rect 17494 11540 17500 11552
rect 17267 11512 17500 11540
rect 17267 11509 17279 11512
rect 17221 11503 17279 11509
rect 17494 11500 17500 11512
rect 17552 11500 17558 11552
rect 18046 11500 18052 11552
rect 18104 11540 18110 11552
rect 18141 11543 18199 11549
rect 18141 11540 18153 11543
rect 18104 11512 18153 11540
rect 18104 11500 18110 11512
rect 18141 11509 18153 11512
rect 18187 11509 18199 11543
rect 18782 11540 18788 11552
rect 18743 11512 18788 11540
rect 18141 11503 18199 11509
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 19242 11540 19248 11552
rect 19203 11512 19248 11540
rect 19242 11500 19248 11512
rect 19300 11500 19306 11552
rect 20717 11543 20775 11549
rect 20717 11509 20729 11543
rect 20763 11540 20775 11543
rect 20990 11540 20996 11552
rect 20763 11512 20996 11540
rect 20763 11509 20775 11512
rect 20717 11503 20775 11509
rect 20990 11500 20996 11512
rect 21048 11500 21054 11552
rect 21726 11500 21732 11552
rect 21784 11540 21790 11552
rect 21821 11543 21879 11549
rect 21821 11540 21833 11543
rect 21784 11512 21833 11540
rect 21784 11500 21790 11512
rect 21821 11509 21833 11512
rect 21867 11509 21879 11543
rect 21821 11503 21879 11509
rect 21910 11500 21916 11552
rect 21968 11540 21974 11552
rect 22281 11543 22339 11549
rect 22281 11540 22293 11543
rect 21968 11512 22293 11540
rect 21968 11500 21974 11512
rect 22281 11509 22293 11512
rect 22327 11509 22339 11543
rect 22281 11503 22339 11509
rect 24854 11500 24860 11552
rect 24912 11540 24918 11552
rect 25041 11543 25099 11549
rect 25041 11540 25053 11543
rect 24912 11512 25053 11540
rect 24912 11500 24918 11512
rect 25041 11509 25053 11512
rect 25087 11509 25099 11543
rect 25041 11503 25099 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1486 11296 1492 11348
rect 1544 11336 1550 11348
rect 1581 11339 1639 11345
rect 1581 11336 1593 11339
rect 1544 11308 1593 11336
rect 1544 11296 1550 11308
rect 1581 11305 1593 11308
rect 1627 11305 1639 11339
rect 2314 11336 2320 11348
rect 2275 11308 2320 11336
rect 1581 11299 1639 11305
rect 2314 11296 2320 11308
rect 2372 11296 2378 11348
rect 2406 11296 2412 11348
rect 2464 11336 2470 11348
rect 2685 11339 2743 11345
rect 2685 11336 2697 11339
rect 2464 11308 2697 11336
rect 2464 11296 2470 11308
rect 2685 11305 2697 11308
rect 2731 11305 2743 11339
rect 2685 11299 2743 11305
rect 4065 11339 4123 11345
rect 4065 11305 4077 11339
rect 4111 11305 4123 11339
rect 4065 11299 4123 11305
rect 2038 11228 2044 11280
rect 2096 11268 2102 11280
rect 4080 11268 4108 11299
rect 4338 11296 4344 11348
rect 4396 11336 4402 11348
rect 4433 11339 4491 11345
rect 4433 11336 4445 11339
rect 4396 11308 4445 11336
rect 4396 11296 4402 11308
rect 4433 11305 4445 11308
rect 4479 11336 4491 11339
rect 6638 11336 6644 11348
rect 4479 11308 6644 11336
rect 4479 11305 4491 11308
rect 4433 11299 4491 11305
rect 6638 11296 6644 11308
rect 6696 11296 6702 11348
rect 7006 11336 7012 11348
rect 6967 11308 7012 11336
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 7377 11339 7435 11345
rect 7377 11305 7389 11339
rect 7423 11336 7435 11339
rect 7558 11336 7564 11348
rect 7423 11308 7564 11336
rect 7423 11305 7435 11308
rect 7377 11299 7435 11305
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 7650 11296 7656 11348
rect 7708 11336 7714 11348
rect 8021 11339 8079 11345
rect 8021 11336 8033 11339
rect 7708 11308 8033 11336
rect 7708 11296 7714 11308
rect 8021 11305 8033 11308
rect 8067 11305 8079 11339
rect 8021 11299 8079 11305
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 9677 11339 9735 11345
rect 9677 11336 9689 11339
rect 9364 11308 9689 11336
rect 9364 11296 9370 11308
rect 9677 11305 9689 11308
rect 9723 11305 9735 11339
rect 9677 11299 9735 11305
rect 11238 11296 11244 11348
rect 11296 11336 11302 11348
rect 12069 11339 12127 11345
rect 12069 11336 12081 11339
rect 11296 11308 12081 11336
rect 11296 11296 11302 11308
rect 12069 11305 12081 11308
rect 12115 11305 12127 11339
rect 12986 11336 12992 11348
rect 12947 11308 12992 11336
rect 12069 11299 12127 11305
rect 12986 11296 12992 11308
rect 13044 11296 13050 11348
rect 13170 11336 13176 11348
rect 13131 11308 13176 11336
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 14642 11336 14648 11348
rect 14603 11308 14648 11336
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 15102 11336 15108 11348
rect 15063 11308 15108 11336
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 16669 11339 16727 11345
rect 16669 11305 16681 11339
rect 16715 11305 16727 11339
rect 17218 11336 17224 11348
rect 17179 11308 17224 11336
rect 16669 11299 16727 11305
rect 4522 11268 4528 11280
rect 2096 11240 4108 11268
rect 4435 11240 4528 11268
rect 2096 11228 2102 11240
rect 4522 11228 4528 11240
rect 4580 11268 4586 11280
rect 6270 11268 6276 11280
rect 4580 11240 6276 11268
rect 4580 11228 4586 11240
rect 6270 11228 6276 11240
rect 6328 11228 6334 11280
rect 7837 11271 7895 11277
rect 7837 11237 7849 11271
rect 7883 11268 7895 11271
rect 8110 11268 8116 11280
rect 7883 11240 8116 11268
rect 7883 11237 7895 11240
rect 7837 11231 7895 11237
rect 8110 11228 8116 11240
rect 8168 11228 8174 11280
rect 8389 11271 8447 11277
rect 8389 11237 8401 11271
rect 8435 11268 8447 11271
rect 9125 11271 9183 11277
rect 9125 11268 9137 11271
rect 8435 11240 9137 11268
rect 8435 11237 8447 11240
rect 8389 11231 8447 11237
rect 9125 11237 9137 11240
rect 9171 11268 9183 11271
rect 9766 11268 9772 11280
rect 9171 11240 9772 11268
rect 9171 11237 9183 11240
rect 9125 11231 9183 11237
rect 9766 11228 9772 11240
rect 9824 11228 9830 11280
rect 10686 11228 10692 11280
rect 10744 11268 10750 11280
rect 10934 11271 10992 11277
rect 10934 11268 10946 11271
rect 10744 11240 10946 11268
rect 10744 11228 10750 11240
rect 10934 11237 10946 11240
rect 10980 11268 10992 11271
rect 11054 11268 11060 11280
rect 10980 11240 11060 11268
rect 10980 11237 10992 11240
rect 10934 11231 10992 11237
rect 11054 11228 11060 11240
rect 11112 11228 11118 11280
rect 12713 11271 12771 11277
rect 12713 11237 12725 11271
rect 12759 11268 12771 11271
rect 13078 11268 13084 11280
rect 12759 11240 13084 11268
rect 12759 11237 12771 11240
rect 12713 11231 12771 11237
rect 13078 11228 13084 11240
rect 13136 11228 13142 11280
rect 13541 11271 13599 11277
rect 13541 11237 13553 11271
rect 13587 11268 13599 11271
rect 13722 11268 13728 11280
rect 13587 11240 13728 11268
rect 13587 11237 13599 11240
rect 13541 11231 13599 11237
rect 13722 11228 13728 11240
rect 13780 11228 13786 11280
rect 15120 11268 15148 11296
rect 15534 11271 15592 11277
rect 15534 11268 15546 11271
rect 15120 11240 15546 11268
rect 15534 11237 15546 11240
rect 15580 11237 15592 11271
rect 15534 11231 15592 11237
rect 16574 11228 16580 11280
rect 16632 11268 16638 11280
rect 16684 11268 16712 11299
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 18138 11336 18144 11348
rect 17328 11308 18144 11336
rect 17328 11268 17356 11308
rect 18138 11296 18144 11308
rect 18196 11296 18202 11348
rect 18782 11296 18788 11348
rect 18840 11336 18846 11348
rect 19429 11339 19487 11345
rect 19429 11336 19441 11339
rect 18840 11308 19441 11336
rect 18840 11296 18846 11308
rect 19429 11305 19441 11308
rect 19475 11305 19487 11339
rect 19429 11299 19487 11305
rect 20717 11339 20775 11345
rect 20717 11305 20729 11339
rect 20763 11336 20775 11339
rect 21082 11336 21088 11348
rect 20763 11308 21088 11336
rect 20763 11305 20775 11308
rect 20717 11299 20775 11305
rect 21082 11296 21088 11308
rect 21140 11336 21146 11348
rect 21726 11336 21732 11348
rect 21140 11308 21732 11336
rect 21140 11296 21146 11308
rect 21726 11296 21732 11308
rect 21784 11296 21790 11348
rect 22278 11336 22284 11348
rect 22239 11308 22284 11336
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 23385 11339 23443 11345
rect 23385 11305 23397 11339
rect 23431 11336 23443 11339
rect 23842 11336 23848 11348
rect 23431 11308 23848 11336
rect 23431 11305 23443 11308
rect 23385 11299 23443 11305
rect 23842 11296 23848 11308
rect 23900 11296 23906 11348
rect 25222 11336 25228 11348
rect 25183 11308 25228 11336
rect 25222 11296 25228 11308
rect 25280 11296 25286 11348
rect 19242 11268 19248 11280
rect 16632 11240 17356 11268
rect 18064 11240 19248 11268
rect 16632 11228 16638 11240
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 2314 11200 2320 11212
rect 1443 11172 2320 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 2314 11160 2320 11172
rect 2372 11160 2378 11212
rect 2489 11203 2547 11209
rect 2489 11200 2501 11203
rect 2424 11172 2501 11200
rect 2424 10996 2452 11172
rect 2489 11169 2501 11172
rect 2535 11169 2547 11203
rect 2489 11163 2547 11169
rect 2866 11160 2872 11212
rect 2924 11200 2930 11212
rect 3050 11200 3056 11212
rect 2924 11172 3056 11200
rect 2924 11160 2930 11172
rect 3050 11160 3056 11172
rect 3108 11160 3114 11212
rect 3142 11160 3148 11212
rect 3200 11200 3206 11212
rect 5997 11203 6055 11209
rect 5997 11200 6009 11203
rect 3200 11172 6009 11200
rect 3200 11160 3206 11172
rect 5997 11169 6009 11172
rect 6043 11200 6055 11203
rect 6454 11200 6460 11212
rect 6043 11172 6460 11200
rect 6043 11169 6055 11172
rect 5997 11163 6055 11169
rect 6454 11160 6460 11172
rect 6512 11160 6518 11212
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11200 8539 11203
rect 9490 11200 9496 11212
rect 8527 11172 9496 11200
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 9490 11160 9496 11172
rect 9548 11160 9554 11212
rect 11238 11200 11244 11212
rect 10704 11172 11244 11200
rect 4614 11132 4620 11144
rect 4575 11104 4620 11132
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 6086 11132 6092 11144
rect 6047 11104 6092 11132
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 6181 11135 6239 11141
rect 6181 11101 6193 11135
rect 6227 11101 6239 11135
rect 8662 11132 8668 11144
rect 8623 11104 8668 11132
rect 6181 11095 6239 11101
rect 2866 11024 2872 11076
rect 2924 11064 2930 11076
rect 3421 11067 3479 11073
rect 3421 11064 3433 11067
rect 2924 11036 3433 11064
rect 2924 11024 2930 11036
rect 3421 11033 3433 11036
rect 3467 11033 3479 11067
rect 3421 11027 3479 11033
rect 3881 11067 3939 11073
rect 3881 11033 3893 11067
rect 3927 11064 3939 11067
rect 4062 11064 4068 11076
rect 3927 11036 4068 11064
rect 3927 11033 3939 11036
rect 3881 11027 3939 11033
rect 4062 11024 4068 11036
rect 4120 11064 4126 11076
rect 4632 11064 4660 11092
rect 4120 11036 4660 11064
rect 5537 11067 5595 11073
rect 4120 11024 4126 11036
rect 5537 11033 5549 11067
rect 5583 11064 5595 11067
rect 5994 11064 6000 11076
rect 5583 11036 6000 11064
rect 5583 11033 5595 11036
rect 5537 11027 5595 11033
rect 5994 11024 6000 11036
rect 6052 11064 6058 11076
rect 6196 11064 6224 11095
rect 8662 11092 8668 11104
rect 8720 11092 8726 11144
rect 10704 11141 10732 11172
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 13630 11200 13636 11212
rect 13591 11172 13636 11200
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 10689 11135 10747 11141
rect 10689 11101 10701 11135
rect 10735 11101 10747 11135
rect 10689 11095 10747 11101
rect 13817 11135 13875 11141
rect 13817 11101 13829 11135
rect 13863 11132 13875 11135
rect 13906 11132 13912 11144
rect 13863 11104 13912 11132
rect 13863 11101 13875 11104
rect 13817 11095 13875 11101
rect 13906 11092 13912 11104
rect 13964 11092 13970 11144
rect 13998 11092 14004 11144
rect 14056 11132 14062 11144
rect 14277 11135 14335 11141
rect 14277 11132 14289 11135
rect 14056 11104 14289 11132
rect 14056 11092 14062 11104
rect 14277 11101 14289 11104
rect 14323 11132 14335 11135
rect 15286 11132 15292 11144
rect 14323 11104 15292 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 17494 11092 17500 11144
rect 17552 11132 17558 11144
rect 18064 11141 18092 11240
rect 19242 11228 19248 11240
rect 19300 11268 19306 11280
rect 22094 11268 22100 11280
rect 19300 11240 22100 11268
rect 19300 11228 19306 11240
rect 18316 11203 18374 11209
rect 18316 11169 18328 11203
rect 18362 11200 18374 11203
rect 19058 11200 19064 11212
rect 18362 11172 19064 11200
rect 18362 11169 18374 11172
rect 18316 11163 18374 11169
rect 19058 11160 19064 11172
rect 19116 11160 19122 11212
rect 20916 11209 20944 11240
rect 22094 11228 22100 11240
rect 22152 11228 22158 11280
rect 22830 11228 22836 11280
rect 22888 11268 22894 11280
rect 23937 11271 23995 11277
rect 23937 11268 23949 11271
rect 22888 11240 23949 11268
rect 22888 11228 22894 11240
rect 23937 11237 23949 11240
rect 23983 11268 23995 11271
rect 24670 11268 24676 11280
rect 23983 11240 24676 11268
rect 23983 11237 23995 11240
rect 23937 11231 23995 11237
rect 24670 11228 24676 11240
rect 24728 11268 24734 11280
rect 24946 11268 24952 11280
rect 24728 11240 24952 11268
rect 24728 11228 24734 11240
rect 24946 11228 24952 11240
rect 25004 11228 25010 11280
rect 20901 11203 20959 11209
rect 20901 11169 20913 11203
rect 20947 11169 20959 11203
rect 20901 11163 20959 11169
rect 20990 11160 20996 11212
rect 21048 11200 21054 11212
rect 21157 11203 21215 11209
rect 21157 11200 21169 11203
rect 21048 11172 21169 11200
rect 21048 11160 21054 11172
rect 21157 11169 21169 11172
rect 21203 11169 21215 11203
rect 22112 11200 22140 11228
rect 22278 11200 22284 11212
rect 22112 11172 22284 11200
rect 21157 11163 21215 11169
rect 22278 11160 22284 11172
rect 22336 11160 22342 11212
rect 25038 11200 25044 11212
rect 24999 11172 25044 11200
rect 25038 11160 25044 11172
rect 25096 11160 25102 11212
rect 18049 11135 18107 11141
rect 18049 11132 18061 11135
rect 17552 11104 18061 11132
rect 17552 11092 17558 11104
rect 18049 11101 18061 11104
rect 18095 11101 18107 11135
rect 18049 11095 18107 11101
rect 24026 11092 24032 11144
rect 24084 11132 24090 11144
rect 24578 11132 24584 11144
rect 24084 11104 24177 11132
rect 24539 11104 24584 11132
rect 24084 11092 24090 11104
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 6052 11036 6224 11064
rect 9493 11067 9551 11073
rect 6052 11024 6058 11036
rect 9493 11033 9505 11067
rect 9539 11064 9551 11067
rect 9582 11064 9588 11076
rect 9539 11036 9588 11064
rect 9539 11033 9551 11036
rect 9493 11027 9551 11033
rect 9582 11024 9588 11036
rect 9640 11024 9646 11076
rect 10042 11064 10048 11076
rect 9692 11036 10048 11064
rect 3145 10999 3203 11005
rect 3145 10996 3157 10999
rect 2424 10968 3157 10996
rect 3145 10965 3157 10968
rect 3191 10996 3203 10999
rect 3602 10996 3608 11008
rect 3191 10968 3608 10996
rect 3191 10965 3203 10968
rect 3145 10959 3203 10965
rect 3602 10956 3608 10968
rect 3660 10956 3666 11008
rect 5166 10996 5172 11008
rect 5127 10968 5172 10996
rect 5166 10956 5172 10968
rect 5224 10956 5230 11008
rect 5442 10956 5448 11008
rect 5500 10996 5506 11008
rect 5629 10999 5687 11005
rect 5629 10996 5641 10999
rect 5500 10968 5641 10996
rect 5500 10956 5506 10968
rect 5629 10965 5641 10968
rect 5675 10996 5687 10999
rect 6086 10996 6092 11008
rect 5675 10968 6092 10996
rect 5675 10965 5687 10968
rect 5629 10959 5687 10965
rect 6086 10956 6092 10968
rect 6144 10956 6150 11008
rect 8938 10956 8944 11008
rect 8996 10996 9002 11008
rect 9692 10996 9720 11036
rect 10042 11024 10048 11036
rect 10100 11064 10106 11076
rect 10226 11064 10232 11076
rect 10100 11036 10232 11064
rect 10100 11024 10106 11036
rect 10226 11024 10232 11036
rect 10284 11024 10290 11076
rect 20349 11067 20407 11073
rect 20349 11033 20361 11067
rect 20395 11064 20407 11067
rect 20714 11064 20720 11076
rect 20395 11036 20720 11064
rect 20395 11033 20407 11036
rect 20349 11027 20407 11033
rect 20714 11024 20720 11036
rect 20772 11024 20778 11076
rect 22462 11064 22468 11076
rect 21836 11036 22468 11064
rect 8996 10968 9720 10996
rect 10597 10999 10655 11005
rect 8996 10956 9002 10968
rect 10597 10965 10609 10999
rect 10643 10996 10655 10999
rect 10686 10996 10692 11008
rect 10643 10968 10692 10996
rect 10643 10965 10655 10968
rect 10597 10959 10655 10965
rect 10686 10956 10692 10968
rect 10744 10956 10750 11008
rect 17954 10996 17960 11008
rect 17915 10968 17960 10996
rect 17954 10956 17960 10968
rect 18012 10956 18018 11008
rect 20070 10956 20076 11008
rect 20128 10996 20134 11008
rect 21836 10996 21864 11036
rect 22462 11024 22468 11036
rect 22520 11024 22526 11076
rect 23017 11067 23075 11073
rect 23017 11033 23029 11067
rect 23063 11064 23075 11067
rect 24044 11064 24072 11092
rect 23063 11036 24072 11064
rect 23063 11033 23075 11036
rect 23017 11027 23075 11033
rect 20128 10968 21864 10996
rect 20128 10956 20134 10968
rect 22094 10956 22100 11008
rect 22152 10996 22158 11008
rect 23477 10999 23535 11005
rect 23477 10996 23489 10999
rect 22152 10968 23489 10996
rect 22152 10956 22158 10968
rect 23477 10965 23489 10968
rect 23523 10965 23535 10999
rect 23477 10959 23535 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 2958 10792 2964 10804
rect 1627 10764 2964 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 2958 10752 2964 10764
rect 3016 10752 3022 10804
rect 3973 10795 4031 10801
rect 3973 10761 3985 10795
rect 4019 10792 4031 10795
rect 4614 10792 4620 10804
rect 4019 10764 4620 10792
rect 4019 10761 4031 10764
rect 3973 10755 4031 10761
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 6454 10792 6460 10804
rect 6415 10764 6460 10792
rect 6454 10752 6460 10764
rect 6512 10752 6518 10804
rect 8478 10752 8484 10804
rect 8536 10792 8542 10804
rect 8938 10792 8944 10804
rect 8536 10764 8944 10792
rect 8536 10752 8542 10764
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 13541 10795 13599 10801
rect 13541 10761 13553 10795
rect 13587 10792 13599 10795
rect 13630 10792 13636 10804
rect 13587 10764 13636 10792
rect 13587 10761 13599 10764
rect 13541 10755 13599 10761
rect 13630 10752 13636 10764
rect 13688 10752 13694 10804
rect 13906 10752 13912 10804
rect 13964 10792 13970 10804
rect 14185 10795 14243 10801
rect 14185 10792 14197 10795
rect 13964 10764 14197 10792
rect 13964 10752 13970 10764
rect 14185 10761 14197 10764
rect 14231 10761 14243 10795
rect 16850 10792 16856 10804
rect 16811 10764 16856 10792
rect 14185 10755 14243 10761
rect 16850 10752 16856 10764
rect 16908 10752 16914 10804
rect 18233 10795 18291 10801
rect 18233 10761 18245 10795
rect 18279 10792 18291 10795
rect 18874 10792 18880 10804
rect 18279 10764 18880 10792
rect 18279 10761 18291 10764
rect 18233 10755 18291 10761
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 20622 10792 20628 10804
rect 20583 10764 20628 10792
rect 20622 10752 20628 10764
rect 20680 10752 20686 10804
rect 22649 10795 22707 10801
rect 22649 10761 22661 10795
rect 22695 10792 22707 10795
rect 23290 10792 23296 10804
rect 22695 10764 23296 10792
rect 22695 10761 22707 10764
rect 22649 10755 22707 10761
rect 23290 10752 23296 10764
rect 23348 10752 23354 10804
rect 24670 10792 24676 10804
rect 24631 10764 24676 10792
rect 24670 10752 24676 10764
rect 24728 10752 24734 10804
rect 25038 10792 25044 10804
rect 24999 10764 25044 10792
rect 25038 10752 25044 10764
rect 25096 10752 25102 10804
rect 25409 10795 25467 10801
rect 25409 10761 25421 10795
rect 25455 10792 25467 10795
rect 25498 10792 25504 10804
rect 25455 10764 25504 10792
rect 25455 10761 25467 10764
rect 25409 10755 25467 10761
rect 25498 10752 25504 10764
rect 25556 10752 25562 10804
rect 10321 10727 10379 10733
rect 10321 10693 10333 10727
rect 10367 10724 10379 10727
rect 11790 10724 11796 10736
rect 10367 10696 11796 10724
rect 10367 10693 10379 10696
rect 10321 10687 10379 10693
rect 11790 10684 11796 10696
rect 11848 10684 11854 10736
rect 20533 10727 20591 10733
rect 20533 10693 20545 10727
rect 20579 10724 20591 10727
rect 20579 10696 21312 10724
rect 20579 10693 20591 10696
rect 20533 10687 20591 10693
rect 2038 10656 2044 10668
rect 1412 10628 2044 10656
rect 1412 10597 1440 10628
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10656 5779 10659
rect 5994 10656 6000 10668
rect 5767 10628 6000 10656
rect 5767 10625 5779 10628
rect 5721 10619 5779 10625
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10656 10287 10659
rect 10873 10659 10931 10665
rect 10873 10656 10885 10659
rect 10275 10628 10885 10656
rect 10275 10625 10287 10628
rect 10229 10619 10287 10625
rect 10873 10625 10885 10628
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10557 1455 10591
rect 1397 10551 1455 10557
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10588 2651 10591
rect 3326 10588 3332 10600
rect 2639 10560 3332 10588
rect 2639 10557 2651 10560
rect 2593 10551 2651 10557
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 3602 10548 3608 10600
rect 3660 10588 3666 10600
rect 4985 10591 5043 10597
rect 4985 10588 4997 10591
rect 3660 10560 4997 10588
rect 3660 10548 3666 10560
rect 4985 10557 4997 10560
rect 5031 10588 5043 10591
rect 5445 10591 5503 10597
rect 5445 10588 5457 10591
rect 5031 10560 5457 10588
rect 5031 10557 5043 10560
rect 4985 10551 5043 10557
rect 5445 10557 5457 10560
rect 5491 10588 5503 10591
rect 5534 10588 5540 10600
rect 5491 10560 5540 10588
rect 5491 10557 5503 10560
rect 5445 10551 5503 10557
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 7282 10548 7288 10600
rect 7340 10588 7346 10600
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 7340 10560 7573 10588
rect 7340 10548 7346 10560
rect 7561 10557 7573 10560
rect 7607 10588 7619 10591
rect 7650 10588 7656 10600
rect 7607 10560 7656 10588
rect 7607 10557 7619 10560
rect 7561 10551 7619 10557
rect 7650 10548 7656 10560
rect 7708 10548 7714 10600
rect 7828 10591 7886 10597
rect 7828 10588 7840 10591
rect 7760 10560 7840 10588
rect 2866 10529 2872 10532
rect 2860 10520 2872 10529
rect 2827 10492 2872 10520
rect 2860 10483 2872 10492
rect 2866 10480 2872 10483
rect 2924 10480 2930 10532
rect 2958 10480 2964 10532
rect 3016 10520 3022 10532
rect 3878 10520 3884 10532
rect 3016 10492 3884 10520
rect 3016 10480 3022 10492
rect 3878 10480 3884 10492
rect 3936 10520 3942 10532
rect 7101 10523 7159 10529
rect 3936 10492 5120 10520
rect 3936 10480 3942 10492
rect 2314 10452 2320 10464
rect 2275 10424 2320 10452
rect 2314 10412 2320 10424
rect 2372 10412 2378 10464
rect 5092 10461 5120 10492
rect 7101 10489 7113 10523
rect 7147 10520 7159 10523
rect 7760 10520 7788 10560
rect 7828 10557 7840 10560
rect 7874 10588 7886 10591
rect 8202 10588 8208 10600
rect 7874 10560 8208 10588
rect 7874 10557 7886 10560
rect 7828 10551 7886 10557
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 10689 10591 10747 10597
rect 10689 10588 10701 10591
rect 9732 10560 10701 10588
rect 9732 10548 9738 10560
rect 10689 10557 10701 10560
rect 10735 10557 10747 10591
rect 10888 10588 10916 10619
rect 11698 10616 11704 10668
rect 11756 10656 11762 10668
rect 11885 10659 11943 10665
rect 11885 10656 11897 10659
rect 11756 10628 11897 10656
rect 11756 10616 11762 10628
rect 11885 10625 11897 10628
rect 11931 10656 11943 10659
rect 11977 10659 12035 10665
rect 11977 10656 11989 10659
rect 11931 10628 11989 10656
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 11977 10625 11989 10628
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 12066 10616 12072 10668
rect 12124 10656 12130 10668
rect 12253 10659 12311 10665
rect 12253 10656 12265 10659
rect 12124 10628 12265 10656
rect 12124 10616 12130 10628
rect 12253 10625 12265 10628
rect 12299 10656 12311 10659
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 12299 10628 13001 10656
rect 12299 10625 12311 10628
rect 12253 10619 12311 10625
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 17497 10659 17555 10665
rect 17497 10625 17509 10659
rect 17543 10656 17555 10659
rect 18782 10656 18788 10668
rect 17543 10628 18788 10656
rect 17543 10625 17555 10628
rect 17497 10619 17555 10625
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 21082 10656 21088 10668
rect 21043 10628 21088 10656
rect 21082 10616 21088 10628
rect 21140 10616 21146 10668
rect 21284 10665 21312 10696
rect 21269 10659 21327 10665
rect 21269 10625 21281 10659
rect 21315 10656 21327 10659
rect 21358 10656 21364 10668
rect 21315 10628 21364 10656
rect 21315 10625 21327 10628
rect 21269 10619 21327 10625
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 24302 10656 24308 10668
rect 24215 10628 24308 10656
rect 24302 10616 24308 10628
rect 24360 10656 24366 10668
rect 24854 10656 24860 10668
rect 24360 10628 24860 10656
rect 24360 10616 24366 10628
rect 24854 10616 24860 10628
rect 24912 10616 24918 10668
rect 10962 10588 10968 10600
rect 10875 10560 10968 10588
rect 10689 10551 10747 10557
rect 10962 10548 10968 10560
rect 11020 10588 11026 10600
rect 12618 10588 12624 10600
rect 11020 10560 12624 10588
rect 11020 10548 11026 10560
rect 12618 10548 12624 10560
rect 12676 10548 12682 10600
rect 12805 10591 12863 10597
rect 12805 10557 12817 10591
rect 12851 10588 12863 10591
rect 13078 10588 13084 10600
rect 12851 10560 13084 10588
rect 12851 10557 12863 10560
rect 12805 10551 12863 10557
rect 13078 10548 13084 10560
rect 13136 10548 13142 10600
rect 15013 10591 15071 10597
rect 15013 10557 15025 10591
rect 15059 10588 15071 10591
rect 15286 10588 15292 10600
rect 15059 10560 15292 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 15286 10548 15292 10560
rect 15344 10588 15350 10600
rect 15473 10591 15531 10597
rect 15473 10588 15485 10591
rect 15344 10560 15485 10588
rect 15344 10548 15350 10560
rect 15473 10557 15485 10560
rect 15519 10557 15531 10591
rect 15473 10551 15531 10557
rect 7147 10492 7788 10520
rect 11977 10523 12035 10529
rect 7147 10489 7159 10492
rect 7101 10483 7159 10489
rect 11977 10489 11989 10523
rect 12023 10520 12035 10523
rect 12897 10523 12955 10529
rect 12897 10520 12909 10523
rect 12023 10492 12909 10520
rect 12023 10489 12035 10492
rect 11977 10483 12035 10489
rect 12897 10489 12909 10492
rect 12943 10489 12955 10523
rect 12897 10483 12955 10489
rect 13722 10480 13728 10532
rect 13780 10520 13786 10532
rect 13909 10523 13967 10529
rect 13909 10520 13921 10523
rect 13780 10492 13921 10520
rect 13780 10480 13786 10492
rect 13909 10489 13921 10492
rect 13955 10520 13967 10523
rect 14550 10520 14556 10532
rect 13955 10492 14556 10520
rect 13955 10489 13967 10492
rect 13909 10483 13967 10489
rect 14550 10480 14556 10492
rect 14608 10480 14614 10532
rect 5077 10455 5135 10461
rect 5077 10421 5089 10455
rect 5123 10421 5135 10455
rect 5077 10415 5135 10421
rect 5166 10412 5172 10464
rect 5224 10452 5230 10464
rect 5537 10455 5595 10461
rect 5537 10452 5549 10455
rect 5224 10424 5549 10452
rect 5224 10412 5230 10424
rect 5537 10421 5549 10424
rect 5583 10421 5595 10455
rect 6178 10452 6184 10464
rect 6139 10424 6184 10452
rect 5537 10415 5595 10421
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 7469 10455 7527 10461
rect 7469 10421 7481 10455
rect 7515 10452 7527 10455
rect 7650 10452 7656 10464
rect 7515 10424 7656 10452
rect 7515 10421 7527 10424
rect 7469 10415 7527 10421
rect 7650 10412 7656 10424
rect 7708 10412 7714 10464
rect 9582 10452 9588 10464
rect 9543 10424 9588 10452
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 10686 10452 10692 10464
rect 9824 10424 10692 10452
rect 9824 10412 9830 10424
rect 10686 10412 10692 10424
rect 10744 10452 10750 10464
rect 10781 10455 10839 10461
rect 10781 10452 10793 10455
rect 10744 10424 10793 10452
rect 10744 10412 10750 10424
rect 10781 10421 10793 10424
rect 10827 10421 10839 10455
rect 10781 10415 10839 10421
rect 11238 10412 11244 10464
rect 11296 10452 11302 10464
rect 11333 10455 11391 10461
rect 11333 10452 11345 10455
rect 11296 10424 11345 10452
rect 11296 10412 11302 10424
rect 11333 10421 11345 10424
rect 11379 10421 11391 10455
rect 11333 10415 11391 10421
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 13630 10452 13636 10464
rect 12483 10424 13636 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 14458 10452 14464 10464
rect 14419 10424 14464 10452
rect 14458 10412 14464 10424
rect 14516 10412 14522 10464
rect 15381 10455 15439 10461
rect 15381 10421 15393 10455
rect 15427 10452 15439 10455
rect 15488 10452 15516 10551
rect 15562 10548 15568 10600
rect 15620 10588 15626 10600
rect 15740 10591 15798 10597
rect 15740 10588 15752 10591
rect 15620 10560 15752 10588
rect 15620 10548 15626 10560
rect 15740 10557 15752 10560
rect 15786 10588 15798 10591
rect 16482 10588 16488 10600
rect 15786 10560 16488 10588
rect 15786 10557 15798 10560
rect 15740 10551 15798 10557
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 20714 10548 20720 10600
rect 20772 10588 20778 10600
rect 20993 10591 21051 10597
rect 20993 10588 21005 10591
rect 20772 10560 21005 10588
rect 20772 10548 20778 10560
rect 20993 10557 21005 10560
rect 21039 10557 21051 10591
rect 22462 10588 22468 10600
rect 22423 10560 22468 10588
rect 20993 10551 21051 10557
rect 22462 10548 22468 10560
rect 22520 10588 22526 10600
rect 23017 10591 23075 10597
rect 23017 10588 23029 10591
rect 22520 10560 23029 10588
rect 22520 10548 22526 10560
rect 23017 10557 23029 10560
rect 23063 10557 23075 10591
rect 23017 10551 23075 10557
rect 23106 10548 23112 10600
rect 23164 10588 23170 10600
rect 24029 10591 24087 10597
rect 24029 10588 24041 10591
rect 23164 10560 24041 10588
rect 23164 10548 23170 10560
rect 24029 10557 24041 10560
rect 24075 10557 24087 10591
rect 25222 10588 25228 10600
rect 25183 10560 25228 10588
rect 24029 10551 24087 10557
rect 25222 10548 25228 10560
rect 25280 10588 25286 10600
rect 25777 10591 25835 10597
rect 25777 10588 25789 10591
rect 25280 10560 25789 10588
rect 25280 10548 25286 10560
rect 25777 10557 25789 10560
rect 25823 10557 25835 10591
rect 25777 10551 25835 10557
rect 17954 10480 17960 10532
rect 18012 10520 18018 10532
rect 18601 10523 18659 10529
rect 18601 10520 18613 10523
rect 18012 10492 18613 10520
rect 18012 10480 18018 10492
rect 18601 10489 18613 10492
rect 18647 10489 18659 10523
rect 19613 10523 19671 10529
rect 19613 10520 19625 10523
rect 18601 10483 18659 10489
rect 18708 10492 19625 10520
rect 18708 10464 18736 10492
rect 19613 10489 19625 10492
rect 19659 10489 19671 10523
rect 19613 10483 19671 10489
rect 21729 10523 21787 10529
rect 21729 10489 21741 10523
rect 21775 10520 21787 10523
rect 22278 10520 22284 10532
rect 21775 10492 22284 10520
rect 21775 10489 21787 10492
rect 21729 10483 21787 10489
rect 22278 10480 22284 10492
rect 22336 10480 22342 10532
rect 23477 10523 23535 10529
rect 23477 10489 23489 10523
rect 23523 10520 23535 10523
rect 23750 10520 23756 10532
rect 23523 10492 23756 10520
rect 23523 10489 23535 10492
rect 23477 10483 23535 10489
rect 23750 10480 23756 10492
rect 23808 10520 23814 10532
rect 24118 10520 24124 10532
rect 23808 10492 24124 10520
rect 23808 10480 23814 10492
rect 24118 10480 24124 10492
rect 24176 10480 24182 10532
rect 17494 10452 17500 10464
rect 15427 10424 17500 10452
rect 15427 10421 15439 10424
rect 15381 10415 15439 10421
rect 17494 10412 17500 10424
rect 17552 10452 17558 10464
rect 17773 10455 17831 10461
rect 17773 10452 17785 10455
rect 17552 10424 17785 10452
rect 17552 10412 17558 10424
rect 17773 10421 17785 10424
rect 17819 10421 17831 10455
rect 18690 10452 18696 10464
rect 18651 10424 18696 10452
rect 17773 10415 17831 10421
rect 18690 10412 18696 10424
rect 18748 10412 18754 10464
rect 19058 10412 19064 10464
rect 19116 10452 19122 10464
rect 19337 10455 19395 10461
rect 19337 10452 19349 10455
rect 19116 10424 19349 10452
rect 19116 10412 19122 10424
rect 19337 10421 19349 10424
rect 19383 10452 19395 10455
rect 19426 10452 19432 10464
rect 19383 10424 19432 10452
rect 19383 10421 19395 10424
rect 19337 10415 19395 10421
rect 19426 10412 19432 10424
rect 19484 10412 19490 10464
rect 20165 10455 20223 10461
rect 20165 10421 20177 10455
rect 20211 10452 20223 10455
rect 20346 10452 20352 10464
rect 20211 10424 20352 10452
rect 20211 10421 20223 10424
rect 20165 10415 20223 10421
rect 20346 10412 20352 10424
rect 20404 10412 20410 10464
rect 22373 10455 22431 10461
rect 22373 10421 22385 10455
rect 22419 10452 22431 10455
rect 22554 10452 22560 10464
rect 22419 10424 22560 10452
rect 22419 10421 22431 10424
rect 22373 10415 22431 10421
rect 22554 10412 22560 10424
rect 22612 10412 22618 10464
rect 23658 10452 23664 10464
rect 23619 10424 23664 10452
rect 23658 10412 23664 10424
rect 23716 10412 23722 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2406 10248 2412 10260
rect 2367 10220 2412 10248
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 7558 10248 7564 10260
rect 7519 10220 7564 10248
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 8662 10248 8668 10260
rect 8623 10220 8668 10248
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 9306 10248 9312 10260
rect 9267 10220 9312 10248
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 11146 10248 11152 10260
rect 11107 10220 11152 10248
rect 11146 10208 11152 10220
rect 11204 10208 11210 10260
rect 11609 10251 11667 10257
rect 11609 10217 11621 10251
rect 11655 10248 11667 10251
rect 11790 10248 11796 10260
rect 11655 10220 11796 10248
rect 11655 10217 11667 10220
rect 11609 10211 11667 10217
rect 11790 10208 11796 10220
rect 11848 10208 11854 10260
rect 14458 10248 14464 10260
rect 14419 10220 14464 10248
rect 14458 10208 14464 10220
rect 14516 10208 14522 10260
rect 15105 10251 15163 10257
rect 15105 10217 15117 10251
rect 15151 10248 15163 10251
rect 15562 10248 15568 10260
rect 15151 10220 15568 10248
rect 15151 10217 15163 10220
rect 15105 10211 15163 10217
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18141 10251 18199 10257
rect 18141 10248 18153 10251
rect 18012 10220 18153 10248
rect 18012 10208 18018 10220
rect 18141 10217 18153 10220
rect 18187 10217 18199 10251
rect 18141 10211 18199 10217
rect 20438 10208 20444 10260
rect 20496 10248 20502 10260
rect 20533 10251 20591 10257
rect 20533 10248 20545 10251
rect 20496 10220 20545 10248
rect 20496 10208 20502 10220
rect 20533 10217 20545 10220
rect 20579 10217 20591 10251
rect 20533 10211 20591 10217
rect 20714 10208 20720 10260
rect 20772 10248 20778 10260
rect 20901 10251 20959 10257
rect 20901 10248 20913 10251
rect 20772 10220 20913 10248
rect 20772 10208 20778 10220
rect 20901 10217 20913 10220
rect 20947 10217 20959 10251
rect 21266 10248 21272 10260
rect 21227 10220 21272 10248
rect 20901 10211 20959 10217
rect 21266 10208 21272 10220
rect 21324 10208 21330 10260
rect 21358 10208 21364 10260
rect 21416 10248 21422 10260
rect 21910 10248 21916 10260
rect 21416 10220 21916 10248
rect 21416 10208 21422 10220
rect 21910 10208 21916 10220
rect 21968 10208 21974 10260
rect 22094 10208 22100 10260
rect 22152 10248 22158 10260
rect 23106 10248 23112 10260
rect 22152 10220 22197 10248
rect 23067 10220 23112 10248
rect 22152 10208 22158 10220
rect 23106 10208 23112 10220
rect 23164 10208 23170 10260
rect 2317 10183 2375 10189
rect 2317 10149 2329 10183
rect 2363 10180 2375 10183
rect 2866 10180 2872 10192
rect 2363 10152 2872 10180
rect 2363 10149 2375 10152
rect 2317 10143 2375 10149
rect 2866 10140 2872 10152
rect 2924 10180 2930 10192
rect 5350 10180 5356 10192
rect 2924 10152 3096 10180
rect 2924 10140 2930 10152
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 1443 10084 1532 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 1504 9988 1532 10084
rect 2774 10072 2780 10124
rect 2832 10112 2838 10124
rect 2832 10084 2877 10112
rect 2832 10072 2838 10084
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10044 2927 10047
rect 2958 10044 2964 10056
rect 2915 10016 2964 10044
rect 2915 10013 2927 10016
rect 2869 10007 2927 10013
rect 2958 10004 2964 10016
rect 3016 10004 3022 10056
rect 3068 10053 3096 10152
rect 4540 10152 5356 10180
rect 3326 10072 3332 10124
rect 3384 10112 3390 10124
rect 4540 10121 4568 10152
rect 5350 10140 5356 10152
rect 5408 10140 5414 10192
rect 6178 10140 6184 10192
rect 6236 10180 6242 10192
rect 8938 10180 8944 10192
rect 6236 10152 8064 10180
rect 8899 10152 8944 10180
rect 6236 10140 6242 10152
rect 3513 10115 3571 10121
rect 3513 10112 3525 10115
rect 3384 10084 3525 10112
rect 3384 10072 3390 10084
rect 3513 10081 3525 10084
rect 3559 10112 3571 10115
rect 4525 10115 4583 10121
rect 4525 10112 4537 10115
rect 3559 10084 4537 10112
rect 3559 10081 3571 10084
rect 3513 10075 3571 10081
rect 4525 10081 4537 10084
rect 4571 10081 4583 10115
rect 4525 10075 4583 10081
rect 4792 10115 4850 10121
rect 4792 10081 4804 10115
rect 4838 10112 4850 10115
rect 5994 10112 6000 10124
rect 4838 10084 6000 10112
rect 4838 10081 4850 10084
rect 4792 10075 4850 10081
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 7558 10072 7564 10124
rect 7616 10112 7622 10124
rect 8036 10121 8064 10152
rect 8938 10140 8944 10152
rect 8996 10140 9002 10192
rect 9858 10140 9864 10192
rect 9916 10180 9922 10192
rect 13173 10183 13231 10189
rect 13173 10180 13185 10183
rect 9916 10152 13185 10180
rect 9916 10140 9922 10152
rect 13173 10149 13185 10152
rect 13219 10149 13231 10183
rect 13173 10143 13231 10149
rect 15286 10140 15292 10192
rect 15344 10180 15350 10192
rect 15749 10183 15807 10189
rect 15749 10180 15761 10183
rect 15344 10152 15761 10180
rect 15344 10140 15350 10152
rect 15749 10149 15761 10152
rect 15795 10149 15807 10183
rect 18046 10180 18052 10192
rect 18007 10152 18052 10180
rect 15749 10143 15807 10149
rect 18046 10140 18052 10152
rect 18104 10180 18110 10192
rect 18509 10183 18567 10189
rect 18509 10180 18521 10183
rect 18104 10152 18521 10180
rect 18104 10140 18110 10152
rect 18509 10149 18521 10152
rect 18555 10149 18567 10183
rect 18509 10143 18567 10149
rect 22833 10183 22891 10189
rect 22833 10149 22845 10183
rect 22879 10180 22891 10183
rect 23658 10180 23664 10192
rect 22879 10152 23664 10180
rect 22879 10149 22891 10152
rect 22833 10143 22891 10149
rect 23658 10140 23664 10152
rect 23716 10140 23722 10192
rect 7929 10115 7987 10121
rect 7929 10112 7941 10115
rect 7616 10084 7941 10112
rect 7616 10072 7622 10084
rect 7929 10081 7941 10084
rect 7975 10081 7987 10115
rect 7929 10075 7987 10081
rect 8021 10115 8079 10121
rect 8021 10081 8033 10115
rect 8067 10112 8079 10115
rect 8386 10112 8392 10124
rect 8067 10084 8392 10112
rect 8067 10081 8079 10084
rect 8021 10075 8079 10081
rect 8386 10072 8392 10084
rect 8444 10072 8450 10124
rect 11054 10112 11060 10124
rect 11015 10084 11060 10112
rect 11054 10072 11060 10084
rect 11112 10072 11118 10124
rect 11517 10115 11575 10121
rect 11517 10081 11529 10115
rect 11563 10112 11575 10115
rect 12342 10112 12348 10124
rect 11563 10084 12348 10112
rect 11563 10081 11575 10084
rect 11517 10075 11575 10081
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 12894 10112 12900 10124
rect 12728 10084 12900 10112
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10044 3111 10047
rect 8202 10044 8208 10056
rect 3099 10016 4476 10044
rect 8163 10016 8208 10044
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 1486 9936 1492 9988
rect 1544 9976 1550 9988
rect 1857 9979 1915 9985
rect 1857 9976 1869 9979
rect 1544 9948 1869 9976
rect 1544 9936 1550 9948
rect 1857 9945 1869 9948
rect 1903 9945 1915 9979
rect 1857 9939 1915 9945
rect 2590 9936 2596 9988
rect 2648 9976 2654 9988
rect 3789 9979 3847 9985
rect 3789 9976 3801 9979
rect 2648 9948 3801 9976
rect 2648 9936 2654 9948
rect 3789 9945 3801 9948
rect 3835 9945 3847 9979
rect 3789 9939 3847 9945
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 1762 9908 1768 9920
rect 1627 9880 1768 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 1762 9868 1768 9880
rect 1820 9868 1826 9920
rect 4448 9917 4476 10016
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 10134 10044 10140 10056
rect 10095 10016 10140 10044
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 11606 10004 11612 10056
rect 11664 10044 11670 10056
rect 11701 10047 11759 10053
rect 11701 10044 11713 10047
rect 11664 10016 11713 10044
rect 11664 10004 11670 10016
rect 11701 10013 11713 10016
rect 11747 10013 11759 10047
rect 11701 10007 11759 10013
rect 7469 9979 7527 9985
rect 7469 9945 7481 9979
rect 7515 9976 7527 9979
rect 7742 9976 7748 9988
rect 7515 9948 7748 9976
rect 7515 9945 7527 9948
rect 7469 9939 7527 9945
rect 7742 9936 7748 9948
rect 7800 9976 7806 9988
rect 8220 9976 8248 10004
rect 12728 9985 12756 10084
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 13078 10112 13084 10124
rect 13039 10084 13084 10112
rect 13078 10072 13084 10084
rect 13136 10072 13142 10124
rect 15657 10115 15715 10121
rect 15657 10081 15669 10115
rect 15703 10112 15715 10115
rect 15930 10112 15936 10124
rect 15703 10084 15936 10112
rect 15703 10081 15715 10084
rect 15657 10075 15715 10081
rect 15930 10072 15936 10084
rect 15988 10072 15994 10124
rect 17770 10072 17776 10124
rect 17828 10112 17834 10124
rect 18601 10115 18659 10121
rect 18601 10112 18613 10115
rect 17828 10084 18613 10112
rect 17828 10072 17834 10084
rect 18601 10081 18613 10084
rect 18647 10081 18659 10115
rect 18601 10075 18659 10081
rect 19334 10072 19340 10124
rect 19392 10112 19398 10124
rect 19797 10115 19855 10121
rect 19797 10112 19809 10115
rect 19392 10084 19809 10112
rect 19392 10072 19398 10084
rect 19797 10081 19809 10084
rect 19843 10112 19855 10115
rect 19886 10112 19892 10124
rect 19843 10084 19892 10112
rect 19843 10081 19855 10084
rect 19797 10075 19855 10081
rect 19886 10072 19892 10084
rect 19944 10072 19950 10124
rect 22554 10072 22560 10124
rect 22612 10112 22618 10124
rect 23106 10112 23112 10124
rect 22612 10084 23112 10112
rect 22612 10072 22618 10084
rect 23106 10072 23112 10084
rect 23164 10112 23170 10124
rect 23560 10115 23618 10121
rect 23560 10112 23572 10115
rect 23164 10084 23572 10112
rect 23164 10072 23170 10084
rect 23560 10081 23572 10084
rect 23606 10112 23618 10115
rect 24302 10112 24308 10124
rect 23606 10084 24308 10112
rect 23606 10081 23618 10084
rect 23560 10075 23618 10081
rect 24302 10072 24308 10084
rect 24360 10072 24366 10124
rect 13262 10044 13268 10056
rect 13223 10016 13268 10044
rect 13262 10004 13268 10016
rect 13320 10004 13326 10056
rect 15378 10004 15384 10056
rect 15436 10044 15442 10056
rect 15841 10047 15899 10053
rect 15841 10044 15853 10047
rect 15436 10016 15853 10044
rect 15436 10004 15442 10016
rect 15841 10013 15853 10016
rect 15887 10013 15899 10047
rect 16666 10044 16672 10056
rect 16627 10016 16672 10044
rect 15841 10007 15899 10013
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 17129 10047 17187 10053
rect 17129 10013 17141 10047
rect 17175 10044 17187 10047
rect 18138 10044 18144 10056
rect 17175 10016 18144 10044
rect 17175 10013 17187 10016
rect 17129 10007 17187 10013
rect 18138 10004 18144 10016
rect 18196 10004 18202 10056
rect 18693 10047 18751 10053
rect 18693 10013 18705 10047
rect 18739 10013 18751 10047
rect 18693 10007 18751 10013
rect 21453 10047 21511 10053
rect 21453 10013 21465 10047
rect 21499 10013 21511 10047
rect 21453 10007 21511 10013
rect 7800 9948 8248 9976
rect 12713 9979 12771 9985
rect 7800 9936 7806 9948
rect 12713 9945 12725 9979
rect 12759 9945 12771 9979
rect 12713 9939 12771 9945
rect 14826 9936 14832 9988
rect 14884 9976 14890 9988
rect 15289 9979 15347 9985
rect 15289 9976 15301 9979
rect 14884 9948 15301 9976
rect 14884 9936 14890 9948
rect 15289 9945 15301 9948
rect 15335 9945 15347 9979
rect 18708 9976 18736 10007
rect 19426 9976 19432 9988
rect 15289 9939 15347 9945
rect 17604 9948 19432 9976
rect 17604 9920 17632 9948
rect 19426 9936 19432 9948
rect 19484 9936 19490 9988
rect 19978 9976 19984 9988
rect 19939 9948 19984 9976
rect 19978 9936 19984 9948
rect 20036 9936 20042 9988
rect 20346 9936 20352 9988
rect 20404 9976 20410 9988
rect 20990 9976 20996 9988
rect 20404 9948 20996 9976
rect 20404 9936 20410 9948
rect 20990 9936 20996 9948
rect 21048 9976 21054 9988
rect 21468 9976 21496 10007
rect 22278 10004 22284 10056
rect 22336 10044 22342 10056
rect 22830 10044 22836 10056
rect 22336 10016 22836 10044
rect 22336 10004 22342 10016
rect 22830 10004 22836 10016
rect 22888 10044 22894 10056
rect 23293 10047 23351 10053
rect 23293 10044 23305 10047
rect 22888 10016 23305 10044
rect 22888 10004 22894 10016
rect 23293 10013 23305 10016
rect 23339 10013 23351 10047
rect 23293 10007 23351 10013
rect 21048 9948 21496 9976
rect 21048 9936 21054 9948
rect 4433 9911 4491 9917
rect 4433 9877 4445 9911
rect 4479 9908 4491 9911
rect 5166 9908 5172 9920
rect 4479 9880 5172 9908
rect 4479 9877 4491 9880
rect 4433 9871 4491 9877
rect 5166 9868 5172 9880
rect 5224 9908 5230 9920
rect 5905 9911 5963 9917
rect 5905 9908 5917 9911
rect 5224 9880 5917 9908
rect 5224 9868 5230 9880
rect 5905 9877 5917 9880
rect 5951 9877 5963 9911
rect 5905 9871 5963 9877
rect 5994 9868 6000 9920
rect 6052 9908 6058 9920
rect 6457 9911 6515 9917
rect 6457 9908 6469 9911
rect 6052 9880 6469 9908
rect 6052 9868 6058 9880
rect 6457 9877 6469 9880
rect 6503 9877 6515 9911
rect 6914 9908 6920 9920
rect 6875 9880 6920 9908
rect 6457 9871 6515 9877
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 9858 9868 9864 9920
rect 9916 9908 9922 9920
rect 9953 9911 10011 9917
rect 9953 9908 9965 9911
rect 9916 9880 9965 9908
rect 9916 9868 9922 9880
rect 9953 9877 9965 9880
rect 9999 9877 10011 9911
rect 10686 9908 10692 9920
rect 10647 9880 10692 9908
rect 9953 9871 10011 9877
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 12529 9911 12587 9917
rect 12529 9877 12541 9911
rect 12575 9908 12587 9911
rect 12618 9908 12624 9920
rect 12575 9880 12624 9908
rect 12575 9877 12587 9880
rect 12529 9871 12587 9877
rect 12618 9868 12624 9880
rect 12676 9908 12682 9920
rect 12986 9908 12992 9920
rect 12676 9880 12992 9908
rect 12676 9868 12682 9880
rect 12986 9868 12992 9880
rect 13044 9868 13050 9920
rect 13817 9911 13875 9917
rect 13817 9877 13829 9911
rect 13863 9908 13875 9911
rect 13906 9908 13912 9920
rect 13863 9880 13912 9908
rect 13863 9877 13875 9880
rect 13817 9871 13875 9877
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 13998 9868 14004 9920
rect 14056 9908 14062 9920
rect 14093 9911 14151 9917
rect 14093 9908 14105 9911
rect 14056 9880 14105 9908
rect 14056 9868 14062 9880
rect 14093 9877 14105 9880
rect 14139 9877 14151 9911
rect 16390 9908 16396 9920
rect 16351 9880 16396 9908
rect 14093 9871 14151 9877
rect 16390 9868 16396 9880
rect 16448 9868 16454 9920
rect 17586 9908 17592 9920
rect 17547 9880 17592 9908
rect 17586 9868 17592 9880
rect 17644 9868 17650 9920
rect 24673 9911 24731 9917
rect 24673 9877 24685 9911
rect 24719 9908 24731 9911
rect 24762 9908 24768 9920
rect 24719 9880 24768 9908
rect 24719 9877 24731 9880
rect 24673 9871 24731 9877
rect 24762 9868 24768 9880
rect 24820 9868 24826 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 8662 9664 8668 9716
rect 8720 9704 8726 9716
rect 9309 9707 9367 9713
rect 9309 9704 9321 9707
rect 8720 9676 9321 9704
rect 8720 9664 8726 9676
rect 9309 9673 9321 9676
rect 9355 9673 9367 9707
rect 9309 9667 9367 9673
rect 10594 9664 10600 9716
rect 10652 9704 10658 9716
rect 10870 9704 10876 9716
rect 10652 9676 10876 9704
rect 10652 9664 10658 9676
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 13262 9664 13268 9716
rect 13320 9704 13326 9716
rect 13449 9707 13507 9713
rect 13449 9704 13461 9707
rect 13320 9676 13461 9704
rect 13320 9664 13326 9676
rect 13449 9673 13461 9676
rect 13495 9673 13507 9707
rect 19426 9704 19432 9716
rect 19387 9676 19432 9704
rect 13449 9667 13507 9673
rect 19426 9664 19432 9676
rect 19484 9664 19490 9716
rect 19886 9664 19892 9716
rect 19944 9704 19950 9716
rect 19981 9707 20039 9713
rect 19981 9704 19993 9707
rect 19944 9676 19993 9704
rect 19944 9664 19950 9676
rect 19981 9673 19993 9676
rect 20027 9673 20039 9707
rect 20346 9704 20352 9716
rect 20307 9676 20352 9704
rect 19981 9667 20039 9673
rect 20346 9664 20352 9676
rect 20404 9664 20410 9716
rect 21266 9664 21272 9716
rect 21324 9704 21330 9716
rect 21453 9707 21511 9713
rect 21453 9704 21465 9707
rect 21324 9676 21465 9704
rect 21324 9664 21330 9676
rect 21453 9673 21465 9676
rect 21499 9673 21511 9707
rect 21453 9667 21511 9673
rect 22002 9664 22008 9716
rect 22060 9704 22066 9716
rect 22646 9704 22652 9716
rect 22060 9676 22652 9704
rect 22060 9664 22066 9676
rect 22646 9664 22652 9676
rect 22704 9664 22710 9716
rect 22830 9664 22836 9716
rect 22888 9704 22894 9716
rect 23293 9707 23351 9713
rect 23293 9704 23305 9707
rect 22888 9676 23305 9704
rect 22888 9664 22894 9676
rect 23293 9673 23305 9676
rect 23339 9673 23351 9707
rect 23293 9667 23351 9673
rect 1578 9636 1584 9648
rect 1539 9608 1584 9636
rect 1578 9596 1584 9608
rect 1636 9596 1642 9648
rect 2409 9639 2467 9645
rect 2409 9605 2421 9639
rect 2455 9636 2467 9639
rect 2590 9636 2596 9648
rect 2455 9608 2596 9636
rect 2455 9605 2467 9608
rect 2409 9599 2467 9605
rect 2590 9596 2596 9608
rect 2648 9596 2654 9648
rect 2777 9639 2835 9645
rect 2777 9605 2789 9639
rect 2823 9636 2835 9639
rect 4062 9636 4068 9648
rect 2823 9608 4068 9636
rect 2823 9605 2835 9608
rect 2777 9599 2835 9605
rect 4062 9596 4068 9608
rect 4120 9596 4126 9648
rect 4338 9636 4344 9648
rect 4299 9608 4344 9636
rect 4338 9596 4344 9608
rect 4396 9596 4402 9648
rect 10505 9639 10563 9645
rect 10505 9605 10517 9639
rect 10551 9636 10563 9639
rect 11146 9636 11152 9648
rect 10551 9608 11152 9636
rect 10551 9605 10563 9608
rect 10505 9599 10563 9605
rect 11146 9596 11152 9608
rect 11204 9596 11210 9648
rect 12158 9636 12164 9648
rect 12119 9608 12164 9636
rect 12158 9596 12164 9608
rect 12216 9596 12222 9648
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 12894 9636 12900 9648
rect 12492 9608 12900 9636
rect 12492 9596 12498 9608
rect 12894 9596 12900 9608
rect 12952 9596 12958 9648
rect 14274 9636 14280 9648
rect 14235 9608 14280 9636
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 17126 9636 17132 9648
rect 16684 9608 17132 9636
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5166 9568 5172 9580
rect 5031 9540 5172 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1578 9500 1584 9512
rect 1443 9472 1584 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1578 9460 1584 9472
rect 1636 9500 1642 9512
rect 2409 9503 2467 9509
rect 2409 9500 2421 9503
rect 1636 9472 2421 9500
rect 1636 9460 1642 9472
rect 2409 9469 2421 9472
rect 2455 9469 2467 9503
rect 2409 9463 2467 9469
rect 2501 9503 2559 9509
rect 2501 9469 2513 9503
rect 2547 9500 2559 9503
rect 3145 9503 3203 9509
rect 3145 9500 3157 9503
rect 2547 9472 3157 9500
rect 2547 9469 2559 9472
rect 2501 9463 2559 9469
rect 3145 9469 3157 9472
rect 3191 9469 3203 9503
rect 3145 9463 3203 9469
rect 1854 9392 1860 9444
rect 1912 9432 1918 9444
rect 2317 9435 2375 9441
rect 2317 9432 2329 9435
rect 1912 9404 2329 9432
rect 1912 9392 1918 9404
rect 2317 9401 2329 9404
rect 2363 9432 2375 9435
rect 2363 9404 2912 9432
rect 2363 9401 2375 9404
rect 2317 9395 2375 9401
rect 1302 9324 1308 9376
rect 1360 9364 1366 9376
rect 2501 9367 2559 9373
rect 2501 9364 2513 9367
rect 1360 9336 2513 9364
rect 1360 9324 1366 9336
rect 2501 9333 2513 9336
rect 2547 9364 2559 9367
rect 2593 9367 2651 9373
rect 2593 9364 2605 9367
rect 2547 9336 2605 9364
rect 2547 9333 2559 9336
rect 2501 9327 2559 9333
rect 2593 9333 2605 9336
rect 2639 9333 2651 9367
rect 2884 9364 2912 9404
rect 2958 9392 2964 9444
rect 3016 9432 3022 9444
rect 3436 9432 3464 9531
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 6687 9540 8064 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 4801 9503 4859 9509
rect 4801 9469 4813 9503
rect 4847 9500 4859 9503
rect 5442 9500 5448 9512
rect 4847 9472 5448 9500
rect 4847 9469 4859 9472
rect 4801 9463 4859 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 7929 9503 7987 9509
rect 7929 9500 7941 9503
rect 7708 9472 7941 9500
rect 7708 9460 7714 9472
rect 7929 9469 7941 9472
rect 7975 9469 7987 9503
rect 8036 9500 8064 9540
rect 10686 9528 10692 9580
rect 10744 9568 10750 9580
rect 10870 9568 10876 9580
rect 10744 9540 10876 9568
rect 10744 9528 10750 9540
rect 10870 9528 10876 9540
rect 10928 9568 10934 9580
rect 11057 9571 11115 9577
rect 11057 9568 11069 9571
rect 10928 9540 11069 9568
rect 10928 9528 10934 9540
rect 11057 9537 11069 9540
rect 11103 9537 11115 9571
rect 12176 9568 12204 9596
rect 16684 9580 16712 9608
rect 17126 9596 17132 9608
rect 17184 9596 17190 9648
rect 17494 9636 17500 9648
rect 17455 9608 17500 9636
rect 17494 9596 17500 9608
rect 17552 9596 17558 9648
rect 17770 9636 17776 9648
rect 17731 9608 17776 9636
rect 17770 9596 17776 9608
rect 17828 9596 17834 9648
rect 20717 9639 20775 9645
rect 20717 9605 20729 9639
rect 20763 9636 20775 9639
rect 21818 9636 21824 9648
rect 20763 9608 21824 9636
rect 20763 9605 20775 9608
rect 20717 9599 20775 9605
rect 21818 9596 21824 9608
rect 21876 9596 21882 9648
rect 22094 9596 22100 9648
rect 22152 9636 22158 9648
rect 22152 9608 22508 9636
rect 22152 9596 22158 9608
rect 12176 9540 12940 9568
rect 11057 9531 11115 9537
rect 12912 9512 12940 9540
rect 12986 9528 12992 9580
rect 13044 9568 13050 9580
rect 13044 9540 13089 9568
rect 13044 9528 13050 9540
rect 13262 9528 13268 9580
rect 13320 9528 13326 9580
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9568 14059 9571
rect 15010 9568 15016 9580
rect 14047 9540 15016 9568
rect 14047 9537 14059 9540
rect 14001 9531 14059 9537
rect 15010 9528 15016 9540
rect 15068 9528 15074 9580
rect 16666 9568 16672 9580
rect 16579 9540 16672 9568
rect 16666 9528 16672 9540
rect 16724 9528 16730 9580
rect 17512 9568 17540 9596
rect 18049 9571 18107 9577
rect 18049 9568 18061 9571
rect 17512 9540 18061 9568
rect 8196 9503 8254 9509
rect 8196 9500 8208 9503
rect 8036 9472 8208 9500
rect 7929 9463 7987 9469
rect 8196 9469 8208 9472
rect 8242 9500 8254 9503
rect 8478 9500 8484 9512
rect 8242 9472 8484 9500
rect 8242 9469 8254 9472
rect 8196 9463 8254 9469
rect 3789 9435 3847 9441
rect 3789 9432 3801 9435
rect 3016 9404 3801 9432
rect 3016 9392 3022 9404
rect 3789 9401 3801 9404
rect 3835 9401 3847 9435
rect 3789 9395 3847 9401
rect 4249 9435 4307 9441
rect 4249 9401 4261 9435
rect 4295 9432 4307 9435
rect 4709 9435 4767 9441
rect 4709 9432 4721 9435
rect 4295 9404 4721 9432
rect 4295 9401 4307 9404
rect 4249 9395 4307 9401
rect 4709 9401 4721 9404
rect 4755 9432 4767 9435
rect 6825 9435 6883 9441
rect 6825 9432 6837 9435
rect 4755 9404 6837 9432
rect 4755 9401 4767 9404
rect 4709 9395 4767 9401
rect 6825 9401 6837 9404
rect 6871 9401 6883 9435
rect 7944 9432 7972 9463
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 12434 9460 12440 9512
rect 12492 9500 12498 9512
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 12492 9472 12817 9500
rect 12492 9460 12498 9472
rect 12805 9469 12817 9472
rect 12851 9469 12863 9503
rect 12805 9463 12863 9469
rect 12894 9460 12900 9512
rect 12952 9500 12958 9512
rect 12952 9472 12997 9500
rect 12952 9460 12958 9472
rect 13280 9444 13308 9528
rect 17788 9512 17816 9540
rect 18049 9537 18061 9540
rect 18095 9537 18107 9571
rect 18049 9531 18107 9537
rect 21177 9571 21235 9577
rect 21177 9537 21189 9571
rect 21223 9568 21235 9571
rect 21358 9568 21364 9580
rect 21223 9540 21364 9568
rect 21223 9537 21235 9540
rect 21177 9531 21235 9537
rect 21358 9528 21364 9540
rect 21416 9528 21422 9580
rect 22480 9577 22508 9608
rect 23474 9596 23480 9648
rect 23532 9636 23538 9648
rect 23661 9639 23719 9645
rect 23661 9636 23673 9639
rect 23532 9608 23673 9636
rect 23532 9596 23538 9608
rect 23661 9605 23673 9608
rect 23707 9605 23719 9639
rect 25406 9636 25412 9648
rect 25367 9608 25412 9636
rect 23661 9599 23719 9605
rect 25406 9596 25412 9608
rect 25464 9596 25470 9648
rect 22465 9571 22523 9577
rect 22465 9537 22477 9571
rect 22511 9537 22523 9571
rect 22465 9531 22523 9537
rect 22649 9571 22707 9577
rect 22649 9537 22661 9571
rect 22695 9568 22707 9571
rect 23106 9568 23112 9580
rect 22695 9540 23112 9568
rect 22695 9537 22707 9540
rect 22649 9531 22707 9537
rect 23106 9528 23112 9540
rect 23164 9528 23170 9580
rect 24305 9571 24363 9577
rect 24305 9537 24317 9571
rect 24351 9537 24363 9571
rect 24305 9531 24363 9537
rect 14458 9460 14464 9512
rect 14516 9500 14522 9512
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 14516 9472 14841 9500
rect 14516 9460 14522 9472
rect 14829 9469 14841 9472
rect 14875 9469 14887 9503
rect 14829 9463 14887 9469
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9500 15623 9503
rect 15930 9500 15936 9512
rect 15611 9472 15936 9500
rect 15611 9469 15623 9472
rect 15565 9463 15623 9469
rect 15930 9460 15936 9472
rect 15988 9460 15994 9512
rect 17770 9460 17776 9512
rect 17828 9460 17834 9512
rect 20438 9460 20444 9512
rect 20496 9500 20502 9512
rect 20533 9503 20591 9509
rect 20533 9500 20545 9503
rect 20496 9472 20545 9500
rect 20496 9460 20502 9472
rect 20533 9469 20545 9472
rect 20579 9469 20591 9503
rect 21910 9500 21916 9512
rect 21823 9472 21916 9500
rect 20533 9463 20591 9469
rect 21910 9460 21916 9472
rect 21968 9500 21974 9512
rect 22373 9503 22431 9509
rect 22373 9500 22385 9503
rect 21968 9472 22385 9500
rect 21968 9460 21974 9472
rect 22373 9469 22385 9472
rect 22419 9469 22431 9503
rect 22373 9463 22431 9469
rect 23658 9460 23664 9512
rect 23716 9500 23722 9512
rect 24029 9503 24087 9509
rect 24029 9500 24041 9503
rect 23716 9472 24041 9500
rect 23716 9460 23722 9472
rect 24029 9469 24041 9472
rect 24075 9469 24087 9503
rect 24320 9500 24348 9531
rect 24762 9500 24768 9512
rect 24320 9472 24768 9500
rect 24029 9463 24087 9469
rect 24762 9460 24768 9472
rect 24820 9460 24826 9512
rect 25222 9500 25228 9512
rect 25183 9472 25228 9500
rect 25222 9460 25228 9472
rect 25280 9500 25286 9512
rect 25777 9503 25835 9509
rect 25777 9500 25789 9503
rect 25280 9472 25789 9500
rect 25280 9460 25286 9472
rect 25777 9469 25789 9472
rect 25823 9469 25835 9503
rect 25777 9463 25835 9469
rect 8570 9432 8576 9444
rect 7944 9404 8576 9432
rect 6825 9395 6883 9401
rect 8570 9392 8576 9404
rect 8628 9392 8634 9444
rect 10965 9435 11023 9441
rect 10965 9432 10977 9435
rect 9968 9404 10977 9432
rect 3237 9367 3295 9373
rect 3237 9364 3249 9367
rect 2884 9336 3249 9364
rect 2593 9327 2651 9333
rect 3237 9333 3249 9336
rect 3283 9364 3295 9367
rect 3418 9364 3424 9376
rect 3283 9336 3424 9364
rect 3283 9333 3295 9336
rect 3237 9327 3295 9333
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 5350 9364 5356 9376
rect 5311 9336 5356 9364
rect 5350 9324 5356 9336
rect 5408 9324 5414 9376
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 5721 9367 5779 9373
rect 5721 9364 5733 9367
rect 5500 9336 5733 9364
rect 5500 9324 5506 9336
rect 5721 9333 5733 9336
rect 5767 9364 5779 9367
rect 5994 9364 6000 9376
rect 5767 9336 6000 9364
rect 5767 9333 5779 9336
rect 5721 9327 5779 9333
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 6181 9367 6239 9373
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 6270 9364 6276 9376
rect 6227 9336 6276 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 7558 9364 7564 9376
rect 7519 9336 7564 9364
rect 7558 9324 7564 9336
rect 7616 9324 7622 9376
rect 9214 9324 9220 9376
rect 9272 9364 9278 9376
rect 9968 9373 9996 9404
rect 10965 9401 10977 9404
rect 11011 9401 11023 9435
rect 10965 9395 11023 9401
rect 13262 9392 13268 9444
rect 13320 9392 13326 9444
rect 14274 9392 14280 9444
rect 14332 9432 14338 9444
rect 14921 9435 14979 9441
rect 14921 9432 14933 9435
rect 14332 9404 14933 9432
rect 14332 9392 14338 9404
rect 14921 9401 14933 9404
rect 14967 9401 14979 9435
rect 16114 9432 16120 9444
rect 14921 9395 14979 9401
rect 15856 9404 16120 9432
rect 15856 9376 15884 9404
rect 16114 9392 16120 9404
rect 16172 9432 16178 9444
rect 16485 9435 16543 9441
rect 16485 9432 16497 9435
rect 16172 9404 16497 9432
rect 16172 9392 16178 9404
rect 16485 9401 16497 9404
rect 16531 9401 16543 9435
rect 16485 9395 16543 9401
rect 17954 9392 17960 9444
rect 18012 9432 18018 9444
rect 18294 9435 18352 9441
rect 18294 9432 18306 9435
rect 18012 9404 18306 9432
rect 18012 9392 18018 9404
rect 18294 9401 18306 9404
rect 18340 9401 18352 9435
rect 24121 9435 24179 9441
rect 24121 9432 24133 9435
rect 18294 9395 18352 9401
rect 22020 9404 24133 9432
rect 9953 9367 10011 9373
rect 9953 9364 9965 9367
rect 9272 9336 9965 9364
rect 9272 9324 9278 9336
rect 9953 9333 9965 9336
rect 9999 9333 10011 9367
rect 9953 9327 10011 9333
rect 10134 9324 10140 9376
rect 10192 9364 10198 9376
rect 10321 9367 10379 9373
rect 10321 9364 10333 9367
rect 10192 9336 10333 9364
rect 10192 9324 10198 9336
rect 10321 9333 10333 9336
rect 10367 9364 10379 9367
rect 10873 9367 10931 9373
rect 10873 9364 10885 9367
rect 10367 9336 10885 9364
rect 10367 9333 10379 9336
rect 10321 9327 10379 9333
rect 10873 9333 10885 9336
rect 10919 9333 10931 9367
rect 11606 9364 11612 9376
rect 11567 9336 11612 9364
rect 10873 9327 10931 9333
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 14458 9364 14464 9376
rect 14419 9336 14464 9364
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 15838 9364 15844 9376
rect 15799 9336 15844 9364
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 16022 9364 16028 9376
rect 15983 9336 16028 9364
rect 16022 9324 16028 9336
rect 16080 9324 16086 9376
rect 16390 9364 16396 9376
rect 16351 9336 16396 9364
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 22020 9373 22048 9404
rect 24121 9401 24133 9404
rect 24167 9432 24179 9435
rect 25041 9435 25099 9441
rect 25041 9432 25053 9435
rect 24167 9404 25053 9432
rect 24167 9401 24179 9404
rect 24121 9395 24179 9401
rect 25041 9401 25053 9404
rect 25087 9401 25099 9435
rect 25041 9395 25099 9401
rect 22005 9367 22063 9373
rect 22005 9333 22017 9367
rect 22051 9333 22063 9367
rect 22005 9327 22063 9333
rect 24765 9367 24823 9373
rect 24765 9333 24777 9367
rect 24811 9364 24823 9367
rect 24854 9364 24860 9376
rect 24811 9336 24860 9364
rect 24811 9333 24823 9336
rect 24765 9327 24823 9333
rect 24854 9324 24860 9336
rect 24912 9324 24918 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1578 9160 1584 9172
rect 1539 9132 1584 9160
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 2222 9120 2228 9172
rect 2280 9160 2286 9172
rect 2317 9163 2375 9169
rect 2317 9160 2329 9163
rect 2280 9132 2329 9160
rect 2280 9120 2286 9132
rect 2317 9129 2329 9132
rect 2363 9160 2375 9163
rect 4062 9160 4068 9172
rect 2363 9132 4068 9160
rect 2363 9129 2375 9132
rect 2317 9123 2375 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 7190 9160 7196 9172
rect 7151 9132 7196 9160
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 8662 9120 8668 9172
rect 8720 9160 8726 9172
rect 8941 9163 8999 9169
rect 8941 9160 8953 9163
rect 8720 9132 8953 9160
rect 8720 9120 8726 9132
rect 8941 9129 8953 9132
rect 8987 9129 8999 9163
rect 8941 9123 8999 9129
rect 11054 9120 11060 9172
rect 11112 9160 11118 9172
rect 11609 9163 11667 9169
rect 11609 9160 11621 9163
rect 11112 9132 11621 9160
rect 11112 9120 11118 9132
rect 11609 9129 11621 9132
rect 11655 9129 11667 9163
rect 11609 9123 11667 9129
rect 12434 9120 12440 9172
rect 12492 9160 12498 9172
rect 15010 9160 15016 9172
rect 12492 9132 12537 9160
rect 14971 9132 15016 9160
rect 12492 9120 12498 9132
rect 15010 9120 15016 9132
rect 15068 9160 15074 9172
rect 15378 9160 15384 9172
rect 15068 9132 15384 9160
rect 15068 9120 15074 9132
rect 15378 9120 15384 9132
rect 15436 9160 15442 9172
rect 16669 9163 16727 9169
rect 16669 9160 16681 9163
rect 15436 9132 16681 9160
rect 15436 9120 15442 9132
rect 16669 9129 16681 9132
rect 16715 9129 16727 9163
rect 17586 9160 17592 9172
rect 17547 9132 17592 9160
rect 16669 9123 16727 9129
rect 17586 9120 17592 9132
rect 17644 9120 17650 9172
rect 18049 9163 18107 9169
rect 18049 9129 18061 9163
rect 18095 9160 18107 9163
rect 18690 9160 18696 9172
rect 18095 9132 18696 9160
rect 18095 9129 18107 9132
rect 18049 9123 18107 9129
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 20254 9160 20260 9172
rect 20215 9132 20260 9160
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 20346 9120 20352 9172
rect 20404 9160 20410 9172
rect 21174 9160 21180 9172
rect 20404 9132 21180 9160
rect 20404 9120 20410 9132
rect 21174 9120 21180 9132
rect 21232 9160 21238 9172
rect 21269 9163 21327 9169
rect 21269 9160 21281 9163
rect 21232 9132 21281 9160
rect 21232 9120 21238 9132
rect 21269 9129 21281 9132
rect 21315 9129 21327 9163
rect 21269 9123 21327 9129
rect 21358 9120 21364 9172
rect 21416 9160 21422 9172
rect 22097 9163 22155 9169
rect 21416 9132 21461 9160
rect 21416 9120 21422 9132
rect 22097 9129 22109 9163
rect 22143 9160 22155 9163
rect 23106 9160 23112 9172
rect 22143 9132 23112 9160
rect 22143 9129 22155 9132
rect 22097 9123 22155 9129
rect 23106 9120 23112 9132
rect 23164 9160 23170 9172
rect 23293 9163 23351 9169
rect 23293 9160 23305 9163
rect 23164 9132 23305 9160
rect 23164 9120 23170 9132
rect 23293 9129 23305 9132
rect 23339 9129 23351 9163
rect 23293 9123 23351 9129
rect 2777 9095 2835 9101
rect 2777 9061 2789 9095
rect 2823 9092 2835 9095
rect 2866 9092 2872 9104
rect 2823 9064 2872 9092
rect 2823 9061 2835 9064
rect 2777 9055 2835 9061
rect 2866 9052 2872 9064
rect 2924 9052 2930 9104
rect 6178 9052 6184 9104
rect 6236 9092 6242 9104
rect 7653 9095 7711 9101
rect 7653 9092 7665 9095
rect 6236 9064 7665 9092
rect 6236 9052 6242 9064
rect 7653 9061 7665 9064
rect 7699 9061 7711 9095
rect 7653 9055 7711 9061
rect 15556 9095 15614 9101
rect 15556 9061 15568 9095
rect 15602 9092 15614 9095
rect 15654 9092 15660 9104
rect 15602 9064 15660 9092
rect 15602 9061 15614 9064
rect 15556 9055 15614 9061
rect 15654 9052 15660 9064
rect 15712 9052 15718 9104
rect 17604 9092 17632 9120
rect 17604 9064 18635 9092
rect 1394 9024 1400 9036
rect 1307 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 9024 1458 9036
rect 1854 9024 1860 9036
rect 1452 8996 1860 9024
rect 1452 8984 1458 8996
rect 1854 8984 1860 8996
rect 1912 8984 1918 9036
rect 4338 9033 4344 9036
rect 4332 9024 4344 9033
rect 4299 8996 4344 9024
rect 4332 8987 4344 8996
rect 4338 8984 4344 8987
rect 4396 8984 4402 9036
rect 7561 9027 7619 9033
rect 7561 8993 7573 9027
rect 7607 9024 7619 9027
rect 8018 9024 8024 9036
rect 7607 8996 8024 9024
rect 7607 8993 7619 8996
rect 7561 8987 7619 8993
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 8297 9027 8355 9033
rect 8297 8993 8309 9027
rect 8343 9024 8355 9027
rect 8386 9024 8392 9036
rect 8343 8996 8392 9024
rect 8343 8993 8355 8996
rect 8297 8987 8355 8993
rect 8386 8984 8392 8996
rect 8444 8984 8450 9036
rect 9582 9024 9588 9036
rect 8496 8996 9588 9024
rect 2590 8916 2596 8968
rect 2648 8956 2654 8968
rect 2869 8959 2927 8965
rect 2869 8956 2881 8959
rect 2648 8928 2881 8956
rect 2648 8916 2654 8928
rect 2869 8925 2881 8928
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 2958 8916 2964 8968
rect 3016 8956 3022 8968
rect 4062 8956 4068 8968
rect 3016 8928 3061 8956
rect 4023 8928 4068 8956
rect 3016 8916 3022 8928
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 7742 8956 7748 8968
rect 7703 8928 7748 8956
rect 7742 8916 7748 8928
rect 7800 8916 7806 8968
rect 8496 8956 8524 8996
rect 9582 8984 9588 8996
rect 9640 8984 9646 9036
rect 10502 9033 10508 9036
rect 10496 9024 10508 9033
rect 10463 8996 10508 9024
rect 10496 8987 10508 8996
rect 10502 8984 10508 8987
rect 10560 8984 10566 9036
rect 12986 9033 12992 9036
rect 12980 9024 12992 9033
rect 12947 8996 12992 9024
rect 12980 8987 12992 8996
rect 12986 8984 12992 8987
rect 13044 8984 13050 9036
rect 14734 8984 14740 9036
rect 14792 9024 14798 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 14792 8996 15301 9024
rect 14792 8984 14798 8996
rect 15289 8993 15301 8996
rect 15335 8993 15347 9027
rect 15289 8987 15347 8993
rect 18046 8984 18052 9036
rect 18104 9024 18110 9036
rect 18230 9024 18236 9036
rect 18104 8996 18236 9024
rect 18104 8984 18110 8996
rect 18230 8984 18236 8996
rect 18288 9024 18294 9036
rect 18417 9027 18475 9033
rect 18417 9024 18429 9027
rect 18288 8996 18429 9024
rect 18288 8984 18294 8996
rect 18417 8993 18429 8996
rect 18463 8993 18475 9027
rect 18417 8987 18475 8993
rect 8220 8928 8524 8956
rect 2409 8891 2467 8897
rect 2409 8857 2421 8891
rect 2455 8888 2467 8891
rect 8220 8888 8248 8928
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 8665 8959 8723 8965
rect 8665 8956 8677 8959
rect 8628 8928 8677 8956
rect 8628 8916 8634 8928
rect 8665 8925 8677 8928
rect 8711 8956 8723 8959
rect 10226 8956 10232 8968
rect 8711 8928 10232 8956
rect 8711 8925 8723 8928
rect 8665 8919 8723 8925
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 12434 8916 12440 8968
rect 12492 8956 12498 8968
rect 18607 8965 18635 9064
rect 20622 9052 20628 9104
rect 20680 9092 20686 9104
rect 21376 9092 21404 9120
rect 20680 9064 21404 9092
rect 24020 9095 24078 9101
rect 20680 9052 20686 9064
rect 24020 9061 24032 9095
rect 24066 9092 24078 9095
rect 24762 9092 24768 9104
rect 24066 9064 24768 9092
rect 24066 9061 24078 9064
rect 24020 9055 24078 9061
rect 24762 9052 24768 9064
rect 24820 9052 24826 9104
rect 19705 9027 19763 9033
rect 19705 8993 19717 9027
rect 19751 9024 19763 9027
rect 20530 9024 20536 9036
rect 19751 8996 20536 9024
rect 19751 8993 19763 8996
rect 19705 8987 19763 8993
rect 20530 8984 20536 8996
rect 20588 8984 20594 9036
rect 22830 8984 22836 9036
rect 22888 9024 22894 9036
rect 23750 9024 23756 9036
rect 22888 8996 23756 9024
rect 22888 8984 22894 8996
rect 23750 8984 23756 8996
rect 23808 8984 23814 9036
rect 12713 8959 12771 8965
rect 12713 8956 12725 8959
rect 12492 8928 12725 8956
rect 12492 8916 12498 8928
rect 12713 8925 12725 8928
rect 12759 8925 12771 8959
rect 12713 8919 12771 8925
rect 18509 8959 18567 8965
rect 18509 8925 18521 8959
rect 18555 8925 18567 8959
rect 18509 8919 18567 8925
rect 18601 8959 18659 8965
rect 18601 8925 18613 8959
rect 18647 8925 18659 8959
rect 18601 8919 18659 8925
rect 20717 8959 20775 8965
rect 20717 8925 20729 8959
rect 20763 8956 20775 8959
rect 20898 8956 20904 8968
rect 20763 8928 20904 8956
rect 20763 8925 20775 8928
rect 20717 8919 20775 8925
rect 2455 8860 4108 8888
rect 2455 8857 2467 8860
rect 2409 8851 2467 8857
rect 1946 8820 1952 8832
rect 1907 8792 1952 8820
rect 1946 8780 1952 8792
rect 2004 8780 2010 8832
rect 3326 8780 3332 8832
rect 3384 8820 3390 8832
rect 3421 8823 3479 8829
rect 3421 8820 3433 8823
rect 3384 8792 3433 8820
rect 3384 8780 3390 8792
rect 3421 8789 3433 8792
rect 3467 8789 3479 8823
rect 3878 8820 3884 8832
rect 3839 8792 3884 8820
rect 3421 8783 3479 8789
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 4080 8820 4108 8860
rect 5276 8860 8248 8888
rect 5276 8820 5304 8860
rect 8294 8848 8300 8900
rect 8352 8888 8358 8900
rect 9309 8891 9367 8897
rect 9309 8888 9321 8891
rect 8352 8860 9321 8888
rect 8352 8848 8358 8860
rect 9309 8857 9321 8860
rect 9355 8857 9367 8891
rect 9309 8851 9367 8857
rect 14737 8891 14795 8897
rect 14737 8857 14749 8891
rect 14783 8888 14795 8891
rect 15102 8888 15108 8900
rect 14783 8860 15108 8888
rect 14783 8857 14795 8860
rect 14737 8851 14795 8857
rect 15102 8848 15108 8860
rect 15160 8848 15166 8900
rect 17494 8848 17500 8900
rect 17552 8888 17558 8900
rect 18524 8888 18552 8919
rect 20898 8916 20904 8928
rect 20956 8916 20962 8968
rect 21453 8959 21511 8965
rect 21453 8925 21465 8959
rect 21499 8925 21511 8959
rect 21453 8919 21511 8925
rect 22741 8959 22799 8965
rect 22741 8925 22753 8959
rect 22787 8956 22799 8959
rect 23198 8956 23204 8968
rect 22787 8928 23204 8956
rect 22787 8925 22799 8928
rect 22741 8919 22799 8925
rect 17552 8860 18552 8888
rect 17552 8848 17558 8860
rect 5442 8820 5448 8832
rect 4080 8792 5304 8820
rect 5403 8792 5448 8820
rect 5442 8780 5448 8792
rect 5500 8780 5506 8832
rect 5994 8820 6000 8832
rect 5955 8792 6000 8820
rect 5994 8780 6000 8792
rect 6052 8780 6058 8832
rect 6362 8820 6368 8832
rect 6323 8792 6368 8820
rect 6362 8780 6368 8792
rect 6420 8780 6426 8832
rect 7098 8820 7104 8832
rect 7059 8792 7104 8820
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 7190 8780 7196 8832
rect 7248 8820 7254 8832
rect 9398 8820 9404 8832
rect 7248 8792 9404 8820
rect 7248 8780 7254 8792
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 9858 8820 9864 8832
rect 9819 8792 9864 8820
rect 9858 8780 9864 8792
rect 9916 8780 9922 8832
rect 10410 8780 10416 8832
rect 10468 8820 10474 8832
rect 10962 8820 10968 8832
rect 10468 8792 10968 8820
rect 10468 8780 10474 8792
rect 10962 8780 10968 8792
rect 11020 8780 11026 8832
rect 14090 8820 14096 8832
rect 14051 8792 14096 8820
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 17954 8820 17960 8832
rect 17915 8792 17960 8820
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 18524 8820 18552 8860
rect 21266 8848 21272 8900
rect 21324 8888 21330 8900
rect 21468 8888 21496 8919
rect 23198 8916 23204 8928
rect 23256 8916 23262 8968
rect 21324 8860 21496 8888
rect 21324 8848 21330 8860
rect 18598 8820 18604 8832
rect 18524 8792 18604 8820
rect 18598 8780 18604 8792
rect 18656 8780 18662 8832
rect 19058 8820 19064 8832
rect 19019 8792 19064 8820
rect 19058 8780 19064 8792
rect 19116 8780 19122 8832
rect 19426 8820 19432 8832
rect 19387 8792 19432 8820
rect 19426 8780 19432 8792
rect 19484 8780 19490 8832
rect 19889 8823 19947 8829
rect 19889 8789 19901 8823
rect 19935 8820 19947 8823
rect 20438 8820 20444 8832
rect 19935 8792 20444 8820
rect 19935 8789 19947 8792
rect 19889 8783 19947 8789
rect 20438 8780 20444 8792
rect 20496 8780 20502 8832
rect 20714 8780 20720 8832
rect 20772 8820 20778 8832
rect 20901 8823 20959 8829
rect 20901 8820 20913 8823
rect 20772 8792 20913 8820
rect 20772 8780 20778 8792
rect 20901 8789 20913 8792
rect 20947 8789 20959 8823
rect 20901 8783 20959 8789
rect 21358 8780 21364 8832
rect 21416 8820 21422 8832
rect 21726 8820 21732 8832
rect 21416 8792 21732 8820
rect 21416 8780 21422 8792
rect 21726 8780 21732 8792
rect 21784 8780 21790 8832
rect 25130 8820 25136 8832
rect 25091 8792 25136 8820
rect 25130 8780 25136 8792
rect 25188 8780 25194 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2133 8619 2191 8625
rect 2133 8585 2145 8619
rect 2179 8616 2191 8619
rect 2590 8616 2596 8628
rect 2179 8588 2596 8616
rect 2179 8585 2191 8588
rect 2133 8579 2191 8585
rect 2590 8576 2596 8588
rect 2648 8616 2654 8628
rect 4614 8616 4620 8628
rect 2648 8588 4620 8616
rect 2648 8576 2654 8588
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 5169 8619 5227 8625
rect 5169 8585 5181 8619
rect 5215 8616 5227 8619
rect 5258 8616 5264 8628
rect 5215 8588 5264 8616
rect 5215 8585 5227 8588
rect 5169 8579 5227 8585
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 7190 8616 7196 8628
rect 7151 8588 7196 8616
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 10137 8619 10195 8625
rect 10137 8616 10149 8619
rect 7760 8588 10149 8616
rect 4062 8508 4068 8560
rect 4120 8548 4126 8560
rect 4249 8551 4307 8557
rect 4249 8548 4261 8551
rect 4120 8520 4261 8548
rect 4120 8508 4126 8520
rect 4249 8517 4261 8520
rect 4295 8548 4307 8551
rect 5350 8548 5356 8560
rect 4295 8520 5356 8548
rect 4295 8517 4307 8520
rect 4249 8511 4307 8517
rect 5350 8508 5356 8520
rect 5408 8548 5414 8560
rect 5534 8548 5540 8560
rect 5408 8520 5540 8548
rect 5408 8508 5414 8520
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 7282 8508 7288 8560
rect 7340 8548 7346 8560
rect 7466 8548 7472 8560
rect 7340 8520 7472 8548
rect 7340 8508 7346 8520
rect 7466 8508 7472 8520
rect 7524 8508 7530 8560
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8480 1823 8483
rect 1811 8452 2360 8480
rect 1811 8449 1823 8452
rect 1765 8443 1823 8449
rect 2222 8412 2228 8424
rect 2183 8384 2228 8412
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 2332 8412 2360 8452
rect 5442 8440 5448 8492
rect 5500 8480 5506 8492
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 5500 8452 5825 8480
rect 5500 8440 5506 8452
rect 5813 8449 5825 8452
rect 5859 8480 5871 8483
rect 6181 8483 6239 8489
rect 6181 8480 6193 8483
rect 5859 8452 6193 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6181 8449 6193 8452
rect 6227 8449 6239 8483
rect 6181 8443 6239 8449
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 7760 8489 7788 8588
rect 10137 8585 10149 8588
rect 10183 8616 10195 8619
rect 10502 8616 10508 8628
rect 10183 8588 10508 8616
rect 10183 8585 10195 8588
rect 10137 8579 10195 8585
rect 10502 8576 10508 8588
rect 10560 8616 10566 8628
rect 10686 8616 10692 8628
rect 10560 8588 10692 8616
rect 10560 8576 10566 8588
rect 10686 8576 10692 8588
rect 10744 8616 10750 8628
rect 11057 8619 11115 8625
rect 11057 8616 11069 8619
rect 10744 8588 11069 8616
rect 10744 8576 10750 8588
rect 11057 8585 11069 8588
rect 11103 8585 11115 8619
rect 11057 8579 11115 8585
rect 14182 8576 14188 8628
rect 14240 8616 14246 8628
rect 16666 8616 16672 8628
rect 14240 8588 16672 8616
rect 14240 8576 14246 8588
rect 16666 8576 16672 8588
rect 16724 8576 16730 8628
rect 17494 8616 17500 8628
rect 17455 8588 17500 8616
rect 17494 8576 17500 8588
rect 17552 8576 17558 8628
rect 17954 8576 17960 8628
rect 18012 8616 18018 8628
rect 19429 8619 19487 8625
rect 19429 8616 19441 8619
rect 18012 8588 19441 8616
rect 18012 8576 18018 8588
rect 19429 8585 19441 8588
rect 19475 8585 19487 8619
rect 19429 8579 19487 8585
rect 20165 8619 20223 8625
rect 20165 8585 20177 8619
rect 20211 8616 20223 8619
rect 20346 8616 20352 8628
rect 20211 8588 20352 8616
rect 20211 8585 20223 8588
rect 20165 8579 20223 8585
rect 20346 8576 20352 8588
rect 20404 8576 20410 8628
rect 20533 8619 20591 8625
rect 20533 8585 20545 8619
rect 20579 8616 20591 8619
rect 20622 8616 20628 8628
rect 20579 8588 20628 8616
rect 20579 8585 20591 8588
rect 20533 8579 20591 8585
rect 20622 8576 20628 8588
rect 20680 8576 20686 8628
rect 24854 8616 24860 8628
rect 24815 8588 24860 8616
rect 24854 8576 24860 8588
rect 24912 8576 24918 8628
rect 25130 8576 25136 8628
rect 25188 8616 25194 8628
rect 25225 8619 25283 8625
rect 25225 8616 25237 8619
rect 25188 8588 25237 8616
rect 25188 8576 25194 8588
rect 25225 8585 25237 8588
rect 25271 8585 25283 8619
rect 25590 8616 25596 8628
rect 25551 8588 25596 8616
rect 25225 8579 25283 8585
rect 25590 8576 25596 8588
rect 25648 8576 25654 8628
rect 8570 8548 8576 8560
rect 8531 8520 8576 8548
rect 8570 8508 8576 8520
rect 8628 8508 8634 8560
rect 16298 8548 16304 8560
rect 16040 8520 16304 8548
rect 7745 8483 7803 8489
rect 7745 8480 7757 8483
rect 7156 8452 7757 8480
rect 7156 8440 7162 8452
rect 7745 8449 7757 8452
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 8018 8440 8024 8492
rect 8076 8480 8082 8492
rect 8297 8483 8355 8489
rect 8297 8480 8309 8483
rect 8076 8452 8309 8480
rect 8076 8440 8082 8452
rect 8297 8449 8309 8452
rect 8343 8480 8355 8483
rect 8343 8452 8892 8480
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 2866 8412 2872 8424
rect 2332 8384 2872 8412
rect 2866 8372 2872 8384
rect 2924 8412 2930 8424
rect 3050 8412 3056 8424
rect 2924 8384 3056 8412
rect 2924 8372 2930 8384
rect 3050 8372 3056 8384
rect 3108 8372 3114 8424
rect 5350 8372 5356 8424
rect 5408 8412 5414 8424
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 5408 8384 5549 8412
rect 5408 8372 5414 8384
rect 5537 8381 5549 8384
rect 5583 8412 5595 8415
rect 8036 8412 8064 8440
rect 5583 8384 8064 8412
rect 5583 8381 5595 8384
rect 5537 8375 5595 8381
rect 8570 8372 8576 8424
rect 8628 8412 8634 8424
rect 8757 8415 8815 8421
rect 8757 8412 8769 8415
rect 8628 8384 8769 8412
rect 8628 8372 8634 8384
rect 8757 8381 8769 8384
rect 8803 8381 8815 8415
rect 8864 8412 8892 8452
rect 10226 8440 10232 8492
rect 10284 8480 10290 8492
rect 10689 8483 10747 8489
rect 10689 8480 10701 8483
rect 10284 8452 10701 8480
rect 10284 8440 10290 8452
rect 10689 8449 10701 8452
rect 10735 8480 10747 8483
rect 11054 8480 11060 8492
rect 10735 8452 11060 8480
rect 10735 8449 10747 8452
rect 10689 8443 10747 8449
rect 11054 8440 11060 8452
rect 11112 8480 11118 8492
rect 11238 8480 11244 8492
rect 11112 8452 11244 8480
rect 11112 8440 11118 8452
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11606 8440 11612 8492
rect 11664 8480 11670 8492
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 11664 8452 11897 8480
rect 11664 8440 11670 8452
rect 11885 8449 11897 8452
rect 11931 8480 11943 8483
rect 11931 8452 12572 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 9306 8412 9312 8424
rect 8864 8384 9312 8412
rect 8757 8375 8815 8381
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 11256 8412 11284 8440
rect 12161 8415 12219 8421
rect 12161 8412 12173 8415
rect 11256 8384 12173 8412
rect 12161 8381 12173 8384
rect 12207 8412 12219 8415
rect 12434 8412 12440 8424
rect 12207 8384 12440 8412
rect 12207 8381 12219 8384
rect 12161 8375 12219 8381
rect 12434 8372 12440 8384
rect 12492 8372 12498 8424
rect 12544 8412 12572 8452
rect 12704 8415 12762 8421
rect 12704 8412 12716 8415
rect 12544 8384 12716 8412
rect 12704 8381 12716 8384
rect 12750 8412 12762 8415
rect 14090 8412 14096 8424
rect 12750 8384 14096 8412
rect 12750 8381 12762 8384
rect 12704 8375 12762 8381
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 14734 8412 14740 8424
rect 14292 8384 14740 8412
rect 1946 8304 1952 8356
rect 2004 8344 2010 8356
rect 2498 8353 2504 8356
rect 2470 8347 2504 8353
rect 2470 8344 2482 8347
rect 2004 8316 2482 8344
rect 2004 8304 2010 8316
rect 2470 8313 2482 8316
rect 2556 8344 2562 8356
rect 4338 8344 4344 8356
rect 2556 8316 2618 8344
rect 2700 8316 4344 8344
rect 2470 8307 2504 8313
rect 2498 8304 2504 8307
rect 2556 8304 2562 8316
rect 2590 8236 2596 8288
rect 2648 8276 2654 8288
rect 2700 8276 2728 8316
rect 3620 8285 3648 8316
rect 4338 8304 4344 8316
rect 4396 8344 4402 8356
rect 4525 8347 4583 8353
rect 4525 8344 4537 8347
rect 4396 8316 4537 8344
rect 4396 8304 4402 8316
rect 4525 8313 4537 8316
rect 4571 8313 4583 8347
rect 4525 8307 4583 8313
rect 5077 8347 5135 8353
rect 5077 8313 5089 8347
rect 5123 8344 5135 8347
rect 5629 8347 5687 8353
rect 5629 8344 5641 8347
rect 5123 8316 5641 8344
rect 5123 8313 5135 8316
rect 5077 8307 5135 8313
rect 5629 8313 5641 8316
rect 5675 8344 5687 8347
rect 6178 8344 6184 8356
rect 5675 8316 6184 8344
rect 5675 8313 5687 8316
rect 5629 8307 5687 8313
rect 6178 8304 6184 8316
rect 6236 8344 6242 8356
rect 6549 8347 6607 8353
rect 6549 8344 6561 8347
rect 6236 8316 6561 8344
rect 6236 8304 6242 8316
rect 6549 8313 6561 8316
rect 6595 8313 6607 8347
rect 7653 8347 7711 8353
rect 7653 8344 7665 8347
rect 6549 8307 6607 8313
rect 7024 8316 7665 8344
rect 2648 8248 2728 8276
rect 3605 8279 3663 8285
rect 2648 8236 2654 8248
rect 3605 8245 3617 8279
rect 3651 8245 3663 8279
rect 3605 8239 3663 8245
rect 5442 8236 5448 8288
rect 5500 8276 5506 8288
rect 7024 8285 7052 8316
rect 7653 8313 7665 8316
rect 7699 8313 7711 8347
rect 7653 8307 7711 8313
rect 8662 8304 8668 8356
rect 8720 8344 8726 8356
rect 9002 8347 9060 8353
rect 9002 8344 9014 8347
rect 8720 8316 9014 8344
rect 8720 8304 8726 8316
rect 9002 8313 9014 8316
rect 9048 8313 9060 8347
rect 12452 8344 12480 8372
rect 12894 8344 12900 8356
rect 12452 8316 12900 8344
rect 9002 8307 9060 8313
rect 12894 8304 12900 8316
rect 12952 8344 12958 8356
rect 14292 8344 14320 8384
rect 14734 8372 14740 8384
rect 14792 8412 14798 8424
rect 15010 8412 15016 8424
rect 14792 8384 15016 8412
rect 14792 8372 14798 8384
rect 15010 8372 15016 8384
rect 15068 8372 15074 8424
rect 15102 8372 15108 8424
rect 15160 8412 15166 8424
rect 15160 8384 15332 8412
rect 15160 8372 15166 8384
rect 15304 8353 15332 8384
rect 15562 8372 15568 8424
rect 15620 8412 15626 8424
rect 16040 8412 16068 8520
rect 16298 8508 16304 8520
rect 16356 8548 16362 8560
rect 16393 8551 16451 8557
rect 16393 8548 16405 8551
rect 16356 8520 16405 8548
rect 16356 8508 16362 8520
rect 16393 8517 16405 8520
rect 16439 8517 16451 8551
rect 16393 8511 16451 8517
rect 17865 8551 17923 8557
rect 17865 8517 17877 8551
rect 17911 8548 17923 8551
rect 18046 8548 18052 8560
rect 17911 8520 18052 8548
rect 17911 8517 17923 8520
rect 17865 8511 17923 8517
rect 18046 8508 18052 8520
rect 18104 8508 18110 8560
rect 21726 8508 21732 8560
rect 21784 8548 21790 8560
rect 22005 8551 22063 8557
rect 22005 8548 22017 8551
rect 21784 8520 22017 8548
rect 21784 8508 21790 8520
rect 22005 8517 22017 8520
rect 22051 8517 22063 8551
rect 22005 8511 22063 8517
rect 24486 8480 24492 8492
rect 24399 8452 24492 8480
rect 24486 8440 24492 8452
rect 24544 8480 24550 8492
rect 25148 8480 25176 8576
rect 24544 8452 25176 8480
rect 24544 8440 24550 8452
rect 15620 8384 16068 8412
rect 15620 8372 15626 8384
rect 17770 8372 17776 8424
rect 17828 8412 17834 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 17828 8384 18061 8412
rect 17828 8372 17834 8384
rect 18049 8381 18061 8384
rect 18095 8412 18107 8415
rect 20622 8412 20628 8424
rect 18095 8384 20628 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 20622 8372 20628 8384
rect 20680 8372 20686 8424
rect 23109 8415 23167 8421
rect 23109 8381 23121 8415
rect 23155 8412 23167 8415
rect 24305 8415 24363 8421
rect 24305 8412 24317 8415
rect 23155 8384 24317 8412
rect 23155 8381 23167 8384
rect 23109 8375 23167 8381
rect 24305 8381 24317 8384
rect 24351 8412 24363 8415
rect 24670 8412 24676 8424
rect 24351 8384 24676 8412
rect 24351 8381 24363 8384
rect 24305 8375 24363 8381
rect 24670 8372 24676 8384
rect 24728 8372 24734 8424
rect 25406 8412 25412 8424
rect 25367 8384 25412 8412
rect 25406 8372 25412 8384
rect 25464 8412 25470 8424
rect 25961 8415 26019 8421
rect 25961 8412 25973 8415
rect 25464 8384 25973 8412
rect 25464 8372 25470 8384
rect 25961 8381 25973 8384
rect 26007 8381 26019 8415
rect 25961 8375 26019 8381
rect 12952 8316 14320 8344
rect 12952 8304 12958 8316
rect 7009 8279 7067 8285
rect 7009 8276 7021 8279
rect 5500 8248 7021 8276
rect 5500 8236 5506 8248
rect 7009 8245 7021 8248
rect 7055 8245 7067 8279
rect 7558 8276 7564 8288
rect 7519 8248 7564 8276
rect 7009 8239 7067 8245
rect 7558 8236 7564 8248
rect 7616 8236 7622 8288
rect 11238 8276 11244 8288
rect 11199 8248 11244 8276
rect 11238 8236 11244 8248
rect 11296 8236 11302 8288
rect 12710 8236 12716 8288
rect 12768 8276 12774 8288
rect 13817 8279 13875 8285
rect 13817 8276 13829 8279
rect 12768 8248 13829 8276
rect 12768 8236 12774 8248
rect 13817 8245 13829 8248
rect 13863 8245 13875 8279
rect 14292 8276 14320 8316
rect 14553 8347 14611 8353
rect 14553 8313 14565 8347
rect 14599 8344 14611 8347
rect 15280 8347 15338 8353
rect 14599 8316 15240 8344
rect 14599 8313 14611 8316
rect 14553 8307 14611 8313
rect 14829 8279 14887 8285
rect 14829 8276 14841 8279
rect 14292 8248 14841 8276
rect 13817 8239 13875 8245
rect 14829 8245 14841 8248
rect 14875 8245 14887 8279
rect 15212 8276 15240 8316
rect 15280 8313 15292 8347
rect 15326 8344 15338 8347
rect 15378 8344 15384 8356
rect 15326 8316 15384 8344
rect 15326 8313 15338 8316
rect 15280 8307 15338 8313
rect 15378 8304 15384 8316
rect 15436 8304 15442 8356
rect 16758 8304 16764 8356
rect 16816 8344 16822 8356
rect 17129 8347 17187 8353
rect 17129 8344 17141 8347
rect 16816 8316 17141 8344
rect 16816 8304 16822 8316
rect 17129 8313 17141 8316
rect 17175 8344 17187 8347
rect 18316 8347 18374 8353
rect 18316 8344 18328 8347
rect 17175 8316 18328 8344
rect 17175 8313 17187 8316
rect 17129 8307 17187 8313
rect 18316 8313 18328 8316
rect 18362 8344 18374 8347
rect 19242 8344 19248 8356
rect 18362 8316 19248 8344
rect 18362 8313 18374 8316
rect 18316 8307 18374 8313
rect 19242 8304 19248 8316
rect 19300 8304 19306 8356
rect 20898 8353 20904 8356
rect 20870 8347 20904 8353
rect 20870 8344 20882 8347
rect 20364 8316 20882 8344
rect 20364 8288 20392 8316
rect 20870 8313 20882 8316
rect 20956 8344 20962 8356
rect 23474 8344 23480 8356
rect 20956 8316 22140 8344
rect 23435 8316 23480 8344
rect 20870 8307 20904 8313
rect 20898 8304 20904 8307
rect 20956 8304 20962 8316
rect 15654 8276 15660 8288
rect 15212 8248 15660 8276
rect 14829 8239 14887 8245
rect 15654 8236 15660 8248
rect 15712 8236 15718 8288
rect 20346 8236 20352 8288
rect 20404 8236 20410 8288
rect 22112 8276 22140 8316
rect 23474 8304 23480 8316
rect 23532 8344 23538 8356
rect 24213 8347 24271 8353
rect 24213 8344 24225 8347
rect 23532 8316 24225 8344
rect 23532 8304 23538 8316
rect 24213 8313 24225 8316
rect 24259 8313 24271 8347
rect 24213 8307 24271 8313
rect 22278 8276 22284 8288
rect 22112 8248 22284 8276
rect 22278 8236 22284 8248
rect 22336 8236 22342 8288
rect 22554 8276 22560 8288
rect 22515 8248 22560 8276
rect 22554 8236 22560 8248
rect 22612 8236 22618 8288
rect 23842 8276 23848 8288
rect 23803 8248 23848 8276
rect 23842 8236 23848 8248
rect 23900 8236 23906 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 2130 8032 2136 8084
rect 2188 8072 2194 8084
rect 2317 8075 2375 8081
rect 2317 8072 2329 8075
rect 2188 8044 2329 8072
rect 2188 8032 2194 8044
rect 2317 8041 2329 8044
rect 2363 8041 2375 8075
rect 2317 8035 2375 8041
rect 2498 8032 2504 8084
rect 2556 8072 2562 8084
rect 2777 8075 2835 8081
rect 2777 8072 2789 8075
rect 2556 8044 2789 8072
rect 2556 8032 2562 8044
rect 2777 8041 2789 8044
rect 2823 8041 2835 8075
rect 2777 8035 2835 8041
rect 5261 8075 5319 8081
rect 5261 8041 5273 8075
rect 5307 8072 5319 8075
rect 5350 8072 5356 8084
rect 5307 8044 5356 8072
rect 5307 8041 5319 8044
rect 5261 8035 5319 8041
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 7837 8075 7895 8081
rect 7837 8072 7849 8075
rect 7800 8044 7849 8072
rect 7800 8032 7806 8044
rect 7837 8041 7849 8044
rect 7883 8041 7895 8075
rect 7837 8035 7895 8041
rect 9214 8032 9220 8084
rect 9272 8072 9278 8084
rect 9582 8072 9588 8084
rect 9272 8044 9588 8072
rect 9272 8032 9278 8044
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 9732 8044 10149 8072
rect 9732 8032 9738 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 11238 8032 11244 8084
rect 11296 8072 11302 8084
rect 12069 8075 12127 8081
rect 12069 8072 12081 8075
rect 11296 8044 12081 8072
rect 11296 8032 11302 8044
rect 12069 8041 12081 8044
rect 12115 8072 12127 8075
rect 12158 8072 12164 8084
rect 12115 8044 12164 8072
rect 12115 8041 12127 8044
rect 12069 8035 12127 8041
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 12805 8075 12863 8081
rect 12805 8041 12817 8075
rect 12851 8072 12863 8075
rect 12894 8072 12900 8084
rect 12851 8044 12900 8072
rect 12851 8041 12863 8044
rect 12805 8035 12863 8041
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 12986 8032 12992 8084
rect 13044 8072 13050 8084
rect 13081 8075 13139 8081
rect 13081 8072 13093 8075
rect 13044 8044 13093 8072
rect 13044 8032 13050 8044
rect 13081 8041 13093 8044
rect 13127 8041 13139 8075
rect 13081 8035 13139 8041
rect 13538 8032 13544 8084
rect 13596 8072 13602 8084
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 13596 8044 13645 8072
rect 13596 8032 13602 8044
rect 13633 8041 13645 8044
rect 13679 8041 13691 8075
rect 13633 8035 13691 8041
rect 14001 8075 14059 8081
rect 14001 8041 14013 8075
rect 14047 8072 14059 8075
rect 14458 8072 14464 8084
rect 14047 8044 14464 8072
rect 14047 8041 14059 8044
rect 14001 8035 14059 8041
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 14737 8075 14795 8081
rect 14737 8041 14749 8075
rect 14783 8072 14795 8075
rect 14826 8072 14832 8084
rect 14783 8044 14832 8072
rect 14783 8041 14795 8044
rect 14737 8035 14795 8041
rect 1670 7964 1676 8016
rect 1728 7964 1734 8016
rect 2222 8004 2228 8016
rect 2183 7976 2228 8004
rect 2222 7964 2228 7976
rect 2280 7964 2286 8016
rect 2406 7964 2412 8016
rect 2464 8004 2470 8016
rect 2682 8004 2688 8016
rect 2464 7976 2688 8004
rect 2464 7964 2470 7976
rect 2682 7964 2688 7976
rect 2740 7964 2746 8016
rect 8389 8007 8447 8013
rect 8389 7973 8401 8007
rect 8435 8004 8447 8007
rect 8662 8004 8668 8016
rect 8435 7976 8668 8004
rect 8435 7973 8447 7976
rect 8389 7967 8447 7973
rect 8662 7964 8668 7976
rect 8720 7964 8726 8016
rect 11606 8004 11612 8016
rect 11519 7976 11612 8004
rect 11606 7964 11612 7976
rect 11664 8004 11670 8016
rect 12342 8004 12348 8016
rect 11664 7976 12348 8004
rect 11664 7964 11670 7976
rect 12342 7964 12348 7976
rect 12400 7964 12406 8016
rect 14093 8007 14151 8013
rect 14093 7973 14105 8007
rect 14139 8004 14151 8007
rect 14752 8004 14780 8035
rect 14826 8032 14832 8044
rect 14884 8032 14890 8084
rect 15102 8072 15108 8084
rect 15063 8044 15108 8072
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 16577 8075 16635 8081
rect 16577 8041 16589 8075
rect 16623 8072 16635 8075
rect 17402 8072 17408 8084
rect 16623 8044 17408 8072
rect 16623 8041 16635 8044
rect 16577 8035 16635 8041
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 17681 8075 17739 8081
rect 17681 8041 17693 8075
rect 17727 8072 17739 8075
rect 17862 8072 17868 8084
rect 17727 8044 17868 8072
rect 17727 8041 17739 8044
rect 17681 8035 17739 8041
rect 17862 8032 17868 8044
rect 17920 8032 17926 8084
rect 18046 8072 18052 8084
rect 17959 8044 18052 8072
rect 18046 8032 18052 8044
rect 18104 8072 18110 8084
rect 19058 8072 19064 8084
rect 18104 8044 19064 8072
rect 18104 8032 18110 8044
rect 19058 8032 19064 8044
rect 19116 8032 19122 8084
rect 19153 8075 19211 8081
rect 19153 8041 19165 8075
rect 19199 8072 19211 8075
rect 19242 8072 19248 8084
rect 19199 8044 19248 8072
rect 19199 8041 19211 8044
rect 19153 8035 19211 8041
rect 19242 8032 19248 8044
rect 19300 8032 19306 8084
rect 19613 8075 19671 8081
rect 19613 8041 19625 8075
rect 19659 8072 19671 8075
rect 20622 8072 20628 8084
rect 19659 8044 20628 8072
rect 19659 8041 19671 8044
rect 19613 8035 19671 8041
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 22278 8072 22284 8084
rect 22239 8044 22284 8072
rect 22278 8032 22284 8044
rect 22336 8032 22342 8084
rect 22738 8032 22744 8084
rect 22796 8072 22802 8084
rect 22833 8075 22891 8081
rect 22833 8072 22845 8075
rect 22796 8044 22845 8072
rect 22796 8032 22802 8044
rect 22833 8041 22845 8044
rect 22879 8041 22891 8075
rect 23750 8072 23756 8084
rect 23711 8044 23756 8072
rect 22833 8035 22891 8041
rect 23750 8032 23756 8044
rect 23808 8032 23814 8084
rect 14139 7976 14780 8004
rect 14139 7973 14151 7976
rect 14093 7967 14151 7973
rect 15010 7964 15016 8016
rect 15068 8004 15074 8016
rect 15473 8007 15531 8013
rect 15473 8004 15485 8007
rect 15068 7976 15485 8004
rect 15068 7964 15074 7976
rect 15473 7973 15485 7976
rect 15519 7973 15531 8007
rect 15473 7967 15531 7973
rect 17770 7964 17776 8016
rect 17828 8004 17834 8016
rect 18693 8007 18751 8013
rect 18693 8004 18705 8007
rect 17828 7976 18705 8004
rect 17828 7964 17834 7976
rect 18693 7973 18705 7976
rect 18739 7973 18751 8007
rect 18693 7967 18751 7973
rect 20349 8007 20407 8013
rect 20349 7973 20361 8007
rect 20395 8004 20407 8007
rect 20530 8004 20536 8016
rect 20395 7976 20536 8004
rect 20395 7973 20407 7976
rect 20349 7967 20407 7973
rect 20530 7964 20536 7976
rect 20588 7964 20594 8016
rect 21168 8007 21226 8013
rect 21168 7973 21180 8007
rect 21214 8004 21226 8007
rect 21266 8004 21272 8016
rect 21214 7976 21272 8004
rect 21214 7973 21226 7976
rect 21168 7967 21226 7973
rect 21266 7964 21272 7976
rect 21324 7964 21330 8016
rect 1688 7936 1716 7964
rect 3602 7936 3608 7948
rect 1688 7908 3608 7936
rect 3602 7896 3608 7908
rect 3660 7896 3666 7948
rect 5804 7939 5862 7945
rect 5804 7905 5816 7939
rect 5850 7936 5862 7939
rect 6086 7936 6092 7948
rect 5850 7908 6092 7936
rect 5850 7905 5862 7908
rect 5804 7899 5862 7905
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 8481 7939 8539 7945
rect 8481 7905 8493 7939
rect 8527 7936 8539 7939
rect 8938 7936 8944 7948
rect 8527 7908 8944 7936
rect 8527 7905 8539 7908
rect 8481 7899 8539 7905
rect 8938 7896 8944 7908
rect 8996 7896 9002 7948
rect 10502 7936 10508 7948
rect 10463 7908 10508 7936
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 15562 7936 15568 7948
rect 14200 7908 15568 7936
rect 1670 7828 1676 7880
rect 1728 7868 1734 7880
rect 2590 7868 2596 7880
rect 1728 7840 2596 7868
rect 1728 7828 1734 7840
rect 2590 7828 2596 7840
rect 2648 7868 2654 7880
rect 2869 7871 2927 7877
rect 2869 7868 2881 7871
rect 2648 7840 2881 7868
rect 2648 7828 2654 7840
rect 2869 7837 2881 7840
rect 2915 7837 2927 7871
rect 4062 7868 4068 7880
rect 4023 7840 4068 7868
rect 2869 7831 2927 7837
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 5534 7868 5540 7880
rect 5495 7840 5540 7868
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 8665 7871 8723 7877
rect 8665 7837 8677 7871
rect 8711 7868 8723 7871
rect 8846 7868 8852 7880
rect 8711 7840 8852 7868
rect 8711 7837 8723 7840
rect 8665 7831 8723 7837
rect 8846 7828 8852 7840
rect 8904 7828 8910 7880
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 9490 7868 9496 7880
rect 9180 7840 9496 7868
rect 9180 7828 9186 7840
rect 9490 7828 9496 7840
rect 9548 7828 9554 7880
rect 10594 7868 10600 7880
rect 10555 7840 10600 7868
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 10686 7828 10692 7880
rect 10744 7868 10750 7880
rect 10744 7840 10789 7868
rect 10744 7828 10750 7840
rect 11790 7828 11796 7880
rect 11848 7868 11854 7880
rect 14200 7877 14228 7908
rect 15562 7896 15568 7908
rect 15620 7896 15626 7948
rect 15838 7896 15844 7948
rect 15896 7936 15902 7948
rect 16485 7939 16543 7945
rect 16485 7936 16497 7939
rect 15896 7908 16497 7936
rect 15896 7896 15902 7908
rect 16485 7905 16497 7908
rect 16531 7905 16543 7939
rect 16485 7899 16543 7905
rect 17589 7939 17647 7945
rect 17589 7905 17601 7939
rect 17635 7936 17647 7939
rect 17954 7936 17960 7948
rect 17635 7908 17960 7936
rect 17635 7905 17647 7908
rect 17589 7899 17647 7905
rect 17954 7896 17960 7908
rect 18012 7936 18018 7948
rect 19705 7939 19763 7945
rect 18012 7908 18276 7936
rect 18012 7896 18018 7908
rect 12161 7871 12219 7877
rect 12161 7868 12173 7871
rect 11848 7840 12173 7868
rect 11848 7828 11854 7840
rect 12161 7837 12173 7840
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 12253 7871 12311 7877
rect 12253 7837 12265 7871
rect 12299 7837 12311 7871
rect 12253 7831 12311 7837
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7868 13599 7871
rect 14185 7871 14243 7877
rect 14185 7868 14197 7871
rect 13587 7840 14197 7868
rect 13587 7837 13599 7840
rect 13541 7831 13599 7837
rect 14185 7837 14197 7840
rect 14231 7837 14243 7871
rect 16758 7868 16764 7880
rect 16719 7840 16764 7868
rect 14185 7831 14243 7837
rect 2958 7760 2964 7812
rect 3016 7800 3022 7812
rect 3697 7803 3755 7809
rect 3697 7800 3709 7803
rect 3016 7772 3709 7800
rect 3016 7760 3022 7772
rect 3697 7769 3709 7772
rect 3743 7769 3755 7803
rect 3697 7763 3755 7769
rect 7282 7760 7288 7812
rect 7340 7800 7346 7812
rect 7926 7800 7932 7812
rect 7340 7772 7932 7800
rect 7340 7760 7346 7772
rect 7926 7760 7932 7772
rect 7984 7760 7990 7812
rect 10870 7760 10876 7812
rect 10928 7800 10934 7812
rect 12268 7800 12296 7831
rect 16758 7828 16764 7840
rect 16816 7828 16822 7880
rect 18248 7877 18276 7908
rect 19705 7905 19717 7939
rect 19751 7936 19763 7939
rect 19978 7936 19984 7948
rect 19751 7908 19984 7936
rect 19751 7905 19763 7908
rect 19705 7899 19763 7905
rect 19978 7896 19984 7908
rect 20036 7896 20042 7948
rect 23768 7936 23796 8032
rect 24204 8007 24262 8013
rect 24204 7973 24216 8007
rect 24250 8004 24262 8007
rect 24486 8004 24492 8016
rect 24250 7976 24492 8004
rect 24250 7973 24262 7976
rect 24204 7967 24262 7973
rect 24486 7964 24492 7976
rect 24544 7964 24550 8016
rect 23937 7939 23995 7945
rect 23937 7936 23949 7939
rect 23768 7908 23949 7936
rect 23937 7905 23949 7908
rect 23983 7905 23995 7939
rect 23937 7899 23995 7905
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7837 18291 7871
rect 19794 7868 19800 7880
rect 19755 7840 19800 7868
rect 18233 7831 18291 7837
rect 12710 7800 12716 7812
rect 10928 7772 12716 7800
rect 10928 7760 10934 7772
rect 12710 7760 12716 7772
rect 12768 7760 12774 7812
rect 15562 7760 15568 7812
rect 15620 7800 15626 7812
rect 16117 7803 16175 7809
rect 16117 7800 16129 7803
rect 15620 7772 16129 7800
rect 15620 7760 15626 7772
rect 16117 7769 16129 7772
rect 16163 7800 16175 7803
rect 18156 7800 18184 7831
rect 19794 7828 19800 7840
rect 19852 7868 19858 7880
rect 20346 7868 20352 7880
rect 19852 7840 20352 7868
rect 19852 7828 19858 7840
rect 20346 7828 20352 7840
rect 20404 7828 20410 7880
rect 20717 7871 20775 7877
rect 20717 7837 20729 7871
rect 20763 7868 20775 7871
rect 20898 7868 20904 7880
rect 20763 7840 20904 7868
rect 20763 7837 20775 7840
rect 20717 7831 20775 7837
rect 20898 7828 20904 7840
rect 20956 7828 20962 7880
rect 16163 7772 18184 7800
rect 16163 7769 16175 7772
rect 16117 7763 16175 7769
rect 18506 7760 18512 7812
rect 18564 7800 18570 7812
rect 19245 7803 19303 7809
rect 19245 7800 19257 7803
rect 18564 7772 19257 7800
rect 18564 7760 18570 7772
rect 19245 7769 19257 7772
rect 19291 7769 19303 7803
rect 19245 7763 19303 7769
rect 1394 7692 1400 7744
rect 1452 7732 1458 7744
rect 1581 7735 1639 7741
rect 1581 7732 1593 7735
rect 1452 7704 1593 7732
rect 1452 7692 1458 7704
rect 1581 7701 1593 7704
rect 1627 7701 1639 7735
rect 1581 7695 1639 7701
rect 2866 7692 2872 7744
rect 2924 7732 2930 7744
rect 3329 7735 3387 7741
rect 3329 7732 3341 7735
rect 2924 7704 3341 7732
rect 2924 7692 2930 7704
rect 3329 7701 3341 7704
rect 3375 7701 3387 7735
rect 4522 7732 4528 7744
rect 4483 7704 4528 7732
rect 3329 7695 3387 7701
rect 4522 7692 4528 7704
rect 4580 7692 4586 7744
rect 6914 7732 6920 7744
rect 6875 7704 6920 7732
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 7558 7732 7564 7744
rect 7519 7704 7564 7732
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 8018 7732 8024 7744
rect 7979 7704 8024 7732
rect 8018 7692 8024 7704
rect 8076 7692 8082 7744
rect 9030 7732 9036 7744
rect 8991 7704 9036 7732
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 9122 7692 9128 7744
rect 9180 7732 9186 7744
rect 9401 7735 9459 7741
rect 9401 7732 9413 7735
rect 9180 7704 9413 7732
rect 9180 7692 9186 7704
rect 9401 7701 9413 7704
rect 9447 7701 9459 7735
rect 10042 7732 10048 7744
rect 10003 7704 10048 7732
rect 9401 7695 9459 7701
rect 10042 7692 10048 7704
rect 10100 7692 10106 7744
rect 11238 7732 11244 7744
rect 11199 7704 11244 7732
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 11698 7732 11704 7744
rect 11659 7704 11704 7732
rect 11698 7692 11704 7704
rect 11756 7692 11762 7744
rect 15654 7692 15660 7744
rect 15712 7732 15718 7744
rect 16025 7735 16083 7741
rect 16025 7732 16037 7735
rect 15712 7704 16037 7732
rect 15712 7692 15718 7704
rect 16025 7701 16037 7704
rect 16071 7732 16083 7735
rect 16850 7732 16856 7744
rect 16071 7704 16856 7732
rect 16071 7701 16083 7704
rect 16025 7695 16083 7701
rect 16850 7692 16856 7704
rect 16908 7692 16914 7744
rect 16942 7692 16948 7744
rect 17000 7732 17006 7744
rect 17129 7735 17187 7741
rect 17129 7732 17141 7735
rect 17000 7704 17141 7732
rect 17000 7692 17006 7704
rect 17129 7701 17141 7704
rect 17175 7701 17187 7735
rect 17129 7695 17187 7701
rect 24670 7692 24676 7744
rect 24728 7732 24734 7744
rect 25317 7735 25375 7741
rect 25317 7732 25329 7735
rect 24728 7704 25329 7732
rect 24728 7692 24734 7704
rect 25317 7701 25329 7704
rect 25363 7701 25375 7735
rect 25317 7695 25375 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1670 7528 1676 7540
rect 1631 7500 1676 7528
rect 1670 7488 1676 7500
rect 1728 7488 1734 7540
rect 3510 7528 3516 7540
rect 3471 7500 3516 7528
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 5166 7528 5172 7540
rect 5127 7500 5172 7528
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 6086 7528 6092 7540
rect 5999 7500 6092 7528
rect 6086 7488 6092 7500
rect 6144 7528 6150 7540
rect 8205 7531 8263 7537
rect 8205 7528 8217 7531
rect 6144 7500 8217 7528
rect 6144 7488 6150 7500
rect 8205 7497 8217 7500
rect 8251 7497 8263 7531
rect 10778 7528 10784 7540
rect 10739 7500 10784 7528
rect 8205 7491 8263 7497
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 11790 7528 11796 7540
rect 11751 7500 11796 7528
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 12158 7528 12164 7540
rect 12119 7500 12164 7528
rect 12158 7488 12164 7500
rect 12216 7488 12222 7540
rect 12710 7528 12716 7540
rect 12671 7500 12716 7528
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 12894 7488 12900 7540
rect 12952 7528 12958 7540
rect 13633 7531 13691 7537
rect 13633 7528 13645 7531
rect 12952 7500 13645 7528
rect 12952 7488 12958 7500
rect 13633 7497 13645 7500
rect 13679 7497 13691 7531
rect 13633 7491 13691 7497
rect 15197 7531 15255 7537
rect 15197 7497 15209 7531
rect 15243 7528 15255 7531
rect 15654 7528 15660 7540
rect 15243 7500 15660 7528
rect 15243 7497 15255 7500
rect 15197 7491 15255 7497
rect 4430 7392 4436 7404
rect 4391 7364 4436 7392
rect 4430 7352 4436 7364
rect 4488 7352 4494 7404
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7392 5135 7395
rect 5626 7392 5632 7404
rect 5123 7364 5632 7392
rect 5123 7361 5135 7364
rect 5077 7355 5135 7361
rect 5626 7352 5632 7364
rect 5684 7392 5690 7404
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5684 7364 5825 7392
rect 5684 7352 5690 7364
rect 5813 7361 5825 7364
rect 5859 7392 5871 7395
rect 6104 7392 6132 7488
rect 9677 7463 9735 7469
rect 9677 7429 9689 7463
rect 9723 7460 9735 7463
rect 10686 7460 10692 7472
rect 9723 7432 10692 7460
rect 9723 7429 9735 7432
rect 9677 7423 9735 7429
rect 10686 7420 10692 7432
rect 10744 7420 10750 7472
rect 13648 7404 13676 7491
rect 15654 7488 15660 7500
rect 15712 7488 15718 7540
rect 15838 7528 15844 7540
rect 15799 7500 15844 7528
rect 15838 7488 15844 7500
rect 15896 7528 15902 7540
rect 16206 7528 16212 7540
rect 15896 7500 16212 7528
rect 15896 7488 15902 7500
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 17402 7528 17408 7540
rect 17363 7500 17408 7528
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 18046 7528 18052 7540
rect 18007 7500 18052 7528
rect 18046 7488 18052 7500
rect 18104 7488 18110 7540
rect 19337 7531 19395 7537
rect 19337 7497 19349 7531
rect 19383 7528 19395 7531
rect 19794 7528 19800 7540
rect 19383 7500 19800 7528
rect 19383 7497 19395 7500
rect 19337 7491 19395 7497
rect 19794 7488 19800 7500
rect 19852 7488 19858 7540
rect 22189 7531 22247 7537
rect 22189 7497 22201 7531
rect 22235 7528 22247 7531
rect 22554 7528 22560 7540
rect 22235 7500 22560 7528
rect 22235 7497 22247 7500
rect 22189 7491 22247 7497
rect 15286 7420 15292 7472
rect 15344 7460 15350 7472
rect 16301 7463 16359 7469
rect 16301 7460 16313 7463
rect 15344 7432 16313 7460
rect 15344 7420 15350 7432
rect 16301 7429 16313 7432
rect 16347 7429 16359 7463
rect 16301 7423 16359 7429
rect 17310 7420 17316 7472
rect 17368 7460 17374 7472
rect 17773 7463 17831 7469
rect 17773 7460 17785 7463
rect 17368 7432 17785 7460
rect 17368 7420 17374 7432
rect 17773 7429 17785 7432
rect 17819 7460 17831 7463
rect 17819 7432 18552 7460
rect 17819 7429 17831 7432
rect 17773 7423 17831 7429
rect 5859 7364 6132 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 9766 7352 9772 7404
rect 9824 7392 9830 7404
rect 10229 7395 10287 7401
rect 10229 7392 10241 7395
rect 9824 7364 10241 7392
rect 9824 7352 9830 7364
rect 10229 7361 10241 7364
rect 10275 7392 10287 7395
rect 10502 7392 10508 7404
rect 10275 7364 10508 7392
rect 10275 7361 10287 7364
rect 10229 7355 10287 7361
rect 10502 7352 10508 7364
rect 10560 7352 10566 7404
rect 11238 7352 11244 7404
rect 11296 7392 11302 7404
rect 11333 7395 11391 7401
rect 11333 7392 11345 7395
rect 11296 7364 11345 7392
rect 11296 7352 11302 7364
rect 11333 7361 11345 7364
rect 11379 7361 11391 7395
rect 13630 7392 13636 7404
rect 13543 7364 13636 7392
rect 11333 7355 11391 7361
rect 13630 7352 13636 7364
rect 13688 7392 13694 7404
rect 13817 7395 13875 7401
rect 13817 7392 13829 7395
rect 13688 7364 13829 7392
rect 13688 7352 13694 7364
rect 13817 7361 13829 7364
rect 13863 7361 13875 7395
rect 16850 7392 16856 7404
rect 16811 7364 16856 7392
rect 13817 7355 13875 7361
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 18524 7401 18552 7432
rect 19978 7420 19984 7472
rect 20036 7460 20042 7472
rect 20717 7463 20775 7469
rect 20717 7460 20729 7463
rect 20036 7432 20729 7460
rect 20036 7420 20042 7432
rect 20717 7429 20729 7432
rect 20763 7429 20775 7463
rect 20717 7423 20775 7429
rect 18509 7395 18567 7401
rect 18509 7361 18521 7395
rect 18555 7361 18567 7395
rect 18509 7355 18567 7361
rect 18693 7395 18751 7401
rect 18693 7361 18705 7395
rect 18739 7392 18751 7395
rect 19242 7392 19248 7404
rect 18739 7364 19248 7392
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 19242 7352 19248 7364
rect 19300 7352 19306 7404
rect 21266 7392 21272 7404
rect 21227 7364 21272 7392
rect 21266 7352 21272 7364
rect 21324 7392 21330 7404
rect 22204 7392 22232 7491
rect 22554 7488 22560 7500
rect 22612 7488 22618 7540
rect 23658 7528 23664 7540
rect 23619 7500 23664 7528
rect 23658 7488 23664 7500
rect 23716 7488 23722 7540
rect 23750 7488 23756 7540
rect 23808 7528 23814 7540
rect 24673 7531 24731 7537
rect 24673 7528 24685 7531
rect 23808 7500 24685 7528
rect 23808 7488 23814 7500
rect 24673 7497 24685 7500
rect 24719 7497 24731 7531
rect 25130 7528 25136 7540
rect 25091 7500 25136 7528
rect 24673 7491 24731 7497
rect 25130 7488 25136 7500
rect 25188 7488 25194 7540
rect 25314 7488 25320 7540
rect 25372 7528 25378 7540
rect 25409 7531 25467 7537
rect 25409 7528 25421 7531
rect 25372 7500 25421 7528
rect 25372 7488 25378 7500
rect 25409 7497 25421 7500
rect 25455 7497 25467 7531
rect 25409 7491 25467 7497
rect 21324 7364 22232 7392
rect 21324 7352 21330 7364
rect 23842 7352 23848 7404
rect 23900 7392 23906 7404
rect 24121 7395 24179 7401
rect 24121 7392 24133 7395
rect 23900 7364 24133 7392
rect 23900 7352 23906 7364
rect 24121 7361 24133 7364
rect 24167 7361 24179 7395
rect 24121 7355 24179 7361
rect 24305 7395 24363 7401
rect 24305 7361 24317 7395
rect 24351 7392 24363 7395
rect 24670 7392 24676 7404
rect 24351 7364 24676 7392
rect 24351 7361 24363 7364
rect 24305 7355 24363 7361
rect 1946 7284 1952 7336
rect 2004 7324 2010 7336
rect 2041 7327 2099 7333
rect 2041 7324 2053 7327
rect 2004 7296 2053 7324
rect 2004 7284 2010 7296
rect 2041 7293 2053 7296
rect 2087 7324 2099 7327
rect 2133 7327 2191 7333
rect 2133 7324 2145 7327
rect 2087 7296 2145 7324
rect 2087 7293 2099 7296
rect 2041 7287 2099 7293
rect 2133 7293 2145 7296
rect 2179 7293 2191 7327
rect 2133 7287 2191 7293
rect 5718 7284 5724 7336
rect 5776 7324 5782 7336
rect 6181 7327 6239 7333
rect 6181 7324 6193 7327
rect 5776 7296 6193 7324
rect 5776 7284 5782 7296
rect 6181 7293 6193 7296
rect 6227 7324 6239 7327
rect 6641 7327 6699 7333
rect 6641 7324 6653 7327
rect 6227 7296 6653 7324
rect 6227 7293 6239 7296
rect 6181 7287 6239 7293
rect 6641 7293 6653 7296
rect 6687 7324 6699 7327
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6687 7296 6837 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 6825 7293 6837 7296
rect 6871 7324 6883 7327
rect 7650 7324 7656 7336
rect 6871 7296 7656 7324
rect 6871 7293 6883 7296
rect 6825 7287 6883 7293
rect 7650 7284 7656 7296
rect 7708 7284 7714 7336
rect 9674 7284 9680 7336
rect 9732 7324 9738 7336
rect 10594 7324 10600 7336
rect 9732 7296 10600 7324
rect 9732 7284 9738 7296
rect 10594 7284 10600 7296
rect 10652 7284 10658 7336
rect 11146 7284 11152 7336
rect 11204 7324 11210 7336
rect 11204 7296 11284 7324
rect 11204 7284 11210 7296
rect 2222 7216 2228 7268
rect 2280 7256 2286 7268
rect 2378 7259 2436 7265
rect 2378 7256 2390 7259
rect 2280 7228 2390 7256
rect 2280 7216 2286 7228
rect 2378 7225 2390 7228
rect 2424 7225 2436 7259
rect 2378 7219 2436 7225
rect 5537 7259 5595 7265
rect 5537 7225 5549 7259
rect 5583 7256 5595 7259
rect 5902 7256 5908 7268
rect 5583 7228 5908 7256
rect 5583 7225 5595 7228
rect 5537 7219 5595 7225
rect 5902 7216 5908 7228
rect 5960 7216 5966 7268
rect 6270 7256 6276 7268
rect 6104 7228 6276 7256
rect 2130 7148 2136 7200
rect 2188 7188 2194 7200
rect 4798 7188 4804 7200
rect 2188 7160 4804 7188
rect 2188 7148 2194 7160
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 5629 7191 5687 7197
rect 5629 7157 5641 7191
rect 5675 7188 5687 7191
rect 6104 7188 6132 7228
rect 6270 7216 6276 7228
rect 6328 7256 6334 7268
rect 6914 7256 6920 7268
rect 6328 7228 6920 7256
rect 6328 7216 6334 7228
rect 6914 7216 6920 7228
rect 6972 7216 6978 7268
rect 7098 7265 7104 7268
rect 7092 7256 7104 7265
rect 7059 7228 7104 7256
rect 7092 7219 7104 7228
rect 7098 7216 7104 7219
rect 7156 7216 7162 7268
rect 8662 7216 8668 7268
rect 8720 7256 8726 7268
rect 9125 7259 9183 7265
rect 9125 7256 9137 7259
rect 8720 7228 9137 7256
rect 8720 7216 8726 7228
rect 9125 7225 9137 7228
rect 9171 7256 9183 7259
rect 9214 7256 9220 7268
rect 9171 7228 9220 7256
rect 9171 7225 9183 7228
rect 9125 7219 9183 7225
rect 9214 7216 9220 7228
rect 9272 7216 9278 7268
rect 9769 7259 9827 7265
rect 9769 7225 9781 7259
rect 9815 7256 9827 7259
rect 10962 7256 10968 7268
rect 9815 7228 10968 7256
rect 9815 7225 9827 7228
rect 9769 7219 9827 7225
rect 10962 7216 10968 7228
rect 11020 7216 11026 7268
rect 11256 7265 11284 7296
rect 12894 7284 12900 7336
rect 12952 7324 12958 7336
rect 13446 7324 13452 7336
rect 12952 7296 13452 7324
rect 12952 7284 12958 7296
rect 13446 7284 13452 7296
rect 13504 7284 13510 7336
rect 18138 7284 18144 7336
rect 18196 7324 18202 7336
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 18196 7296 18429 7324
rect 18196 7284 18202 7296
rect 18417 7293 18429 7296
rect 18463 7293 18475 7327
rect 18417 7287 18475 7293
rect 19613 7327 19671 7333
rect 19613 7293 19625 7327
rect 19659 7324 19671 7327
rect 20254 7324 20260 7336
rect 19659 7296 20260 7324
rect 19659 7293 19671 7296
rect 19613 7287 19671 7293
rect 20254 7284 20260 7296
rect 20312 7284 20318 7336
rect 22281 7327 22339 7333
rect 22281 7293 22293 7327
rect 22327 7324 22339 7327
rect 22738 7324 22744 7336
rect 22327 7296 22744 7324
rect 22327 7293 22339 7296
rect 22281 7287 22339 7293
rect 22738 7284 22744 7296
rect 22796 7284 22802 7336
rect 23106 7324 23112 7336
rect 23019 7296 23112 7324
rect 23106 7284 23112 7296
rect 23164 7324 23170 7336
rect 24320 7324 24348 7355
rect 24670 7352 24676 7364
rect 24728 7352 24734 7404
rect 25222 7324 25228 7336
rect 23164 7296 24348 7324
rect 25183 7296 25228 7324
rect 23164 7284 23170 7296
rect 25222 7284 25228 7296
rect 25280 7324 25286 7336
rect 25777 7327 25835 7333
rect 25777 7324 25789 7327
rect 25280 7296 25789 7324
rect 25280 7284 25286 7296
rect 25777 7293 25789 7296
rect 25823 7293 25835 7327
rect 25777 7287 25835 7293
rect 11241 7259 11299 7265
rect 11241 7225 11253 7259
rect 11287 7225 11299 7259
rect 11241 7219 11299 7225
rect 13357 7259 13415 7265
rect 13357 7225 13369 7259
rect 13403 7256 13415 7259
rect 14062 7259 14120 7265
rect 14062 7256 14074 7259
rect 13403 7228 14074 7256
rect 13403 7225 13415 7228
rect 13357 7219 13415 7225
rect 14062 7225 14074 7228
rect 14108 7256 14120 7259
rect 14366 7256 14372 7268
rect 14108 7228 14372 7256
rect 14108 7225 14120 7228
rect 14062 7219 14120 7225
rect 14366 7216 14372 7228
rect 14424 7216 14430 7268
rect 18966 7256 18972 7268
rect 16684 7228 18972 7256
rect 5675 7160 6132 7188
rect 8849 7191 8907 7197
rect 5675 7157 5687 7160
rect 5629 7151 5687 7157
rect 8849 7157 8861 7191
rect 8895 7188 8907 7191
rect 8938 7188 8944 7200
rect 8895 7160 8944 7188
rect 8895 7157 8907 7160
rect 8849 7151 8907 7157
rect 8938 7148 8944 7160
rect 8996 7148 9002 7200
rect 11149 7191 11207 7197
rect 11149 7157 11161 7191
rect 11195 7188 11207 7191
rect 11698 7188 11704 7200
rect 11195 7160 11704 7188
rect 11195 7157 11207 7160
rect 11149 7151 11207 7157
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 12805 7191 12863 7197
rect 12805 7157 12817 7191
rect 12851 7188 12863 7191
rect 13538 7188 13544 7200
rect 12851 7160 13544 7188
rect 12851 7157 12863 7160
rect 12805 7151 12863 7157
rect 13538 7148 13544 7160
rect 13596 7148 13602 7200
rect 16114 7188 16120 7200
rect 16075 7160 16120 7188
rect 16114 7148 16120 7160
rect 16172 7188 16178 7200
rect 16684 7197 16712 7228
rect 18966 7216 18972 7228
rect 19024 7216 19030 7268
rect 19886 7216 19892 7268
rect 19944 7256 19950 7268
rect 20165 7259 20223 7265
rect 20165 7256 20177 7259
rect 19944 7228 20177 7256
rect 19944 7216 19950 7228
rect 20165 7225 20177 7228
rect 20211 7256 20223 7259
rect 21174 7256 21180 7268
rect 20211 7228 21180 7256
rect 20211 7225 20223 7228
rect 20165 7219 20223 7225
rect 21174 7216 21180 7228
rect 21232 7216 21238 7268
rect 23474 7256 23480 7268
rect 23435 7228 23480 7256
rect 23474 7216 23480 7228
rect 23532 7256 23538 7268
rect 24029 7259 24087 7265
rect 24029 7256 24041 7259
rect 23532 7228 24041 7256
rect 23532 7216 23538 7228
rect 24029 7225 24041 7228
rect 24075 7225 24087 7259
rect 24029 7219 24087 7225
rect 16669 7191 16727 7197
rect 16669 7188 16681 7191
rect 16172 7160 16681 7188
rect 16172 7148 16178 7160
rect 16669 7157 16681 7160
rect 16715 7157 16727 7191
rect 16669 7151 16727 7157
rect 16761 7191 16819 7197
rect 16761 7157 16773 7191
rect 16807 7188 16819 7191
rect 16850 7188 16856 7200
rect 16807 7160 16856 7188
rect 16807 7157 16819 7160
rect 16761 7151 16819 7157
rect 16850 7148 16856 7160
rect 16908 7148 16914 7200
rect 19797 7191 19855 7197
rect 19797 7157 19809 7191
rect 19843 7188 19855 7191
rect 20346 7188 20352 7200
rect 19843 7160 20352 7188
rect 19843 7157 19855 7160
rect 19797 7151 19855 7157
rect 20346 7148 20352 7160
rect 20404 7148 20410 7200
rect 20625 7191 20683 7197
rect 20625 7157 20637 7191
rect 20671 7188 20683 7191
rect 20714 7188 20720 7200
rect 20671 7160 20720 7188
rect 20671 7157 20683 7160
rect 20625 7151 20683 7157
rect 20714 7148 20720 7160
rect 20772 7188 20778 7200
rect 21085 7191 21143 7197
rect 21085 7188 21097 7191
rect 20772 7160 21097 7188
rect 20772 7148 20778 7160
rect 21085 7157 21097 7160
rect 21131 7157 21143 7191
rect 21085 7151 21143 7157
rect 21542 7148 21548 7200
rect 21600 7188 21606 7200
rect 21729 7191 21787 7197
rect 21729 7188 21741 7191
rect 21600 7160 21741 7188
rect 21600 7148 21606 7160
rect 21729 7157 21741 7160
rect 21775 7157 21787 7191
rect 21729 7151 21787 7157
rect 22465 7191 22523 7197
rect 22465 7157 22477 7191
rect 22511 7188 22523 7191
rect 23290 7188 23296 7200
rect 22511 7160 23296 7188
rect 22511 7157 22523 7160
rect 22465 7151 22523 7157
rect 23290 7148 23296 7160
rect 23348 7148 23354 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2406 6984 2412 6996
rect 2367 6956 2412 6984
rect 2406 6944 2412 6956
rect 2464 6944 2470 6996
rect 2590 6944 2596 6996
rect 2648 6984 2654 6996
rect 2777 6987 2835 6993
rect 2777 6984 2789 6987
rect 2648 6956 2789 6984
rect 2648 6944 2654 6956
rect 2777 6953 2789 6956
rect 2823 6984 2835 6987
rect 4062 6984 4068 6996
rect 2823 6956 4068 6984
rect 2823 6953 2835 6956
rect 2777 6947 2835 6953
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 5626 6984 5632 6996
rect 5587 6956 5632 6984
rect 5626 6944 5632 6956
rect 5684 6944 5690 6996
rect 5902 6984 5908 6996
rect 5815 6956 5908 6984
rect 5902 6944 5908 6956
rect 5960 6984 5966 6996
rect 6822 6984 6828 6996
rect 5960 6956 6828 6984
rect 5960 6944 5966 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 8294 6984 8300 6996
rect 8255 6956 8300 6984
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 11054 6984 11060 6996
rect 10796 6956 11060 6984
rect 3510 6916 3516 6928
rect 3471 6888 3516 6916
rect 3510 6876 3516 6888
rect 3568 6876 3574 6928
rect 4709 6919 4767 6925
rect 4709 6885 4721 6919
rect 4755 6916 4767 6919
rect 5166 6916 5172 6928
rect 4755 6888 5172 6916
rect 4755 6885 4767 6888
rect 4709 6879 4767 6885
rect 5166 6876 5172 6888
rect 5224 6876 5230 6928
rect 8110 6876 8116 6928
rect 8168 6916 8174 6928
rect 8205 6919 8263 6925
rect 8205 6916 8217 6919
rect 8168 6888 8217 6916
rect 8168 6876 8174 6888
rect 8205 6885 8217 6888
rect 8251 6885 8263 6919
rect 8205 6879 8263 6885
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 2869 6743 2927 6749
rect 3053 6783 3111 6789
rect 3053 6749 3065 6783
rect 3099 6780 3111 6783
rect 3528 6780 3556 6876
rect 6270 6848 6276 6860
rect 6231 6820 6276 6848
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 9950 6808 9956 6860
rect 10008 6848 10014 6860
rect 10796 6857 10824 6956
rect 11054 6944 11060 6956
rect 11112 6944 11118 6996
rect 11238 6944 11244 6996
rect 11296 6984 11302 6996
rect 12161 6987 12219 6993
rect 12161 6984 12173 6987
rect 11296 6956 12173 6984
rect 11296 6944 11302 6956
rect 12161 6953 12173 6956
rect 12207 6953 12219 6987
rect 13170 6984 13176 6996
rect 13131 6956 13176 6984
rect 12161 6947 12219 6953
rect 13170 6944 13176 6956
rect 13228 6984 13234 6996
rect 13725 6987 13783 6993
rect 13725 6984 13737 6987
rect 13228 6956 13737 6984
rect 13228 6944 13234 6956
rect 13725 6953 13737 6956
rect 13771 6953 13783 6987
rect 13725 6947 13783 6953
rect 14458 6944 14464 6996
rect 14516 6984 14522 6996
rect 14737 6987 14795 6993
rect 14737 6984 14749 6987
rect 14516 6956 14749 6984
rect 14516 6944 14522 6956
rect 14737 6953 14749 6956
rect 14783 6953 14795 6987
rect 15562 6984 15568 6996
rect 15523 6956 15568 6984
rect 14737 6947 14795 6953
rect 15562 6944 15568 6956
rect 15620 6944 15626 6996
rect 15933 6987 15991 6993
rect 15933 6953 15945 6987
rect 15979 6984 15991 6987
rect 16758 6984 16764 6996
rect 15979 6956 16764 6984
rect 15979 6953 15991 6956
rect 15933 6947 15991 6953
rect 16758 6944 16764 6956
rect 16816 6944 16822 6996
rect 18138 6984 18144 6996
rect 18099 6956 18144 6984
rect 18138 6944 18144 6956
rect 18196 6944 18202 6996
rect 19978 6984 19984 6996
rect 19939 6956 19984 6984
rect 19978 6944 19984 6956
rect 20036 6944 20042 6996
rect 20349 6987 20407 6993
rect 20349 6953 20361 6987
rect 20395 6984 20407 6987
rect 20622 6984 20628 6996
rect 20395 6956 20628 6984
rect 20395 6953 20407 6956
rect 20349 6947 20407 6953
rect 20622 6944 20628 6956
rect 20680 6944 20686 6996
rect 20717 6987 20775 6993
rect 20717 6953 20729 6987
rect 20763 6984 20775 6987
rect 21266 6984 21272 6996
rect 20763 6956 21272 6984
rect 20763 6953 20775 6956
rect 20717 6947 20775 6953
rect 21266 6944 21272 6956
rect 21324 6944 21330 6996
rect 22281 6987 22339 6993
rect 22281 6953 22293 6987
rect 22327 6984 22339 6987
rect 22554 6984 22560 6996
rect 22327 6956 22560 6984
rect 22327 6953 22339 6956
rect 22281 6947 22339 6953
rect 22554 6944 22560 6956
rect 22612 6944 22618 6996
rect 23661 6987 23719 6993
rect 23661 6953 23673 6987
rect 23707 6984 23719 6987
rect 23842 6984 23848 6996
rect 23707 6956 23848 6984
rect 23707 6953 23719 6956
rect 23661 6947 23719 6953
rect 23842 6944 23848 6956
rect 23900 6944 23906 6996
rect 13630 6876 13636 6928
rect 13688 6916 13694 6928
rect 14369 6919 14427 6925
rect 14369 6916 14381 6919
rect 13688 6888 14381 6916
rect 13688 6876 13694 6888
rect 14369 6885 14381 6888
rect 14415 6885 14427 6919
rect 14369 6879 14427 6885
rect 18046 6876 18052 6928
rect 18104 6916 18110 6928
rect 19426 6916 19432 6928
rect 18104 6888 19432 6916
rect 18104 6876 18110 6888
rect 19426 6876 19432 6888
rect 19484 6876 19490 6928
rect 24020 6919 24078 6925
rect 24020 6885 24032 6919
rect 24066 6916 24078 6919
rect 24670 6916 24676 6928
rect 24066 6888 24676 6916
rect 24066 6885 24078 6888
rect 24020 6879 24078 6885
rect 24670 6876 24676 6888
rect 24728 6876 24734 6928
rect 10229 6851 10287 6857
rect 10229 6848 10241 6851
rect 10008 6820 10241 6848
rect 10008 6808 10014 6820
rect 10229 6817 10241 6820
rect 10275 6817 10287 6851
rect 10229 6811 10287 6817
rect 10781 6851 10839 6857
rect 10781 6817 10793 6851
rect 10827 6817 10839 6851
rect 10781 6811 10839 6817
rect 10870 6808 10876 6860
rect 10928 6848 10934 6860
rect 16298 6857 16304 6860
rect 11037 6851 11095 6857
rect 11037 6848 11049 6851
rect 10928 6820 11049 6848
rect 10928 6808 10934 6820
rect 11037 6817 11049 6820
rect 11083 6817 11095 6851
rect 16292 6848 16304 6857
rect 16259 6820 16304 6848
rect 11037 6811 11095 6817
rect 16292 6811 16304 6820
rect 16298 6808 16304 6811
rect 16356 6808 16362 6860
rect 18874 6848 18880 6860
rect 18835 6820 18880 6848
rect 18874 6808 18880 6820
rect 18932 6808 18938 6860
rect 20622 6808 20628 6860
rect 20680 6848 20686 6860
rect 21157 6851 21215 6857
rect 21157 6848 21169 6851
rect 20680 6820 21169 6848
rect 20680 6808 20686 6820
rect 21157 6817 21169 6820
rect 21203 6817 21215 6851
rect 23750 6848 23756 6860
rect 23711 6820 23756 6848
rect 21157 6811 21215 6817
rect 23750 6808 23756 6820
rect 23808 6808 23814 6860
rect 4798 6780 4804 6792
rect 3099 6752 3556 6780
rect 4759 6752 4804 6780
rect 3099 6749 3111 6752
rect 3053 6743 3111 6749
rect 1578 6712 1584 6724
rect 1539 6684 1584 6712
rect 1578 6672 1584 6684
rect 1636 6672 1642 6724
rect 2498 6672 2504 6724
rect 2556 6712 2562 6724
rect 2884 6712 2912 6743
rect 4798 6740 4804 6752
rect 4856 6740 4862 6792
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 4948 6752 4993 6780
rect 4948 6740 4954 6752
rect 6086 6740 6092 6792
rect 6144 6780 6150 6792
rect 6365 6783 6423 6789
rect 6365 6780 6377 6783
rect 6144 6752 6377 6780
rect 6144 6740 6150 6752
rect 6365 6749 6377 6752
rect 6411 6780 6423 6783
rect 6454 6780 6460 6792
rect 6411 6752 6460 6780
rect 6411 6749 6423 6752
rect 6365 6743 6423 6749
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6749 6607 6783
rect 8478 6780 8484 6792
rect 8439 6752 8484 6780
rect 6549 6743 6607 6749
rect 3694 6712 3700 6724
rect 2556 6684 3700 6712
rect 2556 6672 2562 6684
rect 3694 6672 3700 6684
rect 3752 6672 3758 6724
rect 3970 6672 3976 6724
rect 4028 6712 4034 6724
rect 4341 6715 4399 6721
rect 4341 6712 4353 6715
rect 4028 6684 4353 6712
rect 4028 6672 4034 6684
rect 4341 6681 4353 6684
rect 4387 6681 4399 6715
rect 6564 6712 6592 6743
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 9766 6780 9772 6792
rect 9727 6752 9772 6780
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 13354 6740 13360 6792
rect 13412 6780 13418 6792
rect 13817 6783 13875 6789
rect 13817 6780 13829 6783
rect 13412 6752 13829 6780
rect 13412 6740 13418 6752
rect 13817 6749 13829 6752
rect 13863 6749 13875 6783
rect 13817 6743 13875 6749
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6749 13967 6783
rect 13909 6743 13967 6749
rect 7009 6715 7067 6721
rect 7009 6712 7021 6715
rect 6564 6684 7021 6712
rect 4341 6675 4399 6681
rect 7009 6681 7021 6684
rect 7055 6712 7067 6715
rect 7098 6712 7104 6724
rect 7055 6684 7104 6712
rect 7055 6681 7067 6684
rect 7009 6675 7067 6681
rect 7098 6672 7104 6684
rect 7156 6712 7162 6724
rect 7377 6715 7435 6721
rect 7377 6712 7389 6715
rect 7156 6684 7389 6712
rect 7156 6672 7162 6684
rect 7377 6681 7389 6684
rect 7423 6712 7435 6715
rect 7745 6715 7803 6721
rect 7745 6712 7757 6715
rect 7423 6684 7757 6712
rect 7423 6681 7435 6684
rect 7377 6675 7435 6681
rect 7745 6681 7757 6684
rect 7791 6712 7803 6715
rect 8496 6712 8524 6740
rect 8754 6712 8760 6724
rect 7791 6684 8524 6712
rect 8588 6684 8760 6712
rect 7791 6681 7803 6684
rect 7745 6675 7803 6681
rect 2222 6644 2228 6656
rect 2183 6616 2228 6644
rect 2222 6604 2228 6616
rect 2280 6604 2286 6656
rect 3786 6644 3792 6656
rect 3747 6616 3792 6644
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 7837 6647 7895 6653
rect 7837 6644 7849 6647
rect 6972 6616 7849 6644
rect 6972 6604 6978 6616
rect 7837 6613 7849 6616
rect 7883 6613 7895 6647
rect 7837 6607 7895 6613
rect 8110 6604 8116 6656
rect 8168 6644 8174 6656
rect 8588 6644 8616 6684
rect 8754 6672 8760 6684
rect 8812 6672 8818 6724
rect 12897 6715 12955 6721
rect 12897 6681 12909 6715
rect 12943 6712 12955 6715
rect 13924 6712 13952 6743
rect 15838 6740 15844 6792
rect 15896 6780 15902 6792
rect 16025 6783 16083 6789
rect 16025 6780 16037 6783
rect 15896 6752 16037 6780
rect 15896 6740 15902 6752
rect 16025 6749 16037 6752
rect 16071 6749 16083 6783
rect 16025 6743 16083 6749
rect 18690 6740 18696 6792
rect 18748 6780 18754 6792
rect 18969 6783 19027 6789
rect 18969 6780 18981 6783
rect 18748 6752 18981 6780
rect 18748 6740 18754 6752
rect 18969 6749 18981 6752
rect 19015 6749 19027 6783
rect 18969 6743 19027 6749
rect 19058 6740 19064 6792
rect 19116 6780 19122 6792
rect 20898 6780 20904 6792
rect 19116 6752 19161 6780
rect 20811 6752 20904 6780
rect 19116 6740 19122 6752
rect 20898 6740 20904 6752
rect 20956 6740 20962 6792
rect 14090 6712 14096 6724
rect 12943 6684 14096 6712
rect 12943 6681 12955 6684
rect 12897 6675 12955 6681
rect 14090 6672 14096 6684
rect 14148 6672 14154 6724
rect 8846 6644 8852 6656
rect 8168 6616 8616 6644
rect 8807 6616 8852 6644
rect 8168 6604 8174 6616
rect 8846 6604 8852 6616
rect 8904 6604 8910 6656
rect 9214 6644 9220 6656
rect 9175 6616 9220 6644
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 10689 6647 10747 6653
rect 10689 6613 10701 6647
rect 10735 6644 10747 6647
rect 11054 6644 11060 6656
rect 10735 6616 11060 6644
rect 10735 6613 10747 6616
rect 10689 6607 10747 6613
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 13170 6604 13176 6656
rect 13228 6644 13234 6656
rect 13357 6647 13415 6653
rect 13357 6644 13369 6647
rect 13228 6616 13369 6644
rect 13228 6604 13234 6616
rect 13357 6613 13369 6616
rect 13403 6644 13415 6647
rect 13814 6644 13820 6656
rect 13403 6616 13820 6644
rect 13403 6613 13415 6616
rect 13357 6607 13415 6613
rect 13814 6604 13820 6616
rect 13872 6604 13878 6656
rect 17402 6644 17408 6656
rect 17363 6616 17408 6644
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 18506 6644 18512 6656
rect 18467 6616 18512 6644
rect 18506 6604 18512 6616
rect 18564 6604 18570 6656
rect 19610 6644 19616 6656
rect 19571 6616 19616 6644
rect 19610 6604 19616 6616
rect 19668 6604 19674 6656
rect 20916 6644 20944 6740
rect 21542 6644 21548 6656
rect 20916 6616 21548 6644
rect 21542 6604 21548 6616
rect 21600 6604 21606 6656
rect 22738 6604 22744 6656
rect 22796 6644 22802 6656
rect 22833 6647 22891 6653
rect 22833 6644 22845 6647
rect 22796 6616 22845 6644
rect 22796 6604 22802 6616
rect 22833 6613 22845 6616
rect 22879 6613 22891 6647
rect 25130 6644 25136 6656
rect 25091 6616 25136 6644
rect 22833 6607 22891 6613
rect 25130 6604 25136 6616
rect 25188 6604 25194 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2498 6440 2504 6452
rect 2459 6412 2504 6440
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 2832 6412 2877 6440
rect 2832 6400 2838 6412
rect 3602 6400 3608 6452
rect 3660 6440 3666 6452
rect 3789 6443 3847 6449
rect 3789 6440 3801 6443
rect 3660 6412 3801 6440
rect 3660 6400 3666 6412
rect 3789 6409 3801 6412
rect 3835 6440 3847 6443
rect 4065 6443 4123 6449
rect 4065 6440 4077 6443
rect 3835 6412 4077 6440
rect 3835 6409 3847 6412
rect 3789 6403 3847 6409
rect 4065 6409 4077 6412
rect 4111 6409 4123 6443
rect 4065 6403 4123 6409
rect 5997 6443 6055 6449
rect 5997 6409 6009 6443
rect 6043 6440 6055 6443
rect 6086 6440 6092 6452
rect 6043 6412 6092 6440
rect 6043 6409 6055 6412
rect 5997 6403 6055 6409
rect 6086 6400 6092 6412
rect 6144 6400 6150 6452
rect 6270 6440 6276 6452
rect 6231 6412 6276 6440
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 8478 6400 8484 6452
rect 8536 6440 8542 6452
rect 9493 6443 9551 6449
rect 9493 6440 9505 6443
rect 8536 6412 9505 6440
rect 8536 6400 8542 6412
rect 9493 6409 9505 6412
rect 9539 6409 9551 6443
rect 9493 6403 9551 6409
rect 10686 6400 10692 6452
rect 10744 6440 10750 6452
rect 13078 6440 13084 6452
rect 10744 6412 13084 6440
rect 10744 6400 10750 6412
rect 13078 6400 13084 6412
rect 13136 6400 13142 6452
rect 13354 6440 13360 6452
rect 13315 6412 13360 6440
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 14366 6400 14372 6452
rect 14424 6440 14430 6452
rect 15105 6443 15163 6449
rect 15105 6440 15117 6443
rect 14424 6412 15117 6440
rect 14424 6400 14430 6412
rect 15105 6409 15117 6412
rect 15151 6409 15163 6443
rect 15105 6403 15163 6409
rect 17402 6400 17408 6452
rect 17460 6440 17466 6452
rect 17497 6443 17555 6449
rect 17497 6440 17509 6443
rect 17460 6412 17509 6440
rect 17460 6400 17466 6412
rect 17497 6409 17509 6412
rect 17543 6440 17555 6443
rect 17865 6443 17923 6449
rect 17865 6440 17877 6443
rect 17543 6412 17877 6440
rect 17543 6409 17555 6412
rect 17497 6403 17555 6409
rect 17865 6409 17877 6412
rect 17911 6440 17923 6443
rect 19058 6440 19064 6452
rect 17911 6412 19064 6440
rect 17911 6409 17923 6412
rect 17865 6403 17923 6409
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 23106 6440 23112 6452
rect 23067 6412 23112 6440
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 23477 6443 23535 6449
rect 23477 6409 23489 6443
rect 23523 6440 23535 6443
rect 23750 6440 23756 6452
rect 23523 6412 23756 6440
rect 23523 6409 23535 6412
rect 23477 6403 23535 6409
rect 23750 6400 23756 6412
rect 23808 6440 23814 6452
rect 23937 6443 23995 6449
rect 23937 6440 23949 6443
rect 23808 6412 23949 6440
rect 23808 6400 23814 6412
rect 23937 6409 23949 6412
rect 23983 6409 23995 6443
rect 23937 6403 23995 6409
rect 2133 6375 2191 6381
rect 2133 6341 2145 6375
rect 2179 6372 2191 6375
rect 2590 6372 2596 6384
rect 2179 6344 2596 6372
rect 2179 6341 2191 6344
rect 2133 6335 2191 6341
rect 2590 6332 2596 6344
rect 2648 6332 2654 6384
rect 4341 6375 4399 6381
rect 4341 6372 4353 6375
rect 3252 6344 4353 6372
rect 3252 6316 3280 6344
rect 4341 6341 4353 6344
rect 4387 6341 4399 6375
rect 4341 6335 4399 6341
rect 4798 6332 4804 6384
rect 4856 6372 4862 6384
rect 5353 6375 5411 6381
rect 5353 6372 5365 6375
rect 4856 6344 5365 6372
rect 4856 6332 4862 6344
rect 5353 6341 5365 6344
rect 5399 6372 5411 6375
rect 5442 6372 5448 6384
rect 5399 6344 5448 6372
rect 5399 6341 5411 6344
rect 5353 6335 5411 6341
rect 5442 6332 5448 6344
rect 5500 6332 5506 6384
rect 3234 6304 3240 6316
rect 3195 6276 3240 6304
rect 3234 6264 3240 6276
rect 3292 6264 3298 6316
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6304 3479 6307
rect 3510 6304 3516 6316
rect 3467 6276 3516 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 4890 6304 4896 6316
rect 4851 6276 4896 6304
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 6288 6304 6316 6400
rect 9766 6332 9772 6384
rect 9824 6372 9830 6384
rect 10321 6375 10379 6381
rect 10321 6372 10333 6375
rect 9824 6344 10333 6372
rect 9824 6332 9830 6344
rect 10321 6341 10333 6344
rect 10367 6372 10379 6375
rect 10413 6375 10471 6381
rect 10413 6372 10425 6375
rect 10367 6344 10425 6372
rect 10367 6341 10379 6344
rect 10321 6335 10379 6341
rect 10413 6341 10425 6344
rect 10459 6341 10471 6375
rect 10413 6335 10471 6341
rect 10962 6332 10968 6384
rect 11020 6372 11026 6384
rect 11609 6375 11667 6381
rect 11609 6372 11621 6375
rect 11020 6344 11621 6372
rect 11020 6332 11026 6344
rect 11609 6341 11621 6344
rect 11655 6372 11667 6375
rect 12710 6372 12716 6384
rect 11655 6344 12716 6372
rect 11655 6341 11667 6344
rect 11609 6335 11667 6341
rect 12710 6332 12716 6344
rect 12768 6372 12774 6384
rect 12768 6344 13768 6372
rect 12768 6332 12774 6344
rect 13740 6313 13768 6344
rect 6825 6307 6883 6313
rect 6825 6304 6837 6307
rect 6288 6276 6837 6304
rect 6825 6273 6837 6276
rect 6871 6273 6883 6307
rect 11149 6307 11207 6313
rect 11149 6304 11161 6307
rect 6825 6267 6883 6273
rect 10060 6276 11161 6304
rect 3145 6239 3203 6245
rect 3145 6205 3157 6239
rect 3191 6236 3203 6239
rect 3970 6236 3976 6248
rect 3191 6208 3976 6236
rect 3191 6205 3203 6208
rect 3145 6199 3203 6205
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6236 4307 6239
rect 4706 6236 4712 6248
rect 4295 6208 4712 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 8018 6196 8024 6248
rect 8076 6236 8082 6248
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 8076 6208 8125 6236
rect 8076 6196 8082 6208
rect 8113 6205 8125 6208
rect 8159 6205 8171 6239
rect 8113 6199 8171 6205
rect 4065 6171 4123 6177
rect 4065 6137 4077 6171
rect 4111 6168 4123 6171
rect 4801 6171 4859 6177
rect 4801 6168 4813 6171
rect 4111 6140 4813 6168
rect 4111 6137 4123 6140
rect 4065 6131 4123 6137
rect 4801 6137 4813 6140
rect 4847 6168 4859 6171
rect 7558 6168 7564 6180
rect 4847 6140 7564 6168
rect 4847 6137 4859 6140
rect 4801 6131 4859 6137
rect 7558 6128 7564 6140
rect 7616 6128 7622 6180
rect 8386 6177 8392 6180
rect 7653 6171 7711 6177
rect 7653 6137 7665 6171
rect 7699 6168 7711 6171
rect 8380 6168 8392 6177
rect 7699 6140 8392 6168
rect 7699 6137 7711 6140
rect 7653 6131 7711 6137
rect 8380 6131 8392 6140
rect 8386 6128 8392 6131
rect 8444 6128 8450 6180
rect 1397 6103 1455 6109
rect 1397 6069 1409 6103
rect 1443 6100 1455 6103
rect 1578 6100 1584 6112
rect 1443 6072 1584 6100
rect 1443 6069 1455 6072
rect 1397 6063 1455 6069
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 8018 6100 8024 6112
rect 7979 6072 8024 6100
rect 8018 6060 8024 6072
rect 8076 6060 8082 6112
rect 8846 6060 8852 6112
rect 8904 6100 8910 6112
rect 10060 6109 10088 6276
rect 11149 6273 11161 6276
rect 11195 6273 11207 6307
rect 11149 6267 11207 6273
rect 13725 6307 13783 6313
rect 13725 6273 13737 6307
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 10321 6239 10379 6245
rect 10321 6205 10333 6239
rect 10367 6236 10379 6239
rect 10778 6236 10784 6248
rect 10367 6208 10784 6236
rect 10367 6205 10379 6208
rect 10321 6199 10379 6205
rect 10778 6196 10784 6208
rect 10836 6236 10842 6248
rect 11057 6239 11115 6245
rect 11057 6236 11069 6239
rect 10836 6208 11069 6236
rect 10836 6196 10842 6208
rect 11057 6205 11069 6208
rect 11103 6205 11115 6239
rect 11057 6199 11115 6205
rect 12253 6239 12311 6245
rect 12253 6205 12265 6239
rect 12299 6236 12311 6239
rect 12526 6236 12532 6248
rect 12299 6208 12532 6236
rect 12299 6205 12311 6208
rect 12253 6199 12311 6205
rect 12526 6196 12532 6208
rect 12584 6236 12590 6248
rect 12621 6239 12679 6245
rect 12621 6236 12633 6239
rect 12584 6208 12633 6236
rect 12584 6196 12590 6208
rect 12621 6205 12633 6208
rect 12667 6205 12679 6239
rect 13740 6236 13768 6267
rect 16482 6264 16488 6316
rect 16540 6304 16546 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16540 6276 16865 6304
rect 16540 6264 16546 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 17034 6304 17040 6316
rect 16947 6276 17040 6304
rect 16853 6267 16911 6273
rect 17034 6264 17040 6276
rect 17092 6304 17098 6316
rect 17420 6304 17448 6400
rect 18690 6372 18696 6384
rect 18651 6344 18696 6372
rect 18690 6332 18696 6344
rect 18748 6332 18754 6384
rect 17092 6276 17448 6304
rect 22649 6307 22707 6313
rect 17092 6264 17098 6276
rect 22649 6273 22661 6307
rect 22695 6304 22707 6307
rect 22738 6304 22744 6316
rect 22695 6276 22744 6304
rect 22695 6273 22707 6276
rect 22649 6267 22707 6273
rect 22738 6264 22744 6276
rect 22796 6264 22802 6316
rect 23952 6304 23980 6403
rect 24121 6307 24179 6313
rect 24121 6304 24133 6307
rect 23952 6276 24133 6304
rect 24121 6273 24133 6276
rect 24167 6273 24179 6307
rect 24121 6267 24179 6273
rect 15838 6236 15844 6248
rect 13740 6208 15844 6236
rect 12621 6199 12679 6205
rect 15838 6196 15844 6208
rect 15896 6196 15902 6248
rect 18141 6239 18199 6245
rect 18141 6205 18153 6239
rect 18187 6236 18199 6239
rect 18322 6236 18328 6248
rect 18187 6208 18328 6236
rect 18187 6205 18199 6208
rect 18141 6199 18199 6205
rect 18322 6196 18328 6208
rect 18380 6196 18386 6248
rect 19245 6239 19303 6245
rect 19245 6205 19257 6239
rect 19291 6205 19303 6239
rect 19245 6199 19303 6205
rect 13992 6171 14050 6177
rect 13992 6137 14004 6171
rect 14038 6168 14050 6171
rect 14090 6168 14096 6180
rect 14038 6140 14096 6168
rect 14038 6137 14050 6140
rect 13992 6131 14050 6137
rect 14090 6128 14096 6140
rect 14148 6128 14154 6180
rect 16301 6171 16359 6177
rect 16301 6137 16313 6171
rect 16347 6168 16359 6171
rect 16347 6140 16804 6168
rect 16347 6137 16359 6140
rect 16301 6131 16359 6137
rect 10045 6103 10103 6109
rect 10045 6100 10057 6103
rect 8904 6072 10057 6100
rect 8904 6060 8910 6072
rect 10045 6069 10057 6072
rect 10091 6069 10103 6103
rect 10045 6063 10103 6069
rect 10597 6103 10655 6109
rect 10597 6069 10609 6103
rect 10643 6100 10655 6103
rect 10686 6100 10692 6112
rect 10643 6072 10692 6100
rect 10643 6069 10655 6072
rect 10597 6063 10655 6069
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 10965 6103 11023 6109
rect 10965 6069 10977 6103
rect 11011 6100 11023 6103
rect 11054 6100 11060 6112
rect 11011 6072 11060 6100
rect 11011 6069 11023 6072
rect 10965 6063 11023 6069
rect 11054 6060 11060 6072
rect 11112 6060 11118 6112
rect 12805 6103 12863 6109
rect 12805 6069 12817 6103
rect 12851 6100 12863 6103
rect 13538 6100 13544 6112
rect 12851 6072 13544 6100
rect 12851 6069 12863 6072
rect 12805 6063 12863 6069
rect 13538 6060 13544 6072
rect 13596 6060 13602 6112
rect 16393 6103 16451 6109
rect 16393 6069 16405 6103
rect 16439 6100 16451 6103
rect 16574 6100 16580 6112
rect 16439 6072 16580 6100
rect 16439 6069 16451 6072
rect 16393 6063 16451 6069
rect 16574 6060 16580 6072
rect 16632 6060 16638 6112
rect 16776 6109 16804 6140
rect 17770 6128 17776 6180
rect 17828 6168 17834 6180
rect 19061 6171 19119 6177
rect 19061 6168 19073 6171
rect 17828 6140 19073 6168
rect 17828 6128 17834 6140
rect 19061 6137 19073 6140
rect 19107 6168 19119 6171
rect 19260 6168 19288 6199
rect 21726 6196 21732 6248
rect 21784 6236 21790 6248
rect 22373 6239 22431 6245
rect 22373 6236 22385 6239
rect 21784 6208 22385 6236
rect 21784 6196 21790 6208
rect 22373 6205 22385 6208
rect 22419 6205 22431 6239
rect 22373 6199 22431 6205
rect 22465 6239 22523 6245
rect 22465 6205 22477 6239
rect 22511 6236 22523 6239
rect 23382 6236 23388 6248
rect 22511 6208 23388 6236
rect 22511 6205 22523 6208
rect 22465 6199 22523 6205
rect 19107 6140 19288 6168
rect 19512 6171 19570 6177
rect 19107 6137 19119 6140
rect 19061 6131 19119 6137
rect 19512 6137 19524 6171
rect 19558 6168 19570 6171
rect 19610 6168 19616 6180
rect 19558 6140 19616 6168
rect 19558 6137 19570 6140
rect 19512 6131 19570 6137
rect 19610 6128 19616 6140
rect 19668 6168 19674 6180
rect 19978 6168 19984 6180
rect 19668 6140 19984 6168
rect 19668 6128 19674 6140
rect 19978 6128 19984 6140
rect 20036 6128 20042 6180
rect 21545 6171 21603 6177
rect 21545 6137 21557 6171
rect 21591 6168 21603 6171
rect 22480 6168 22508 6199
rect 23382 6196 23388 6208
rect 23440 6196 23446 6248
rect 24394 6245 24400 6248
rect 24388 6236 24400 6245
rect 24307 6208 24400 6236
rect 24388 6199 24400 6208
rect 24452 6236 24458 6248
rect 25130 6236 25136 6248
rect 24452 6208 25136 6236
rect 24394 6196 24400 6199
rect 24452 6196 24458 6208
rect 25130 6196 25136 6208
rect 25188 6196 25194 6248
rect 21591 6140 22508 6168
rect 21591 6137 21603 6140
rect 21545 6131 21603 6137
rect 16761 6103 16819 6109
rect 16761 6069 16773 6103
rect 16807 6100 16819 6103
rect 16850 6100 16856 6112
rect 16807 6072 16856 6100
rect 16807 6069 16819 6072
rect 16761 6063 16819 6069
rect 16850 6060 16856 6072
rect 16908 6060 16914 6112
rect 18325 6103 18383 6109
rect 18325 6069 18337 6103
rect 18371 6100 18383 6103
rect 18414 6100 18420 6112
rect 18371 6072 18420 6100
rect 18371 6069 18383 6072
rect 18325 6063 18383 6069
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 20622 6100 20628 6112
rect 20583 6072 20628 6100
rect 20622 6060 20628 6072
rect 20680 6060 20686 6112
rect 21726 6060 21732 6112
rect 21784 6100 21790 6112
rect 21821 6103 21879 6109
rect 21821 6100 21833 6103
rect 21784 6072 21833 6100
rect 21784 6060 21790 6072
rect 21821 6069 21833 6072
rect 21867 6069 21879 6103
rect 21821 6063 21879 6069
rect 21910 6060 21916 6112
rect 21968 6100 21974 6112
rect 22005 6103 22063 6109
rect 22005 6100 22017 6103
rect 21968 6072 22017 6100
rect 21968 6060 21974 6072
rect 22005 6069 22017 6072
rect 22051 6069 22063 6103
rect 22005 6063 22063 6069
rect 25130 6060 25136 6112
rect 25188 6100 25194 6112
rect 25501 6103 25559 6109
rect 25501 6100 25513 6103
rect 25188 6072 25513 6100
rect 25188 6060 25194 6072
rect 25501 6069 25513 6072
rect 25547 6069 25559 6103
rect 25501 6063 25559 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1578 5896 1584 5908
rect 1539 5868 1584 5896
rect 1578 5856 1584 5868
rect 1636 5856 1642 5908
rect 2317 5899 2375 5905
rect 2317 5865 2329 5899
rect 2363 5896 2375 5899
rect 2406 5896 2412 5908
rect 2363 5868 2412 5896
rect 2363 5865 2375 5868
rect 2317 5859 2375 5865
rect 2406 5856 2412 5868
rect 2464 5896 2470 5908
rect 2682 5896 2688 5908
rect 2464 5868 2688 5896
rect 2464 5856 2470 5868
rect 2682 5856 2688 5868
rect 2740 5856 2746 5908
rect 3421 5899 3479 5905
rect 3421 5865 3433 5899
rect 3467 5896 3479 5899
rect 3510 5896 3516 5908
rect 3467 5868 3516 5896
rect 3467 5865 3479 5868
rect 3421 5859 3479 5865
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 3878 5856 3884 5908
rect 3936 5896 3942 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 3936 5868 4077 5896
rect 3936 5856 3942 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 4246 5856 4252 5908
rect 4304 5896 4310 5908
rect 4525 5899 4583 5905
rect 4525 5896 4537 5899
rect 4304 5868 4537 5896
rect 4304 5856 4310 5868
rect 4525 5865 4537 5868
rect 4571 5865 4583 5899
rect 4525 5859 4583 5865
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5629 5899 5687 5905
rect 5629 5896 5641 5899
rect 5592 5868 5641 5896
rect 5592 5856 5598 5868
rect 5629 5865 5641 5868
rect 5675 5896 5687 5899
rect 6362 5896 6368 5908
rect 5675 5868 6368 5896
rect 5675 5865 5687 5868
rect 5629 5859 5687 5865
rect 6362 5856 6368 5868
rect 6420 5856 6426 5908
rect 8021 5899 8079 5905
rect 8021 5865 8033 5899
rect 8067 5896 8079 5899
rect 8202 5896 8208 5908
rect 8067 5868 8208 5896
rect 8067 5865 8079 5868
rect 8021 5859 8079 5865
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 9677 5899 9735 5905
rect 9677 5865 9689 5899
rect 9723 5896 9735 5899
rect 9858 5896 9864 5908
rect 9723 5868 9864 5896
rect 9723 5865 9735 5868
rect 9677 5859 9735 5865
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 10870 5896 10876 5908
rect 10831 5868 10876 5896
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 11330 5896 11336 5908
rect 11291 5868 11336 5896
rect 11330 5856 11336 5868
rect 11388 5856 11394 5908
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 12529 5899 12587 5905
rect 12529 5896 12541 5899
rect 12492 5868 12541 5896
rect 12492 5856 12498 5868
rect 12529 5865 12541 5868
rect 12575 5896 12587 5899
rect 13722 5896 13728 5908
rect 12575 5868 13728 5896
rect 12575 5865 12587 5868
rect 12529 5859 12587 5865
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 14090 5896 14096 5908
rect 14051 5868 14096 5896
rect 14090 5856 14096 5868
rect 14148 5896 14154 5908
rect 14645 5899 14703 5905
rect 14645 5896 14657 5899
rect 14148 5868 14657 5896
rect 14148 5856 14154 5868
rect 14645 5865 14657 5868
rect 14691 5865 14703 5899
rect 14645 5859 14703 5865
rect 14734 5856 14740 5908
rect 14792 5896 14798 5908
rect 15013 5899 15071 5905
rect 15013 5896 15025 5899
rect 14792 5868 15025 5896
rect 14792 5856 14798 5868
rect 15013 5865 15025 5868
rect 15059 5865 15071 5899
rect 15013 5859 15071 5865
rect 16117 5899 16175 5905
rect 16117 5865 16129 5899
rect 16163 5896 16175 5899
rect 16298 5896 16304 5908
rect 16163 5868 16304 5896
rect 16163 5865 16175 5868
rect 16117 5859 16175 5865
rect 2222 5788 2228 5840
rect 2280 5828 2286 5840
rect 3789 5831 3847 5837
rect 3789 5828 3801 5831
rect 2280 5800 3801 5828
rect 2280 5788 2286 5800
rect 3789 5797 3801 5800
rect 3835 5828 3847 5831
rect 4890 5828 4896 5840
rect 3835 5800 4896 5828
rect 3835 5797 3847 5800
rect 3789 5791 3847 5797
rect 4890 5788 4896 5800
rect 4948 5788 4954 5840
rect 5997 5831 6055 5837
rect 5997 5797 6009 5831
rect 6043 5828 6055 5831
rect 6270 5828 6276 5840
rect 6043 5800 6276 5828
rect 6043 5797 6055 5800
rect 5997 5791 6055 5797
rect 6270 5788 6276 5800
rect 6328 5828 6334 5840
rect 6730 5828 6736 5840
rect 6328 5800 6736 5828
rect 6328 5788 6334 5800
rect 6730 5788 6736 5800
rect 6788 5788 6794 5840
rect 8110 5788 8116 5840
rect 8168 5828 8174 5840
rect 8389 5831 8447 5837
rect 8389 5828 8401 5831
rect 8168 5800 8401 5828
rect 8168 5788 8174 5800
rect 8389 5797 8401 5800
rect 8435 5797 8447 5831
rect 8389 5791 8447 5797
rect 12980 5831 13038 5837
rect 12980 5797 12992 5831
rect 13026 5828 13038 5831
rect 13170 5828 13176 5840
rect 13026 5800 13176 5828
rect 13026 5797 13038 5800
rect 12980 5791 13038 5797
rect 13170 5788 13176 5800
rect 13228 5788 13234 5840
rect 2682 5760 2688 5772
rect 2643 5732 2688 5760
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 4062 5720 4068 5772
rect 4120 5760 4126 5772
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 4120 5732 4445 5760
rect 4120 5720 4126 5732
rect 4433 5729 4445 5732
rect 4479 5729 4491 5763
rect 5166 5760 5172 5772
rect 5079 5732 5172 5760
rect 4433 5723 4491 5729
rect 5166 5720 5172 5732
rect 5224 5760 5230 5772
rect 7742 5760 7748 5772
rect 5224 5732 7748 5760
rect 5224 5720 5230 5732
rect 7742 5720 7748 5732
rect 7800 5720 7806 5772
rect 10042 5760 10048 5772
rect 10003 5732 10048 5760
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 10870 5760 10876 5772
rect 10152 5732 10876 5760
rect 2498 5652 2504 5704
rect 2556 5692 2562 5704
rect 2777 5695 2835 5701
rect 2777 5692 2789 5695
rect 2556 5664 2789 5692
rect 2556 5652 2562 5664
rect 2777 5661 2789 5664
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 6086 5692 6092 5704
rect 6047 5664 6092 5692
rect 4709 5655 4767 5661
rect 1854 5584 1860 5636
rect 1912 5624 1918 5636
rect 1949 5627 2007 5633
rect 1949 5624 1961 5627
rect 1912 5596 1961 5624
rect 1912 5584 1918 5596
rect 1949 5593 1961 5596
rect 1995 5624 2007 5627
rect 2884 5624 2912 5655
rect 1995 5596 2912 5624
rect 4724 5624 4752 5655
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 6273 5695 6331 5701
rect 6273 5661 6285 5695
rect 6319 5692 6331 5695
rect 6730 5692 6736 5704
rect 6319 5664 6736 5692
rect 6319 5661 6331 5664
rect 6273 5655 6331 5661
rect 5258 5624 5264 5636
rect 4724 5596 5264 5624
rect 1995 5593 2007 5596
rect 1949 5587 2007 5593
rect 5258 5584 5264 5596
rect 5316 5624 5322 5636
rect 5537 5627 5595 5633
rect 5537 5624 5549 5627
rect 5316 5596 5549 5624
rect 5316 5584 5322 5596
rect 5537 5593 5549 5596
rect 5583 5624 5595 5627
rect 6288 5624 6316 5655
rect 6730 5652 6736 5664
rect 6788 5652 6794 5704
rect 6917 5695 6975 5701
rect 6917 5661 6929 5695
rect 6963 5692 6975 5695
rect 7098 5692 7104 5704
rect 6963 5664 7104 5692
rect 6963 5661 6975 5664
rect 6917 5655 6975 5661
rect 7098 5652 7104 5664
rect 7156 5652 7162 5704
rect 8481 5695 8539 5701
rect 8481 5692 8493 5695
rect 7208 5664 8493 5692
rect 7208 5624 7236 5664
rect 8481 5661 8493 5664
rect 8527 5692 8539 5695
rect 8570 5692 8576 5704
rect 8527 5664 8576 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 8570 5652 8576 5664
rect 8628 5652 8634 5704
rect 8665 5695 8723 5701
rect 8665 5661 8677 5695
rect 8711 5661 8723 5695
rect 8665 5655 8723 5661
rect 5583 5596 6316 5624
rect 6380 5596 7236 5624
rect 7929 5627 7987 5633
rect 5583 5593 5595 5596
rect 5537 5587 5595 5593
rect 3418 5516 3424 5568
rect 3476 5556 3482 5568
rect 6380 5556 6408 5596
rect 7929 5593 7941 5627
rect 7975 5624 7987 5627
rect 8386 5624 8392 5636
rect 7975 5596 8392 5624
rect 7975 5593 7987 5596
rect 7929 5587 7987 5593
rect 8386 5584 8392 5596
rect 8444 5624 8450 5636
rect 8680 5624 8708 5655
rect 8754 5652 8760 5704
rect 8812 5692 8818 5704
rect 9674 5692 9680 5704
rect 8812 5664 9680 5692
rect 8812 5652 8818 5664
rect 9674 5652 9680 5664
rect 9732 5692 9738 5704
rect 10152 5701 10180 5732
rect 10870 5720 10876 5732
rect 10928 5720 10934 5772
rect 11606 5760 11612 5772
rect 11567 5732 11612 5760
rect 11606 5720 11612 5732
rect 11664 5720 11670 5772
rect 11974 5720 11980 5772
rect 12032 5760 12038 5772
rect 14182 5760 14188 5772
rect 12032 5732 14188 5760
rect 12032 5720 12038 5732
rect 14182 5720 14188 5732
rect 14240 5720 14246 5772
rect 15028 5760 15056 5859
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 16482 5896 16488 5908
rect 16443 5868 16488 5896
rect 16482 5856 16488 5868
rect 16540 5856 16546 5908
rect 18785 5899 18843 5905
rect 18785 5865 18797 5899
rect 18831 5896 18843 5899
rect 18874 5896 18880 5908
rect 18831 5868 18880 5896
rect 18831 5865 18843 5868
rect 18785 5859 18843 5865
rect 18874 5856 18880 5868
rect 18932 5856 18938 5908
rect 18966 5856 18972 5908
rect 19024 5896 19030 5908
rect 19061 5899 19119 5905
rect 19061 5896 19073 5899
rect 19024 5868 19073 5896
rect 19024 5856 19030 5868
rect 19061 5865 19073 5868
rect 19107 5865 19119 5899
rect 19061 5859 19119 5865
rect 17034 5837 17040 5840
rect 17028 5828 17040 5837
rect 16995 5800 17040 5828
rect 17028 5791 17040 5800
rect 17034 5788 17040 5791
rect 17092 5788 17098 5840
rect 19076 5828 19104 5859
rect 19518 5856 19524 5908
rect 19576 5896 19582 5908
rect 19705 5899 19763 5905
rect 19705 5896 19717 5899
rect 19576 5868 19717 5896
rect 19576 5856 19582 5868
rect 19705 5865 19717 5868
rect 19751 5865 19763 5899
rect 21542 5896 21548 5908
rect 21503 5868 21548 5896
rect 19705 5859 19763 5865
rect 21542 5856 21548 5868
rect 21600 5856 21606 5908
rect 22005 5899 22063 5905
rect 22005 5865 22017 5899
rect 22051 5896 22063 5899
rect 22094 5896 22100 5908
rect 22051 5868 22100 5896
rect 22051 5865 22063 5868
rect 22005 5859 22063 5865
rect 19613 5831 19671 5837
rect 19613 5828 19625 5831
rect 19076 5800 19625 5828
rect 19613 5797 19625 5800
rect 19659 5797 19671 5831
rect 19613 5791 19671 5797
rect 15289 5763 15347 5769
rect 15289 5760 15301 5763
rect 15028 5732 15301 5760
rect 15289 5729 15301 5732
rect 15335 5729 15347 5763
rect 15289 5723 15347 5729
rect 15838 5720 15844 5772
rect 15896 5760 15902 5772
rect 16761 5763 16819 5769
rect 16761 5760 16773 5763
rect 15896 5732 16773 5760
rect 15896 5720 15902 5732
rect 16761 5729 16773 5732
rect 16807 5760 16819 5763
rect 16850 5760 16856 5772
rect 16807 5732 16856 5760
rect 16807 5729 16819 5732
rect 16761 5723 16819 5729
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 18322 5720 18328 5772
rect 18380 5760 18386 5772
rect 20257 5763 20315 5769
rect 20257 5760 20269 5763
rect 18380 5732 20269 5760
rect 18380 5720 18386 5732
rect 20257 5729 20269 5732
rect 20303 5729 20315 5763
rect 20257 5723 20315 5729
rect 20993 5763 21051 5769
rect 20993 5729 21005 5763
rect 21039 5760 21051 5763
rect 22020 5760 22048 5859
rect 22094 5856 22100 5868
rect 22152 5856 22158 5908
rect 24121 5899 24179 5905
rect 24121 5865 24133 5899
rect 24167 5896 24179 5899
rect 24394 5896 24400 5908
rect 24167 5868 24400 5896
rect 24167 5865 24179 5868
rect 24121 5859 24179 5865
rect 24394 5856 24400 5868
rect 24452 5896 24458 5908
rect 24670 5896 24676 5908
rect 24452 5868 24676 5896
rect 24452 5856 24458 5868
rect 24670 5856 24676 5868
rect 24728 5856 24734 5908
rect 24946 5896 24952 5908
rect 24907 5868 24952 5896
rect 24946 5856 24952 5868
rect 25004 5856 25010 5908
rect 23750 5828 23756 5840
rect 22112 5800 23756 5828
rect 22112 5769 22140 5800
rect 23750 5788 23756 5800
rect 23808 5788 23814 5840
rect 22370 5769 22376 5772
rect 21039 5732 22048 5760
rect 22097 5763 22155 5769
rect 21039 5729 21051 5732
rect 20993 5723 21051 5729
rect 22097 5729 22109 5763
rect 22143 5729 22155 5763
rect 22364 5760 22376 5769
rect 22331 5732 22376 5760
rect 22097 5723 22155 5729
rect 22364 5723 22376 5732
rect 10137 5695 10195 5701
rect 10137 5692 10149 5695
rect 9732 5664 10149 5692
rect 9732 5652 9738 5664
rect 10137 5661 10149 5664
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10321 5695 10379 5701
rect 10321 5661 10333 5695
rect 10367 5692 10379 5695
rect 10778 5692 10784 5704
rect 10367 5664 10784 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 10336 5624 10364 5655
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 12710 5692 12716 5704
rect 12671 5664 12716 5692
rect 12710 5652 12716 5664
rect 12768 5652 12774 5704
rect 19886 5692 19892 5704
rect 19847 5664 19892 5692
rect 19886 5652 19892 5664
rect 19944 5652 19950 5704
rect 8444 5596 10364 5624
rect 8444 5584 8450 5596
rect 22002 5584 22008 5636
rect 22060 5624 22066 5636
rect 22112 5624 22140 5723
rect 22370 5720 22376 5723
rect 22428 5720 22434 5772
rect 24762 5652 24768 5704
rect 24820 5692 24826 5704
rect 25041 5695 25099 5701
rect 25041 5692 25053 5695
rect 24820 5664 25053 5692
rect 24820 5652 24826 5664
rect 25041 5661 25053 5664
rect 25087 5661 25099 5695
rect 25041 5655 25099 5661
rect 25130 5652 25136 5704
rect 25188 5692 25194 5704
rect 25188 5664 25233 5692
rect 25188 5652 25194 5664
rect 22060 5596 22140 5624
rect 22060 5584 22066 5596
rect 23934 5584 23940 5636
rect 23992 5624 23998 5636
rect 24581 5627 24639 5633
rect 24581 5624 24593 5627
rect 23992 5596 24593 5624
rect 23992 5584 23998 5596
rect 24581 5593 24593 5596
rect 24627 5593 24639 5627
rect 24581 5587 24639 5593
rect 3476 5528 6408 5556
rect 3476 5516 3482 5528
rect 6914 5516 6920 5568
rect 6972 5556 6978 5568
rect 7193 5559 7251 5565
rect 7193 5556 7205 5559
rect 6972 5528 7205 5556
rect 6972 5516 6978 5528
rect 7193 5525 7205 5528
rect 7239 5525 7251 5559
rect 9398 5556 9404 5568
rect 9359 5528 9404 5556
rect 7193 5519 7251 5525
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 11698 5516 11704 5568
rect 11756 5556 11762 5568
rect 11793 5559 11851 5565
rect 11793 5556 11805 5559
rect 11756 5528 11805 5556
rect 11756 5516 11762 5528
rect 11793 5525 11805 5528
rect 11839 5525 11851 5559
rect 11793 5519 11851 5525
rect 12894 5516 12900 5568
rect 12952 5556 12958 5568
rect 13722 5556 13728 5568
rect 12952 5528 13728 5556
rect 12952 5516 12958 5528
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 15473 5559 15531 5565
rect 15473 5525 15485 5559
rect 15519 5556 15531 5559
rect 15930 5556 15936 5568
rect 15519 5528 15936 5556
rect 15519 5525 15531 5528
rect 15473 5519 15531 5525
rect 15930 5516 15936 5528
rect 15988 5516 15994 5568
rect 18138 5556 18144 5568
rect 18099 5528 18144 5556
rect 18138 5516 18144 5528
rect 18196 5516 18202 5568
rect 19245 5559 19303 5565
rect 19245 5525 19257 5559
rect 19291 5556 19303 5559
rect 19334 5556 19340 5568
rect 19291 5528 19340 5556
rect 19291 5525 19303 5528
rect 19245 5519 19303 5525
rect 19334 5516 19340 5528
rect 19392 5516 19398 5568
rect 20622 5556 20628 5568
rect 20583 5528 20628 5556
rect 20622 5516 20628 5528
rect 20680 5516 20686 5568
rect 21177 5559 21235 5565
rect 21177 5525 21189 5559
rect 21223 5556 21235 5559
rect 21450 5556 21456 5568
rect 21223 5528 21456 5556
rect 21223 5525 21235 5528
rect 21177 5519 21235 5525
rect 21450 5516 21456 5528
rect 21508 5516 21514 5568
rect 22738 5516 22744 5568
rect 22796 5556 22802 5568
rect 23477 5559 23535 5565
rect 23477 5556 23489 5559
rect 22796 5528 23489 5556
rect 22796 5516 22802 5528
rect 23477 5525 23489 5528
rect 23523 5525 23535 5559
rect 23477 5519 23535 5525
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1397 5355 1455 5361
rect 1397 5321 1409 5355
rect 1443 5352 1455 5355
rect 2222 5352 2228 5364
rect 1443 5324 2228 5352
rect 1443 5321 1455 5324
rect 1397 5315 1455 5321
rect 2222 5312 2228 5324
rect 2280 5352 2286 5364
rect 2958 5352 2964 5364
rect 2280 5324 2964 5352
rect 2280 5312 2286 5324
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 3789 5355 3847 5361
rect 3789 5352 3801 5355
rect 3252 5324 3801 5352
rect 1854 5176 1860 5228
rect 1912 5216 1918 5228
rect 3252 5225 3280 5324
rect 3789 5321 3801 5324
rect 3835 5352 3847 5355
rect 4062 5352 4068 5364
rect 3835 5324 4068 5352
rect 3835 5321 3847 5324
rect 3789 5315 3847 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4157 5355 4215 5361
rect 4157 5321 4169 5355
rect 4203 5352 4215 5355
rect 4246 5352 4252 5364
rect 4203 5324 4252 5352
rect 4203 5321 4215 5324
rect 4157 5315 4215 5321
rect 4246 5312 4252 5324
rect 4304 5312 4310 5364
rect 5350 5312 5356 5364
rect 5408 5352 5414 5364
rect 5629 5355 5687 5361
rect 5629 5352 5641 5355
rect 5408 5324 5641 5352
rect 5408 5312 5414 5324
rect 5629 5321 5641 5324
rect 5675 5352 5687 5355
rect 7098 5352 7104 5364
rect 5675 5324 7104 5352
rect 5675 5321 5687 5324
rect 5629 5315 5687 5321
rect 7098 5312 7104 5324
rect 7156 5312 7162 5364
rect 10870 5312 10876 5364
rect 10928 5352 10934 5364
rect 11241 5355 11299 5361
rect 11241 5352 11253 5355
rect 10928 5324 11253 5352
rect 10928 5312 10934 5324
rect 11241 5321 11253 5324
rect 11287 5321 11299 5355
rect 11241 5315 11299 5321
rect 12802 5312 12808 5364
rect 12860 5352 12866 5364
rect 13449 5355 13507 5361
rect 12860 5324 13308 5352
rect 12860 5312 12866 5324
rect 8294 5244 8300 5296
rect 8352 5284 8358 5296
rect 8757 5287 8815 5293
rect 8757 5284 8769 5287
rect 8352 5256 8769 5284
rect 8352 5244 8358 5256
rect 8757 5253 8769 5256
rect 8803 5284 8815 5287
rect 9214 5284 9220 5296
rect 8803 5256 9220 5284
rect 8803 5253 8815 5256
rect 8757 5247 8815 5253
rect 9214 5244 9220 5256
rect 9272 5244 9278 5296
rect 10689 5287 10747 5293
rect 10689 5253 10701 5287
rect 10735 5284 10747 5287
rect 12161 5287 12219 5293
rect 12161 5284 12173 5287
rect 10735 5256 12173 5284
rect 10735 5253 10747 5256
rect 10689 5247 10747 5253
rect 12161 5253 12173 5256
rect 12207 5284 12219 5287
rect 13170 5284 13176 5296
rect 12207 5256 13176 5284
rect 12207 5253 12219 5256
rect 12161 5247 12219 5253
rect 13170 5244 13176 5256
rect 13228 5244 13234 5296
rect 13280 5284 13308 5324
rect 13449 5321 13461 5355
rect 13495 5352 13507 5355
rect 14366 5352 14372 5364
rect 13495 5324 14372 5352
rect 13495 5321 13507 5324
rect 13449 5315 13507 5321
rect 13541 5287 13599 5293
rect 13541 5284 13553 5287
rect 13280 5256 13553 5284
rect 13541 5253 13553 5256
rect 13587 5253 13599 5287
rect 13541 5247 13599 5253
rect 1949 5219 2007 5225
rect 1949 5216 1961 5219
rect 1912 5188 1961 5216
rect 1912 5176 1918 5188
rect 1949 5185 1961 5188
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5185 3295 5219
rect 3237 5179 3295 5185
rect 12710 5176 12716 5228
rect 12768 5216 12774 5228
rect 12989 5219 13047 5225
rect 12989 5216 13001 5219
rect 12768 5188 13001 5216
rect 12768 5176 12774 5188
rect 12989 5185 13001 5188
rect 13035 5185 13047 5219
rect 13998 5216 14004 5228
rect 13959 5188 14004 5216
rect 12989 5179 13047 5185
rect 1578 5108 1584 5160
rect 1636 5148 1642 5160
rect 1765 5151 1823 5157
rect 1765 5148 1777 5151
rect 1636 5120 1777 5148
rect 1636 5108 1642 5120
rect 1765 5117 1777 5120
rect 1811 5117 1823 5151
rect 4246 5148 4252 5160
rect 4207 5120 4252 5148
rect 1765 5111 1823 5117
rect 4246 5108 4252 5120
rect 4304 5148 4310 5160
rect 7098 5157 7104 5160
rect 6549 5151 6607 5157
rect 6549 5148 6561 5151
rect 4304 5120 6561 5148
rect 4304 5108 4310 5120
rect 6549 5117 6561 5120
rect 6595 5148 6607 5151
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6595 5120 6837 5148
rect 6595 5117 6607 5120
rect 6549 5111 6607 5117
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 7092 5148 7104 5157
rect 7059 5120 7104 5148
rect 6825 5111 6883 5117
rect 7092 5111 7104 5120
rect 1394 5040 1400 5092
rect 1452 5080 1458 5092
rect 2409 5083 2467 5089
rect 2409 5080 2421 5083
rect 1452 5052 2421 5080
rect 1452 5040 1458 5052
rect 2409 5049 2421 5052
rect 2455 5080 2467 5083
rect 2498 5080 2504 5092
rect 2455 5052 2504 5080
rect 2455 5049 2467 5052
rect 2409 5043 2467 5049
rect 2498 5040 2504 5052
rect 2556 5040 2562 5092
rect 4516 5083 4574 5089
rect 4516 5049 4528 5083
rect 4562 5080 4574 5083
rect 5258 5080 5264 5092
rect 4562 5052 5264 5080
rect 4562 5049 4574 5052
rect 4516 5043 4574 5049
rect 5258 5040 5264 5052
rect 5316 5040 5322 5092
rect 6840 5080 6868 5111
rect 7098 5108 7104 5111
rect 7156 5108 7162 5160
rect 8478 5148 8484 5160
rect 8128 5120 8484 5148
rect 8018 5080 8024 5092
rect 6840 5052 8024 5080
rect 8018 5040 8024 5052
rect 8076 5080 8082 5092
rect 8128 5080 8156 5120
rect 8478 5108 8484 5120
rect 8536 5148 8542 5160
rect 9214 5148 9220 5160
rect 8536 5120 9220 5148
rect 8536 5108 8542 5120
rect 9214 5108 9220 5120
rect 9272 5148 9278 5160
rect 9309 5151 9367 5157
rect 9309 5148 9321 5151
rect 9272 5120 9321 5148
rect 9272 5108 9278 5120
rect 9309 5117 9321 5120
rect 9355 5117 9367 5151
rect 9309 5111 9367 5117
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 13004 5148 13032 5179
rect 13998 5176 14004 5188
rect 14056 5176 14062 5228
rect 14108 5225 14136 5324
rect 14366 5312 14372 5324
rect 14424 5312 14430 5364
rect 16850 5312 16856 5364
rect 16908 5352 16914 5364
rect 17037 5355 17095 5361
rect 17037 5352 17049 5355
rect 16908 5324 17049 5352
rect 16908 5312 16914 5324
rect 17037 5321 17049 5324
rect 17083 5352 17095 5355
rect 17770 5352 17776 5364
rect 17083 5324 17776 5352
rect 17083 5321 17095 5324
rect 17037 5315 17095 5321
rect 17770 5312 17776 5324
rect 17828 5352 17834 5364
rect 17828 5324 18092 5352
rect 17828 5312 17834 5324
rect 18064 5225 18092 5324
rect 19518 5312 19524 5364
rect 19576 5352 19582 5364
rect 19981 5355 20039 5361
rect 19981 5352 19993 5355
rect 19576 5324 19993 5352
rect 19576 5312 19582 5324
rect 19981 5321 19993 5324
rect 20027 5321 20039 5355
rect 19981 5315 20039 5321
rect 20438 5312 20444 5364
rect 20496 5352 20502 5364
rect 21542 5352 21548 5364
rect 20496 5324 21548 5352
rect 20496 5312 20502 5324
rect 21542 5312 21548 5324
rect 21600 5312 21606 5364
rect 22922 5312 22928 5364
rect 22980 5352 22986 5364
rect 23017 5355 23075 5361
rect 23017 5352 23029 5355
rect 22980 5324 23029 5352
rect 22980 5312 22986 5324
rect 23017 5321 23029 5324
rect 23063 5321 23075 5355
rect 23017 5315 23075 5321
rect 23937 5355 23995 5361
rect 23937 5321 23949 5355
rect 23983 5352 23995 5355
rect 24397 5355 24455 5361
rect 24397 5352 24409 5355
rect 23983 5324 24409 5352
rect 23983 5321 23995 5324
rect 23937 5315 23995 5321
rect 24397 5321 24409 5324
rect 24443 5352 24455 5355
rect 24762 5352 24768 5364
rect 24443 5324 24768 5352
rect 24443 5321 24455 5324
rect 24397 5315 24455 5321
rect 24762 5312 24768 5324
rect 24820 5312 24826 5364
rect 24946 5312 24952 5364
rect 25004 5352 25010 5364
rect 25409 5355 25467 5361
rect 25409 5352 25421 5355
rect 25004 5324 25421 5352
rect 25004 5312 25010 5324
rect 25409 5321 25421 5324
rect 25455 5321 25467 5355
rect 25409 5315 25467 5321
rect 19058 5244 19064 5296
rect 19116 5284 19122 5296
rect 19429 5287 19487 5293
rect 19429 5284 19441 5287
rect 19116 5256 19441 5284
rect 19116 5244 19122 5256
rect 19429 5253 19441 5256
rect 19475 5284 19487 5287
rect 24210 5284 24216 5296
rect 19475 5256 19932 5284
rect 24171 5256 24216 5284
rect 19475 5253 19487 5256
rect 19429 5247 19487 5253
rect 19904 5228 19932 5256
rect 24210 5244 24216 5256
rect 24268 5244 24274 5296
rect 14093 5219 14151 5225
rect 14093 5185 14105 5219
rect 14139 5185 14151 5219
rect 14093 5179 14151 5185
rect 18049 5219 18107 5225
rect 18049 5185 18061 5219
rect 18095 5185 18107 5219
rect 18049 5179 18107 5185
rect 19886 5176 19892 5228
rect 19944 5216 19950 5228
rect 21177 5219 21235 5225
rect 21177 5216 21189 5219
rect 19944 5188 21189 5216
rect 19944 5176 19950 5188
rect 21177 5185 21189 5188
rect 21223 5216 21235 5219
rect 21545 5219 21603 5225
rect 21545 5216 21557 5219
rect 21223 5188 21557 5216
rect 21223 5185 21235 5188
rect 21177 5179 21235 5185
rect 21545 5185 21557 5188
rect 21591 5185 21603 5219
rect 21545 5179 21603 5185
rect 24670 5176 24676 5228
rect 24728 5216 24734 5228
rect 24949 5219 25007 5225
rect 24949 5216 24961 5219
rect 24728 5188 24961 5216
rect 24728 5176 24734 5188
rect 24949 5185 24961 5188
rect 24995 5185 25007 5219
rect 24949 5179 25007 5185
rect 14921 5151 14979 5157
rect 14921 5148 14933 5151
rect 12492 5120 12537 5148
rect 13004 5120 14933 5148
rect 12492 5108 12498 5120
rect 14921 5117 14933 5120
rect 14967 5148 14979 5151
rect 15105 5151 15163 5157
rect 15105 5148 15117 5151
rect 14967 5120 15117 5148
rect 14967 5117 14979 5120
rect 14921 5111 14979 5117
rect 15105 5117 15117 5120
rect 15151 5117 15163 5151
rect 15105 5111 15163 5117
rect 18138 5108 18144 5160
rect 18196 5148 18202 5160
rect 18305 5151 18363 5157
rect 18305 5148 18317 5151
rect 18196 5120 18317 5148
rect 18196 5108 18202 5120
rect 18305 5117 18317 5120
rect 18351 5117 18363 5151
rect 20901 5151 20959 5157
rect 20901 5148 20913 5151
rect 18305 5111 18363 5117
rect 20364 5120 20913 5148
rect 9398 5080 9404 5092
rect 8076 5052 8156 5080
rect 8220 5052 9404 5080
rect 8076 5040 8082 5052
rect 8220 5024 8248 5052
rect 9398 5040 9404 5052
rect 9456 5080 9462 5092
rect 9554 5083 9612 5089
rect 9554 5080 9566 5083
rect 9456 5052 9566 5080
rect 9456 5040 9462 5052
rect 9554 5049 9566 5052
rect 9600 5049 9612 5083
rect 9554 5043 9612 5049
rect 13814 5040 13820 5092
rect 13872 5080 13878 5092
rect 13909 5083 13967 5089
rect 13909 5080 13921 5083
rect 13872 5052 13921 5080
rect 13872 5040 13878 5052
rect 13909 5049 13921 5052
rect 13955 5049 13967 5083
rect 13909 5043 13967 5049
rect 14645 5083 14703 5089
rect 14645 5049 14657 5083
rect 14691 5080 14703 5083
rect 15350 5083 15408 5089
rect 15350 5080 15362 5083
rect 14691 5052 15362 5080
rect 14691 5049 14703 5052
rect 14645 5043 14703 5049
rect 15350 5049 15362 5052
rect 15396 5080 15408 5083
rect 15838 5080 15844 5092
rect 15396 5052 15844 5080
rect 15396 5049 15408 5052
rect 15350 5043 15408 5049
rect 15838 5040 15844 5052
rect 15896 5040 15902 5092
rect 17494 5080 17500 5092
rect 17407 5052 17500 5080
rect 17494 5040 17500 5052
rect 17552 5080 17558 5092
rect 18156 5080 18184 5108
rect 17552 5052 18184 5080
rect 17552 5040 17558 5052
rect 1486 4972 1492 5024
rect 1544 5012 1550 5024
rect 1857 5015 1915 5021
rect 1857 5012 1869 5015
rect 1544 4984 1869 5012
rect 1544 4972 1550 4984
rect 1857 4981 1869 4984
rect 1903 4981 1915 5015
rect 1857 4975 1915 4981
rect 2682 4972 2688 5024
rect 2740 5012 2746 5024
rect 2774 5012 2780 5024
rect 2740 4984 2780 5012
rect 2740 4972 2746 4984
rect 2774 4972 2780 4984
rect 2832 5012 2838 5024
rect 2869 5015 2927 5021
rect 2869 5012 2881 5015
rect 2832 4984 2881 5012
rect 2832 4972 2838 4984
rect 2869 4981 2881 4984
rect 2915 5012 2927 5015
rect 4062 5012 4068 5024
rect 2915 4984 4068 5012
rect 2915 4981 2927 4984
rect 2869 4975 2927 4981
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 5166 4972 5172 5024
rect 5224 5012 5230 5024
rect 6086 5012 6092 5024
rect 5224 4984 6092 5012
rect 5224 4972 5230 4984
rect 6086 4972 6092 4984
rect 6144 5012 6150 5024
rect 6181 5015 6239 5021
rect 6181 5012 6193 5015
rect 6144 4984 6193 5012
rect 6144 4972 6150 4984
rect 6181 4981 6193 4984
rect 6227 4981 6239 5015
rect 8202 5012 8208 5024
rect 8163 4984 8208 5012
rect 6181 4975 6239 4981
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 8570 4972 8576 5024
rect 8628 5012 8634 5024
rect 9030 5012 9036 5024
rect 8628 4984 9036 5012
rect 8628 4972 8634 4984
rect 9030 4972 9036 4984
rect 9088 5012 9094 5024
rect 9125 5015 9183 5021
rect 9125 5012 9137 5015
rect 9088 4984 9137 5012
rect 9088 4972 9094 4984
rect 9125 4981 9137 4984
rect 9171 4981 9183 5015
rect 9125 4975 9183 4981
rect 11885 5015 11943 5021
rect 11885 4981 11897 5015
rect 11931 5012 11943 5015
rect 12434 5012 12440 5024
rect 11931 4984 12440 5012
rect 11931 4981 11943 4984
rect 11885 4975 11943 4981
rect 12434 4972 12440 4984
rect 12492 4972 12498 5024
rect 12621 5015 12679 5021
rect 12621 4981 12633 5015
rect 12667 5012 12679 5015
rect 12986 5012 12992 5024
rect 12667 4984 12992 5012
rect 12667 4981 12679 4984
rect 12621 4975 12679 4981
rect 12986 4972 12992 4984
rect 13044 4972 13050 5024
rect 16482 5012 16488 5024
rect 16443 4984 16488 5012
rect 16482 4972 16488 4984
rect 16540 4972 16546 5024
rect 20254 4972 20260 5024
rect 20312 5012 20318 5024
rect 20364 5021 20392 5120
rect 20901 5117 20913 5120
rect 20947 5148 20959 5151
rect 21726 5148 21732 5160
rect 20947 5120 21732 5148
rect 20947 5117 20959 5120
rect 20901 5111 20959 5117
rect 21726 5108 21732 5120
rect 21784 5108 21790 5160
rect 22465 5151 22523 5157
rect 22465 5117 22477 5151
rect 22511 5148 22523 5151
rect 22922 5148 22928 5160
rect 22511 5120 22928 5148
rect 22511 5117 22523 5120
rect 22465 5111 22523 5117
rect 22922 5108 22928 5120
rect 22980 5108 22986 5160
rect 24854 5148 24860 5160
rect 24815 5120 24860 5148
rect 24854 5108 24860 5120
rect 24912 5108 24918 5160
rect 20438 5040 20444 5092
rect 20496 5080 20502 5092
rect 20993 5083 21051 5089
rect 20993 5080 21005 5083
rect 20496 5052 21005 5080
rect 20496 5040 20502 5052
rect 20993 5049 21005 5052
rect 21039 5049 21051 5083
rect 20993 5043 21051 5049
rect 24210 5040 24216 5092
rect 24268 5080 24274 5092
rect 24765 5083 24823 5089
rect 24765 5080 24777 5083
rect 24268 5052 24777 5080
rect 24268 5040 24274 5052
rect 24765 5049 24777 5052
rect 24811 5049 24823 5083
rect 24765 5043 24823 5049
rect 20349 5015 20407 5021
rect 20349 5012 20361 5015
rect 20312 4984 20361 5012
rect 20312 4972 20318 4984
rect 20349 4981 20361 4984
rect 20395 4981 20407 5015
rect 20530 5012 20536 5024
rect 20491 4984 20536 5012
rect 20349 4975 20407 4981
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 22002 4972 22008 5024
rect 22060 5012 22066 5024
rect 22097 5015 22155 5021
rect 22097 5012 22109 5015
rect 22060 4984 22109 5012
rect 22060 4972 22066 4984
rect 22097 4981 22109 4984
rect 22143 4981 22155 5015
rect 22646 5012 22652 5024
rect 22607 4984 22652 5012
rect 22097 4975 22155 4981
rect 22646 4972 22652 4984
rect 22704 4972 22710 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1486 4768 1492 4820
rect 1544 4808 1550 4820
rect 1581 4811 1639 4817
rect 1581 4808 1593 4811
rect 1544 4780 1593 4808
rect 1544 4768 1550 4780
rect 1581 4777 1593 4780
rect 1627 4777 1639 4811
rect 2038 4808 2044 4820
rect 1999 4780 2044 4808
rect 1581 4771 1639 4777
rect 2038 4768 2044 4780
rect 2096 4768 2102 4820
rect 2406 4808 2412 4820
rect 2367 4780 2412 4808
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 5169 4811 5227 4817
rect 5169 4808 5181 4811
rect 4212 4780 5181 4808
rect 4212 4768 4218 4780
rect 5169 4777 5181 4780
rect 5215 4777 5227 4811
rect 5169 4771 5227 4777
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5442 4808 5448 4820
rect 5307 4780 5448 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 6362 4808 6368 4820
rect 6323 4780 6368 4808
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 6638 4768 6644 4820
rect 6696 4808 6702 4820
rect 6733 4811 6791 4817
rect 6733 4808 6745 4811
rect 6696 4780 6745 4808
rect 6696 4768 6702 4780
rect 6733 4777 6745 4780
rect 6779 4777 6791 4811
rect 7926 4808 7932 4820
rect 7887 4780 7932 4808
rect 6733 4771 6791 4777
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 9309 4811 9367 4817
rect 9309 4808 9321 4811
rect 9272 4780 9321 4808
rect 9272 4768 9278 4780
rect 9309 4777 9321 4780
rect 9355 4777 9367 4811
rect 9309 4771 9367 4777
rect 10689 4811 10747 4817
rect 10689 4777 10701 4811
rect 10735 4808 10747 4811
rect 10778 4808 10784 4820
rect 10735 4780 10784 4808
rect 10735 4777 10747 4780
rect 10689 4771 10747 4777
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 12526 4808 12532 4820
rect 12487 4780 12532 4808
rect 12526 4768 12532 4780
rect 12584 4808 12590 4820
rect 12802 4808 12808 4820
rect 12584 4780 12808 4808
rect 12584 4768 12590 4780
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 13633 4811 13691 4817
rect 13633 4777 13645 4811
rect 13679 4808 13691 4811
rect 13998 4808 14004 4820
rect 13679 4780 14004 4808
rect 13679 4777 13691 4780
rect 13633 4771 13691 4777
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 14642 4768 14648 4820
rect 14700 4808 14706 4820
rect 15013 4811 15071 4817
rect 15013 4808 15025 4811
rect 14700 4780 15025 4808
rect 14700 4768 14706 4780
rect 15013 4777 15025 4780
rect 15059 4808 15071 4811
rect 15749 4811 15807 4817
rect 15749 4808 15761 4811
rect 15059 4780 15761 4808
rect 15059 4777 15071 4780
rect 15013 4771 15071 4777
rect 15749 4777 15761 4780
rect 15795 4777 15807 4811
rect 15749 4771 15807 4777
rect 16022 4768 16028 4820
rect 16080 4808 16086 4820
rect 16301 4811 16359 4817
rect 16301 4808 16313 4811
rect 16080 4780 16313 4808
rect 16080 4768 16086 4780
rect 16301 4777 16313 4780
rect 16347 4808 16359 4811
rect 16482 4808 16488 4820
rect 16347 4780 16488 4808
rect 16347 4777 16359 4780
rect 16301 4771 16359 4777
rect 16482 4768 16488 4780
rect 16540 4768 16546 4820
rect 16761 4811 16819 4817
rect 16761 4777 16773 4811
rect 16807 4808 16819 4811
rect 17034 4808 17040 4820
rect 16807 4780 17040 4808
rect 16807 4777 16819 4780
rect 16761 4771 16819 4777
rect 17034 4768 17040 4780
rect 17092 4768 17098 4820
rect 17221 4811 17279 4817
rect 17221 4777 17233 4811
rect 17267 4808 17279 4811
rect 17957 4811 18015 4817
rect 17957 4808 17969 4811
rect 17267 4780 17969 4808
rect 17267 4777 17279 4780
rect 17221 4771 17279 4777
rect 17957 4777 17969 4780
rect 18003 4808 18015 4811
rect 18506 4808 18512 4820
rect 18003 4780 18512 4808
rect 18003 4777 18015 4780
rect 17957 4771 18015 4777
rect 18506 4768 18512 4780
rect 18564 4768 18570 4820
rect 19150 4808 19156 4820
rect 19111 4780 19156 4808
rect 19150 4768 19156 4780
rect 19208 4768 19214 4820
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 19521 4811 19579 4817
rect 19521 4808 19533 4811
rect 19392 4780 19533 4808
rect 19392 4768 19398 4780
rect 19521 4777 19533 4780
rect 19567 4808 19579 4811
rect 20165 4811 20223 4817
rect 20165 4808 20177 4811
rect 19567 4780 20177 4808
rect 19567 4777 19579 4780
rect 19521 4771 19579 4777
rect 20165 4777 20177 4780
rect 20211 4777 20223 4811
rect 20165 4771 20223 4777
rect 20438 4768 20444 4820
rect 20496 4808 20502 4820
rect 20625 4811 20683 4817
rect 20625 4808 20637 4811
rect 20496 4780 20637 4808
rect 20496 4768 20502 4780
rect 20625 4777 20637 4780
rect 20671 4777 20683 4811
rect 20625 4771 20683 4777
rect 20806 4768 20812 4820
rect 20864 4808 20870 4820
rect 20901 4811 20959 4817
rect 20901 4808 20913 4811
rect 20864 4780 20913 4808
rect 20864 4768 20870 4780
rect 20901 4777 20913 4780
rect 20947 4777 20959 4811
rect 20901 4771 20959 4777
rect 21269 4811 21327 4817
rect 21269 4777 21281 4811
rect 21315 4808 21327 4811
rect 21634 4808 21640 4820
rect 21315 4780 21640 4808
rect 21315 4777 21327 4780
rect 21269 4771 21327 4777
rect 21634 4768 21640 4780
rect 21692 4768 21698 4820
rect 22189 4811 22247 4817
rect 22189 4777 22201 4811
rect 22235 4808 22247 4811
rect 22370 4808 22376 4820
rect 22235 4780 22376 4808
rect 22235 4777 22247 4780
rect 22189 4771 22247 4777
rect 22370 4768 22376 4780
rect 22428 4768 22434 4820
rect 24489 4811 24547 4817
rect 24489 4777 24501 4811
rect 24535 4808 24547 4811
rect 24762 4808 24768 4820
rect 24535 4780 24768 4808
rect 24535 4777 24547 4780
rect 24489 4771 24547 4777
rect 24762 4768 24768 4780
rect 24820 4768 24826 4820
rect 2501 4743 2559 4749
rect 2501 4709 2513 4743
rect 2547 4740 2559 4743
rect 3786 4740 3792 4752
rect 2547 4712 3792 4740
rect 2547 4709 2559 4712
rect 2501 4703 2559 4709
rect 3786 4700 3792 4712
rect 3844 4740 3850 4752
rect 3844 4712 5580 4740
rect 3844 4700 3850 4712
rect 5552 4684 5580 4712
rect 6546 4700 6552 4752
rect 6604 4740 6610 4752
rect 6825 4743 6883 4749
rect 6825 4740 6837 4743
rect 6604 4712 6837 4740
rect 6604 4700 6610 4712
rect 6825 4709 6837 4712
rect 6871 4709 6883 4743
rect 6825 4703 6883 4709
rect 7190 4700 7196 4752
rect 7248 4740 7254 4752
rect 8018 4740 8024 4752
rect 7248 4712 8024 4740
rect 7248 4700 7254 4712
rect 8018 4700 8024 4712
rect 8076 4740 8082 4752
rect 8389 4743 8447 4749
rect 8389 4740 8401 4743
rect 8076 4712 8401 4740
rect 8076 4700 8082 4712
rect 8389 4709 8401 4712
rect 8435 4709 8447 4743
rect 8389 4703 8447 4709
rect 11238 4700 11244 4752
rect 11296 4740 11302 4752
rect 11394 4743 11452 4749
rect 11394 4740 11406 4743
rect 11296 4712 11406 4740
rect 11296 4700 11302 4712
rect 11394 4709 11406 4712
rect 11440 4709 11452 4743
rect 11394 4703 11452 4709
rect 11514 4700 11520 4752
rect 11572 4700 11578 4752
rect 13906 4700 13912 4752
rect 13964 4740 13970 4752
rect 14093 4743 14151 4749
rect 14093 4740 14105 4743
rect 13964 4712 14105 4740
rect 13964 4700 13970 4712
rect 14093 4709 14105 4712
rect 14139 4709 14151 4743
rect 14093 4703 14151 4709
rect 16574 4700 16580 4752
rect 16632 4740 16638 4752
rect 17313 4743 17371 4749
rect 17313 4740 17325 4743
rect 16632 4712 17325 4740
rect 16632 4700 16638 4712
rect 17313 4709 17325 4712
rect 17359 4740 17371 4743
rect 17402 4740 17408 4752
rect 17359 4712 17408 4740
rect 17359 4709 17371 4712
rect 17313 4703 17371 4709
rect 17402 4700 17408 4712
rect 17460 4700 17466 4752
rect 19058 4740 19064 4752
rect 19019 4712 19064 4740
rect 19058 4700 19064 4712
rect 19116 4700 19122 4752
rect 19613 4743 19671 4749
rect 19613 4709 19625 4743
rect 19659 4740 19671 4743
rect 20530 4740 20536 4752
rect 19659 4712 20536 4740
rect 19659 4709 19671 4712
rect 19613 4703 19671 4709
rect 3881 4675 3939 4681
rect 3881 4641 3893 4675
rect 3927 4672 3939 4675
rect 4709 4675 4767 4681
rect 4709 4672 4721 4675
rect 3927 4644 4721 4672
rect 3927 4641 3939 4644
rect 3881 4635 3939 4641
rect 4709 4641 4721 4644
rect 4755 4672 4767 4675
rect 5258 4672 5264 4684
rect 4755 4644 5264 4672
rect 4755 4641 4767 4644
rect 4709 4635 4767 4641
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 5534 4632 5540 4684
rect 5592 4632 5598 4684
rect 8294 4672 8300 4684
rect 8255 4644 8300 4672
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 9950 4632 9956 4684
rect 10008 4672 10014 4684
rect 10045 4675 10103 4681
rect 10045 4672 10057 4675
rect 10008 4644 10057 4672
rect 10008 4632 10014 4644
rect 10045 4641 10057 4644
rect 10091 4641 10103 4675
rect 10045 4635 10103 4641
rect 10870 4632 10876 4684
rect 10928 4672 10934 4684
rect 11149 4675 11207 4681
rect 11149 4672 11161 4675
rect 10928 4644 11161 4672
rect 10928 4632 10934 4644
rect 11149 4641 11161 4644
rect 11195 4641 11207 4675
rect 11532 4672 11560 4700
rect 13998 4672 14004 4684
rect 11532 4644 14004 4672
rect 11149 4635 11207 4641
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 15657 4675 15715 4681
rect 15657 4641 15669 4675
rect 15703 4672 15715 4675
rect 16206 4672 16212 4684
rect 15703 4644 16212 4672
rect 15703 4641 15715 4644
rect 15657 4635 15715 4641
rect 16206 4632 16212 4644
rect 16264 4632 16270 4684
rect 19518 4632 19524 4684
rect 19576 4672 19582 4684
rect 19628 4672 19656 4703
rect 20530 4700 20536 4712
rect 20588 4700 20594 4752
rect 20990 4700 20996 4752
rect 21048 4740 21054 4752
rect 21361 4743 21419 4749
rect 21361 4740 21373 4743
rect 21048 4712 21373 4740
rect 21048 4700 21054 4712
rect 21361 4709 21373 4712
rect 21407 4740 21419 4743
rect 21910 4740 21916 4752
rect 21407 4712 21916 4740
rect 21407 4709 21419 4712
rect 21361 4703 21419 4709
rect 21910 4700 21916 4712
rect 21968 4700 21974 4752
rect 22388 4740 22416 4768
rect 24857 4743 24915 4749
rect 24857 4740 24869 4743
rect 22388 4712 24869 4740
rect 24857 4709 24869 4712
rect 24903 4740 24915 4743
rect 25130 4740 25136 4752
rect 24903 4712 25136 4740
rect 24903 4709 24915 4712
rect 24857 4703 24915 4709
rect 25130 4700 25136 4712
rect 25188 4700 25194 4752
rect 19576 4644 19656 4672
rect 19576 4632 19582 4644
rect 22002 4632 22008 4684
rect 22060 4672 22066 4684
rect 22738 4681 22744 4684
rect 22465 4675 22523 4681
rect 22465 4672 22477 4675
rect 22060 4644 22477 4672
rect 22060 4632 22066 4644
rect 22465 4641 22477 4644
rect 22511 4641 22523 4675
rect 22732 4672 22744 4681
rect 22699 4644 22744 4672
rect 22465 4635 22523 4641
rect 22732 4635 22744 4644
rect 22738 4632 22744 4635
rect 22796 4632 22802 4684
rect 24946 4672 24952 4684
rect 24907 4644 24952 4672
rect 24946 4632 24952 4644
rect 25004 4632 25010 4684
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 3234 4604 3240 4616
rect 2731 4576 3240 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 3234 4564 3240 4576
rect 3292 4604 3298 4616
rect 3421 4607 3479 4613
rect 3421 4604 3433 4607
rect 3292 4576 3433 4604
rect 3292 4564 3298 4576
rect 3421 4573 3433 4576
rect 3467 4573 3479 4607
rect 5350 4604 5356 4616
rect 5311 4576 5356 4604
rect 3421 4567 3479 4573
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 6638 4604 6644 4616
rect 6196 4576 6644 4604
rect 4801 4539 4859 4545
rect 4801 4505 4813 4539
rect 4847 4536 4859 4539
rect 6196 4536 6224 4576
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4604 6975 4607
rect 8202 4604 8208 4616
rect 6963 4576 8208 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 4847 4508 6224 4536
rect 6273 4539 6331 4545
rect 4847 4505 4859 4508
rect 4801 4499 4859 4505
rect 6273 4505 6285 4539
rect 6319 4536 6331 4539
rect 6932 4536 6960 4567
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8481 4607 8539 4613
rect 8481 4573 8493 4607
rect 8527 4573 8539 4607
rect 8481 4567 8539 4573
rect 7466 4536 7472 4548
rect 6319 4508 6960 4536
rect 7379 4508 7472 4536
rect 6319 4505 6331 4508
rect 6273 4499 6331 4505
rect 7466 4496 7472 4508
rect 7524 4536 7530 4548
rect 7837 4539 7895 4545
rect 7837 4536 7849 4539
rect 7524 4508 7849 4536
rect 7524 4496 7530 4508
rect 7837 4505 7849 4508
rect 7883 4536 7895 4539
rect 8496 4536 8524 4567
rect 14090 4564 14096 4616
rect 14148 4604 14154 4616
rect 14185 4607 14243 4613
rect 14185 4604 14197 4607
rect 14148 4576 14197 4604
rect 14148 4564 14154 4576
rect 14185 4573 14197 4576
rect 14231 4573 14243 4607
rect 14185 4567 14243 4573
rect 15841 4607 15899 4613
rect 15841 4573 15853 4607
rect 15887 4573 15899 4607
rect 17494 4604 17500 4616
rect 17455 4576 17500 4604
rect 15841 4567 15899 4573
rect 7883 4508 8524 4536
rect 10229 4539 10287 4545
rect 7883 4505 7895 4508
rect 7837 4499 7895 4505
rect 10229 4505 10241 4539
rect 10275 4536 10287 4539
rect 10778 4536 10784 4548
rect 10275 4508 10784 4536
rect 10275 4505 10287 4508
rect 10229 4499 10287 4505
rect 10778 4496 10784 4508
rect 10836 4496 10842 4548
rect 10888 4508 11192 4536
rect 3050 4468 3056 4480
rect 3011 4440 3056 4468
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4249 4471 4307 4477
rect 4249 4468 4261 4471
rect 4212 4440 4261 4468
rect 4212 4428 4218 4440
rect 4249 4437 4261 4440
rect 4295 4437 4307 4471
rect 4249 4431 4307 4437
rect 5442 4428 5448 4480
rect 5500 4468 5506 4480
rect 5813 4471 5871 4477
rect 5813 4468 5825 4471
rect 5500 4440 5825 4468
rect 5500 4428 5506 4440
rect 5813 4437 5825 4440
rect 5859 4468 5871 4471
rect 6362 4468 6368 4480
rect 5859 4440 6368 4468
rect 5859 4437 5871 4440
rect 5813 4431 5871 4437
rect 6362 4428 6368 4440
rect 6420 4428 6426 4480
rect 6638 4428 6644 4480
rect 6696 4468 6702 4480
rect 7006 4468 7012 4480
rect 6696 4440 7012 4468
rect 6696 4428 6702 4440
rect 7006 4428 7012 4440
rect 7064 4428 7070 4480
rect 8846 4428 8852 4480
rect 8904 4468 8910 4480
rect 9033 4471 9091 4477
rect 9033 4468 9045 4471
rect 8904 4440 9045 4468
rect 8904 4428 8910 4440
rect 9033 4437 9045 4440
rect 9079 4468 9091 4471
rect 9122 4468 9128 4480
rect 9079 4440 9128 4468
rect 9079 4437 9091 4440
rect 9033 4431 9091 4437
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 9953 4471 10011 4477
rect 9953 4437 9965 4471
rect 9999 4468 10011 4471
rect 10042 4468 10048 4480
rect 9999 4440 10048 4468
rect 9999 4437 10011 4440
rect 9953 4431 10011 4437
rect 10042 4428 10048 4440
rect 10100 4468 10106 4480
rect 10888 4468 10916 4508
rect 11054 4468 11060 4480
rect 10100 4440 10916 4468
rect 11015 4440 11060 4468
rect 10100 4428 10106 4440
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 11164 4468 11192 4508
rect 15654 4496 15660 4548
rect 15712 4536 15718 4548
rect 15856 4536 15884 4567
rect 17494 4564 17500 4576
rect 17552 4564 17558 4616
rect 19702 4604 19708 4616
rect 19663 4576 19708 4604
rect 19702 4564 19708 4576
rect 19760 4604 19766 4616
rect 20622 4604 20628 4616
rect 19760 4576 20628 4604
rect 19760 4564 19766 4576
rect 20622 4564 20628 4576
rect 20680 4564 20686 4616
rect 21545 4607 21603 4613
rect 21545 4573 21557 4607
rect 21591 4604 21603 4607
rect 22278 4604 22284 4616
rect 21591 4576 22284 4604
rect 21591 4573 21603 4576
rect 21545 4567 21603 4573
rect 22278 4564 22284 4576
rect 22336 4564 22342 4616
rect 15712 4508 15884 4536
rect 16853 4539 16911 4545
rect 15712 4496 15718 4508
rect 16853 4505 16865 4539
rect 16899 4536 16911 4539
rect 17678 4536 17684 4548
rect 16899 4508 17684 4536
rect 16899 4505 16911 4508
rect 16853 4499 16911 4505
rect 17678 4496 17684 4508
rect 17736 4496 17742 4548
rect 12526 4468 12532 4480
rect 11164 4440 12532 4468
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 13170 4468 13176 4480
rect 13131 4440 13176 4468
rect 13170 4428 13176 4440
rect 13228 4428 13234 4480
rect 13538 4468 13544 4480
rect 13499 4440 13544 4468
rect 13538 4428 13544 4440
rect 13596 4428 13602 4480
rect 14734 4468 14740 4480
rect 14695 4440 14740 4468
rect 14734 4428 14740 4440
rect 14792 4428 14798 4480
rect 15286 4468 15292 4480
rect 15247 4440 15292 4468
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 18322 4468 18328 4480
rect 18283 4440 18328 4468
rect 18322 4428 18328 4440
rect 18380 4428 18386 4480
rect 18693 4471 18751 4477
rect 18693 4437 18705 4471
rect 18739 4468 18751 4471
rect 18874 4468 18880 4480
rect 18739 4440 18880 4468
rect 18739 4437 18751 4440
rect 18693 4431 18751 4437
rect 18874 4428 18880 4440
rect 18932 4428 18938 4480
rect 23842 4468 23848 4480
rect 23803 4440 23848 4468
rect 23842 4428 23848 4440
rect 23900 4428 23906 4480
rect 25133 4471 25191 4477
rect 25133 4437 25145 4471
rect 25179 4468 25191 4471
rect 27062 4468 27068 4480
rect 25179 4440 27068 4468
rect 25179 4437 25191 4440
rect 25133 4431 25191 4437
rect 27062 4428 27068 4440
rect 27120 4428 27126 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 5169 4267 5227 4273
rect 5169 4233 5181 4267
rect 5215 4264 5227 4267
rect 6546 4264 6552 4276
rect 5215 4236 6552 4264
rect 5215 4233 5227 4236
rect 5169 4227 5227 4233
rect 6546 4224 6552 4236
rect 6604 4224 6610 4276
rect 9953 4267 10011 4273
rect 9953 4233 9965 4267
rect 9999 4264 10011 4267
rect 10226 4264 10232 4276
rect 9999 4236 10232 4264
rect 9999 4233 10011 4236
rect 9953 4227 10011 4233
rect 10226 4224 10232 4236
rect 10284 4264 10290 4276
rect 11054 4264 11060 4276
rect 10284 4236 11060 4264
rect 10284 4224 10290 4236
rect 11054 4224 11060 4236
rect 11112 4224 11118 4276
rect 13081 4267 13139 4273
rect 13081 4233 13093 4267
rect 13127 4264 13139 4267
rect 13906 4264 13912 4276
rect 13127 4236 13912 4264
rect 13127 4233 13139 4236
rect 13081 4227 13139 4233
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 13998 4224 14004 4276
rect 14056 4264 14062 4276
rect 14093 4267 14151 4273
rect 14093 4264 14105 4267
rect 14056 4236 14105 4264
rect 14056 4224 14062 4236
rect 14093 4233 14105 4236
rect 14139 4233 14151 4267
rect 16206 4264 16212 4276
rect 16167 4236 16212 4264
rect 14093 4227 14151 4233
rect 16206 4224 16212 4236
rect 16264 4224 16270 4276
rect 17313 4267 17371 4273
rect 17313 4233 17325 4267
rect 17359 4264 17371 4267
rect 17494 4264 17500 4276
rect 17359 4236 17500 4264
rect 17359 4233 17371 4236
rect 17313 4227 17371 4233
rect 17494 4224 17500 4236
rect 17552 4224 17558 4276
rect 19337 4267 19395 4273
rect 19337 4233 19349 4267
rect 19383 4264 19395 4267
rect 19702 4264 19708 4276
rect 19383 4236 19708 4264
rect 19383 4233 19395 4236
rect 19337 4227 19395 4233
rect 19702 4224 19708 4236
rect 19760 4224 19766 4276
rect 21634 4224 21640 4276
rect 21692 4264 21698 4276
rect 21729 4267 21787 4273
rect 21729 4264 21741 4267
rect 21692 4236 21741 4264
rect 21692 4224 21698 4236
rect 21729 4233 21741 4236
rect 21775 4233 21787 4267
rect 21729 4227 21787 4233
rect 22738 4224 22744 4276
rect 22796 4264 22802 4276
rect 23385 4267 23443 4273
rect 23385 4264 23397 4267
rect 22796 4236 23397 4264
rect 22796 4224 22802 4236
rect 23385 4233 23397 4236
rect 23431 4233 23443 4267
rect 23385 4227 23443 4233
rect 24946 4224 24952 4276
rect 25004 4264 25010 4276
rect 25869 4267 25927 4273
rect 25869 4264 25881 4267
rect 25004 4236 25881 4264
rect 25004 4224 25010 4236
rect 25869 4233 25881 4236
rect 25915 4233 25927 4267
rect 25869 4227 25927 4233
rect 4525 4199 4583 4205
rect 4525 4165 4537 4199
rect 4571 4196 4583 4199
rect 4893 4199 4951 4205
rect 4893 4196 4905 4199
rect 4571 4168 4905 4196
rect 4571 4165 4583 4168
rect 4525 4159 4583 4165
rect 4893 4165 4905 4168
rect 4939 4196 4951 4199
rect 5350 4196 5356 4208
rect 4939 4168 5356 4196
rect 4939 4165 4951 4168
rect 4893 4159 4951 4165
rect 5350 4156 5356 4168
rect 5408 4196 5414 4208
rect 5408 4168 5764 4196
rect 5408 4156 5414 4168
rect 1946 4128 1952 4140
rect 1907 4100 1952 4128
rect 1946 4088 1952 4100
rect 2004 4128 2010 4140
rect 5736 4137 5764 4168
rect 6730 4156 6736 4208
rect 6788 4196 6794 4208
rect 7466 4196 7472 4208
rect 6788 4168 7472 4196
rect 6788 4156 6794 4168
rect 7392 4137 7420 4168
rect 7466 4156 7472 4168
rect 7524 4156 7530 4208
rect 9122 4196 9128 4208
rect 9048 4168 9128 4196
rect 2041 4131 2099 4137
rect 2041 4128 2053 4131
rect 2004 4100 2053 4128
rect 2004 4088 2010 4100
rect 2041 4097 2053 4100
rect 2087 4097 2099 4131
rect 2041 4091 2099 4097
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4097 5779 4131
rect 5721 4091 5779 4097
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 9048 4137 9076 4168
rect 9122 4156 9128 4168
rect 9180 4156 9186 4208
rect 10870 4156 10876 4208
rect 10928 4196 10934 4208
rect 11149 4199 11207 4205
rect 11149 4196 11161 4199
rect 10928 4168 11161 4196
rect 10928 4156 10934 4168
rect 11149 4165 11161 4168
rect 11195 4165 11207 4199
rect 11149 4159 11207 4165
rect 11238 4156 11244 4208
rect 11296 4196 11302 4208
rect 11517 4199 11575 4205
rect 11517 4196 11529 4199
rect 11296 4168 11529 4196
rect 11296 4156 11302 4168
rect 11517 4165 11529 4168
rect 11563 4165 11575 4199
rect 11517 4159 11575 4165
rect 13170 4156 13176 4208
rect 13228 4196 13234 4208
rect 13228 4168 13676 4196
rect 13228 4156 13234 4168
rect 8849 4131 8907 4137
rect 8849 4128 8861 4131
rect 7616 4100 8861 4128
rect 7616 4088 7622 4100
rect 8849 4097 8861 4100
rect 8895 4097 8907 4131
rect 8849 4091 8907 4097
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4097 9091 4131
rect 9858 4128 9864 4140
rect 9771 4100 9864 4128
rect 9033 4091 9091 4097
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4060 5687 4063
rect 5994 4060 6000 4072
rect 5675 4032 6000 4060
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 6362 4020 6368 4072
rect 6420 4060 6426 4072
rect 7285 4063 7343 4069
rect 7285 4060 7297 4063
rect 6420 4032 7297 4060
rect 6420 4020 6426 4032
rect 7285 4029 7297 4032
rect 7331 4060 7343 4063
rect 7926 4060 7932 4072
rect 7331 4032 7932 4060
rect 7331 4029 7343 4032
rect 7285 4023 7343 4029
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 8864 4060 8892 4091
rect 9858 4088 9864 4100
rect 9916 4128 9922 4140
rect 10505 4131 10563 4137
rect 10505 4128 10517 4131
rect 9916 4100 10517 4128
rect 9916 4088 9922 4100
rect 10505 4097 10517 4100
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 13354 4088 13360 4140
rect 13412 4128 13418 4140
rect 13648 4137 13676 4168
rect 13541 4131 13599 4137
rect 13541 4128 13553 4131
rect 13412 4100 13553 4128
rect 13412 4088 13418 4100
rect 13541 4097 13553 4100
rect 13587 4097 13599 4131
rect 13541 4091 13599 4097
rect 13633 4131 13691 4137
rect 13633 4097 13645 4131
rect 13679 4097 13691 4131
rect 14550 4128 14556 4140
rect 14511 4100 14556 4128
rect 13633 4091 13691 4097
rect 14550 4088 14556 4100
rect 14608 4088 14614 4140
rect 14734 4088 14740 4140
rect 14792 4128 14798 4140
rect 15197 4131 15255 4137
rect 15197 4128 15209 4131
rect 14792 4100 15209 4128
rect 14792 4088 14798 4100
rect 15197 4097 15209 4100
rect 15243 4097 15255 4131
rect 16761 4131 16819 4137
rect 16761 4128 16773 4131
rect 15197 4091 15255 4097
rect 16040 4100 16773 4128
rect 9398 4060 9404 4072
rect 8864 4032 9404 4060
rect 9398 4020 9404 4032
rect 9456 4020 9462 4072
rect 10413 4063 10471 4069
rect 10413 4029 10425 4063
rect 10459 4060 10471 4063
rect 10686 4060 10692 4072
rect 10459 4032 10692 4060
rect 10459 4029 10471 4032
rect 10413 4023 10471 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 11422 4060 11428 4072
rect 10796 4032 11428 4060
rect 2308 3995 2366 4001
rect 2308 3961 2320 3995
rect 2354 3992 2366 3995
rect 3234 3992 3240 4004
rect 2354 3964 3240 3992
rect 2354 3961 2366 3964
rect 2308 3955 2366 3961
rect 3234 3952 3240 3964
rect 3292 3952 3298 4004
rect 5537 3995 5595 4001
rect 5537 3961 5549 3995
rect 5583 3992 5595 3995
rect 8757 3995 8815 4001
rect 8757 3992 8769 3995
rect 5583 3964 6868 3992
rect 5583 3961 5595 3964
rect 5537 3955 5595 3961
rect 6840 3936 6868 3964
rect 8220 3964 8769 3992
rect 8220 3936 8248 3964
rect 8757 3961 8769 3964
rect 8803 3961 8815 3995
rect 8757 3955 8815 3961
rect 2866 3884 2872 3936
rect 2924 3924 2930 3936
rect 3421 3927 3479 3933
rect 3421 3924 3433 3927
rect 2924 3896 3433 3924
rect 2924 3884 2930 3896
rect 3421 3893 3433 3896
rect 3467 3924 3479 3927
rect 4062 3924 4068 3936
rect 3467 3896 4068 3924
rect 3467 3893 3479 3896
rect 3421 3887 3479 3893
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 6086 3884 6092 3936
rect 6144 3924 6150 3936
rect 6181 3927 6239 3933
rect 6181 3924 6193 3927
rect 6144 3896 6193 3924
rect 6144 3884 6150 3896
rect 6181 3893 6193 3896
rect 6227 3893 6239 3927
rect 6181 3887 6239 3893
rect 6362 3884 6368 3936
rect 6420 3924 6426 3936
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 6420 3896 6561 3924
rect 6420 3884 6426 3896
rect 6549 3893 6561 3896
rect 6595 3893 6607 3927
rect 6822 3924 6828 3936
rect 6783 3896 6828 3924
rect 6549 3887 6607 3893
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 7190 3924 7196 3936
rect 7151 3896 7196 3924
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 8202 3924 8208 3936
rect 8067 3896 8208 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8386 3924 8392 3936
rect 8347 3896 8392 3924
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 10100 3896 10333 3924
rect 10100 3884 10106 3896
rect 10321 3893 10333 3896
rect 10367 3924 10379 3927
rect 10796 3924 10824 4032
rect 11422 4020 11428 4032
rect 11480 4020 11486 4072
rect 12158 4060 12164 4072
rect 12119 4032 12164 4060
rect 12158 4020 12164 4032
rect 12216 4020 12222 4072
rect 12710 4020 12716 4072
rect 12768 4060 12774 4072
rect 12989 4063 13047 4069
rect 12989 4060 13001 4063
rect 12768 4032 13001 4060
rect 12768 4020 12774 4032
rect 12989 4029 13001 4032
rect 13035 4029 13047 4063
rect 12989 4023 13047 4029
rect 13004 3992 13032 4023
rect 13170 4020 13176 4072
rect 13228 4060 13234 4072
rect 13372 4060 13400 4088
rect 13228 4032 13400 4060
rect 14568 4060 14596 4088
rect 15105 4063 15163 4069
rect 15105 4060 15117 4063
rect 14568 4032 15117 4060
rect 13228 4020 13234 4032
rect 15105 4029 15117 4032
rect 15151 4029 15163 4063
rect 15933 4063 15991 4069
rect 15933 4060 15945 4063
rect 15105 4023 15163 4029
rect 15488 4032 15945 4060
rect 13449 3995 13507 4001
rect 13449 3992 13461 3995
rect 13004 3964 13461 3992
rect 13449 3961 13461 3964
rect 13495 3961 13507 3995
rect 15010 3992 15016 4004
rect 14971 3964 15016 3992
rect 13449 3955 13507 3961
rect 15010 3952 15016 3964
rect 15068 3952 15074 4004
rect 10367 3896 10824 3924
rect 10367 3893 10379 3896
rect 10321 3887 10379 3893
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 14645 3927 14703 3933
rect 14645 3924 14657 3927
rect 12492 3896 14657 3924
rect 12492 3884 12498 3896
rect 14645 3893 14657 3896
rect 14691 3924 14703 3927
rect 15488 3924 15516 4032
rect 15933 4029 15945 4032
rect 15979 4029 15991 4063
rect 15933 4023 15991 4029
rect 15562 3952 15568 4004
rect 15620 3992 15626 4004
rect 16040 4001 16068 4100
rect 16761 4097 16773 4100
rect 16807 4097 16819 4131
rect 16761 4091 16819 4097
rect 17678 4088 17684 4140
rect 17736 4128 17742 4140
rect 17865 4131 17923 4137
rect 17865 4128 17877 4131
rect 17736 4100 17877 4128
rect 17736 4088 17742 4100
rect 17865 4097 17877 4100
rect 17911 4128 17923 4131
rect 18230 4128 18236 4140
rect 17911 4100 18236 4128
rect 17911 4097 17923 4100
rect 17865 4091 17923 4097
rect 18230 4088 18236 4100
rect 18288 4088 18294 4140
rect 18322 4088 18328 4140
rect 18380 4128 18386 4140
rect 18690 4128 18696 4140
rect 18380 4100 18696 4128
rect 18380 4088 18386 4100
rect 18690 4088 18696 4100
rect 18748 4088 18754 4140
rect 18874 4128 18880 4140
rect 18835 4100 18880 4128
rect 18874 4088 18880 4100
rect 18932 4088 18938 4140
rect 19889 4131 19947 4137
rect 19889 4097 19901 4131
rect 19935 4128 19947 4131
rect 21269 4131 21327 4137
rect 21269 4128 21281 4131
rect 19935 4100 21281 4128
rect 19935 4097 19947 4100
rect 19889 4091 19947 4097
rect 21269 4097 21281 4100
rect 21315 4128 21327 4131
rect 21910 4128 21916 4140
rect 21315 4100 21916 4128
rect 21315 4097 21327 4100
rect 21269 4091 21327 4097
rect 21910 4088 21916 4100
rect 21968 4088 21974 4140
rect 22094 4088 22100 4140
rect 22152 4128 22158 4140
rect 23017 4131 23075 4137
rect 23017 4128 23029 4131
rect 22152 4100 23029 4128
rect 22152 4088 22158 4100
rect 23017 4097 23029 4100
rect 23063 4128 23075 4131
rect 23566 4128 23572 4140
rect 23063 4100 23572 4128
rect 23063 4097 23075 4100
rect 23017 4091 23075 4097
rect 23566 4088 23572 4100
rect 23624 4088 23630 4140
rect 24765 4131 24823 4137
rect 24765 4097 24777 4131
rect 24811 4128 24823 4131
rect 25130 4128 25136 4140
rect 24811 4100 25136 4128
rect 24811 4097 24823 4100
rect 24765 4091 24823 4097
rect 25130 4088 25136 4100
rect 25188 4088 25194 4140
rect 16574 4060 16580 4072
rect 16535 4032 16580 4060
rect 16574 4020 16580 4032
rect 16632 4020 16638 4072
rect 18248 4060 18276 4088
rect 18601 4063 18659 4069
rect 18601 4060 18613 4063
rect 18248 4032 18613 4060
rect 18601 4029 18613 4032
rect 18647 4029 18659 4063
rect 18601 4023 18659 4029
rect 20530 4020 20536 4072
rect 20588 4060 20594 4072
rect 21085 4063 21143 4069
rect 21085 4060 21097 4063
rect 20588 4032 21097 4060
rect 20588 4020 20594 4032
rect 21085 4029 21097 4032
rect 21131 4029 21143 4063
rect 22462 4060 22468 4072
rect 22423 4032 22468 4060
rect 21085 4023 21143 4029
rect 22462 4020 22468 4032
rect 22520 4020 22526 4072
rect 23658 4020 23664 4072
rect 23716 4060 23722 4072
rect 23716 4032 23980 4060
rect 23716 4020 23722 4032
rect 16025 3995 16083 4001
rect 16025 3992 16037 3995
rect 15620 3964 16037 3992
rect 15620 3952 15626 3964
rect 16025 3961 16037 3964
rect 16071 3961 16083 3995
rect 16025 3955 16083 3961
rect 16390 3952 16396 4004
rect 16448 3992 16454 4004
rect 16669 3995 16727 4001
rect 16669 3992 16681 3995
rect 16448 3964 16681 3992
rect 16448 3952 16454 3964
rect 16669 3961 16681 3964
rect 16715 3961 16727 3995
rect 16669 3955 16727 3961
rect 20257 3995 20315 4001
rect 20257 3961 20269 3995
rect 20303 3992 20315 3995
rect 22189 3995 22247 4001
rect 20303 3964 21220 3992
rect 20303 3961 20315 3964
rect 20257 3955 20315 3961
rect 21192 3936 21220 3964
rect 22189 3961 22201 3995
rect 22235 3992 22247 3995
rect 22278 3992 22284 4004
rect 22235 3964 22284 3992
rect 22235 3961 22247 3964
rect 22189 3955 22247 3961
rect 22278 3952 22284 3964
rect 22336 3992 22342 4004
rect 23842 3992 23848 4004
rect 22336 3964 23848 3992
rect 22336 3952 22342 3964
rect 23842 3952 23848 3964
rect 23900 3952 23906 4004
rect 23952 3992 23980 4032
rect 24026 4020 24032 4072
rect 24084 4060 24090 4072
rect 24489 4063 24547 4069
rect 24489 4060 24501 4063
rect 24084 4032 24501 4060
rect 24084 4020 24090 4032
rect 24489 4029 24501 4032
rect 24535 4029 24547 4063
rect 24489 4023 24547 4029
rect 23952 3964 24164 3992
rect 15654 3924 15660 3936
rect 14691 3896 15516 3924
rect 15615 3896 15660 3924
rect 14691 3893 14703 3896
rect 14645 3887 14703 3893
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 15930 3924 15936 3936
rect 15891 3896 15936 3924
rect 15930 3884 15936 3896
rect 15988 3884 15994 3936
rect 18230 3924 18236 3936
rect 18191 3896 18236 3924
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 20530 3924 20536 3936
rect 20491 3896 20536 3924
rect 20530 3884 20536 3896
rect 20588 3884 20594 3936
rect 20714 3924 20720 3936
rect 20675 3896 20720 3924
rect 20714 3884 20720 3896
rect 20772 3884 20778 3936
rect 21174 3884 21180 3936
rect 21232 3924 21238 3936
rect 22646 3924 22652 3936
rect 21232 3896 21277 3924
rect 22607 3896 22652 3924
rect 21232 3884 21238 3896
rect 22646 3884 22652 3896
rect 22704 3884 22710 3936
rect 23198 3884 23204 3936
rect 23256 3924 23262 3936
rect 23937 3927 23995 3933
rect 23937 3924 23949 3927
rect 23256 3896 23949 3924
rect 23256 3884 23262 3896
rect 23937 3893 23949 3896
rect 23983 3924 23995 3927
rect 24026 3924 24032 3936
rect 23983 3896 24032 3924
rect 23983 3893 23995 3896
rect 23937 3887 23995 3893
rect 24026 3884 24032 3896
rect 24084 3884 24090 3936
rect 24136 3933 24164 3964
rect 24210 3952 24216 4004
rect 24268 3992 24274 4004
rect 24581 3995 24639 4001
rect 24581 3992 24593 3995
rect 24268 3964 24593 3992
rect 24268 3952 24274 3964
rect 24581 3961 24593 3964
rect 24627 3992 24639 3995
rect 25501 3995 25559 4001
rect 25501 3992 25513 3995
rect 24627 3964 25513 3992
rect 24627 3961 24639 3964
rect 24581 3955 24639 3961
rect 25501 3961 25513 3964
rect 25547 3961 25559 3995
rect 25501 3955 25559 3961
rect 24121 3927 24179 3933
rect 24121 3893 24133 3927
rect 24167 3893 24179 3927
rect 25130 3924 25136 3936
rect 25091 3896 25136 3924
rect 24121 3887 24179 3893
rect 25130 3884 25136 3896
rect 25188 3884 25194 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 2038 3680 2044 3732
rect 2096 3720 2102 3732
rect 2501 3723 2559 3729
rect 2501 3720 2513 3723
rect 2096 3692 2513 3720
rect 2096 3680 2102 3692
rect 2501 3689 2513 3692
rect 2547 3689 2559 3723
rect 2501 3683 2559 3689
rect 3145 3723 3203 3729
rect 3145 3689 3157 3723
rect 3191 3720 3203 3723
rect 3234 3720 3240 3732
rect 3191 3692 3240 3720
rect 3191 3689 3203 3692
rect 3145 3683 3203 3689
rect 3234 3680 3240 3692
rect 3292 3720 3298 3732
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 3292 3692 3433 3720
rect 3292 3680 3298 3692
rect 3421 3689 3433 3692
rect 3467 3689 3479 3723
rect 3421 3683 3479 3689
rect 5258 3680 5264 3732
rect 5316 3720 5322 3732
rect 5445 3723 5503 3729
rect 5445 3720 5457 3723
rect 5316 3692 5457 3720
rect 5316 3680 5322 3692
rect 5445 3689 5457 3692
rect 5491 3689 5503 3723
rect 5445 3683 5503 3689
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 6549 3723 6607 3729
rect 6549 3720 6561 3723
rect 5592 3692 6561 3720
rect 5592 3680 5598 3692
rect 6549 3689 6561 3692
rect 6595 3689 6607 3723
rect 8018 3720 8024 3732
rect 7979 3692 8024 3720
rect 6549 3683 6607 3689
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 9493 3723 9551 3729
rect 9493 3689 9505 3723
rect 9539 3720 9551 3723
rect 10042 3720 10048 3732
rect 9539 3692 10048 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 10686 3720 10692 3732
rect 10647 3692 10692 3720
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 12158 3720 12164 3732
rect 12119 3692 12164 3720
rect 12158 3680 12164 3692
rect 12216 3680 12222 3732
rect 12618 3680 12624 3732
rect 12676 3720 12682 3732
rect 12713 3723 12771 3729
rect 12713 3720 12725 3723
rect 12676 3692 12725 3720
rect 12676 3680 12682 3692
rect 12713 3689 12725 3692
rect 12759 3689 12771 3723
rect 13262 3720 13268 3732
rect 13223 3692 13268 3720
rect 12713 3683 12771 3689
rect 13262 3680 13268 3692
rect 13320 3680 13326 3732
rect 14090 3680 14096 3732
rect 14148 3720 14154 3732
rect 14277 3723 14335 3729
rect 14277 3720 14289 3723
rect 14148 3692 14289 3720
rect 14148 3680 14154 3692
rect 14277 3689 14289 3692
rect 14323 3689 14335 3723
rect 14277 3683 14335 3689
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 14792 3692 15025 3720
rect 14792 3680 14798 3692
rect 15013 3689 15025 3692
rect 15059 3689 15071 3723
rect 15013 3683 15071 3689
rect 15289 3723 15347 3729
rect 15289 3689 15301 3723
rect 15335 3720 15347 3723
rect 15378 3720 15384 3732
rect 15335 3692 15384 3720
rect 15335 3689 15347 3692
rect 15289 3683 15347 3689
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 15749 3723 15807 3729
rect 15749 3689 15761 3723
rect 15795 3720 15807 3723
rect 15930 3720 15936 3732
rect 15795 3692 15936 3720
rect 15795 3689 15807 3692
rect 15749 3683 15807 3689
rect 15930 3680 15936 3692
rect 15988 3680 15994 3732
rect 16206 3680 16212 3732
rect 16264 3720 16270 3732
rect 16669 3723 16727 3729
rect 16669 3720 16681 3723
rect 16264 3692 16681 3720
rect 16264 3680 16270 3692
rect 16669 3689 16681 3692
rect 16715 3689 16727 3723
rect 16669 3683 16727 3689
rect 17037 3723 17095 3729
rect 17037 3689 17049 3723
rect 17083 3720 17095 3723
rect 17218 3720 17224 3732
rect 17083 3692 17224 3720
rect 17083 3689 17095 3692
rect 17037 3683 17095 3689
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 17402 3720 17408 3732
rect 17363 3692 17408 3720
rect 17402 3680 17408 3692
rect 17460 3680 17466 3732
rect 18046 3720 18052 3732
rect 18007 3692 18052 3720
rect 18046 3680 18052 3692
rect 18104 3680 18110 3732
rect 18230 3680 18236 3732
rect 18288 3720 18294 3732
rect 18509 3723 18567 3729
rect 18509 3720 18521 3723
rect 18288 3692 18521 3720
rect 18288 3680 18294 3692
rect 18509 3689 18521 3692
rect 18555 3689 18567 3723
rect 18509 3683 18567 3689
rect 18690 3680 18696 3732
rect 18748 3720 18754 3732
rect 18874 3720 18880 3732
rect 18748 3692 18880 3720
rect 18748 3680 18754 3692
rect 18874 3680 18880 3692
rect 18932 3720 18938 3732
rect 19061 3723 19119 3729
rect 19061 3720 19073 3723
rect 18932 3692 19073 3720
rect 18932 3680 18938 3692
rect 19061 3689 19073 3692
rect 19107 3720 19119 3723
rect 19426 3720 19432 3732
rect 19107 3692 19432 3720
rect 19107 3689 19119 3692
rect 19061 3683 19119 3689
rect 19426 3680 19432 3692
rect 19484 3680 19490 3732
rect 19518 3680 19524 3732
rect 19576 3720 19582 3732
rect 19576 3692 19621 3720
rect 19576 3680 19582 3692
rect 20714 3680 20720 3732
rect 20772 3720 20778 3732
rect 21358 3720 21364 3732
rect 20772 3692 21364 3720
rect 20772 3680 20778 3692
rect 21358 3680 21364 3692
rect 21416 3680 21422 3732
rect 21910 3720 21916 3732
rect 21871 3692 21916 3720
rect 21910 3680 21916 3692
rect 21968 3680 21974 3732
rect 22186 3680 22192 3732
rect 22244 3720 22250 3732
rect 22281 3723 22339 3729
rect 22281 3720 22293 3723
rect 22244 3692 22293 3720
rect 22244 3680 22250 3692
rect 22281 3689 22293 3692
rect 22327 3689 22339 3723
rect 22281 3683 22339 3689
rect 2406 3652 2412 3664
rect 2319 3624 2412 3652
rect 2406 3612 2412 3624
rect 2464 3652 2470 3664
rect 3326 3652 3332 3664
rect 2464 3624 3332 3652
rect 2464 3612 2470 3624
rect 3326 3612 3332 3624
rect 3384 3612 3390 3664
rect 4062 3612 4068 3664
rect 4120 3652 4126 3664
rect 4310 3655 4368 3661
rect 4310 3652 4322 3655
rect 4120 3624 4322 3652
rect 4120 3612 4126 3624
rect 4310 3621 4322 3624
rect 4356 3621 4368 3655
rect 9950 3652 9956 3664
rect 4310 3615 4368 3621
rect 9692 3624 9956 3652
rect 4154 3584 4160 3596
rect 4080 3556 4160 3584
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3516 2743 3519
rect 2866 3516 2872 3528
rect 2731 3488 2872 3516
rect 2731 3485 2743 3488
rect 2685 3479 2743 3485
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 3878 3476 3884 3528
rect 3936 3516 3942 3528
rect 4080 3525 4108 3556
rect 4154 3544 4160 3556
rect 4212 3544 4218 3596
rect 6546 3544 6552 3596
rect 6604 3584 6610 3596
rect 9692 3593 9720 3624
rect 9950 3612 9956 3624
rect 10008 3652 10014 3664
rect 11054 3661 11060 3664
rect 10229 3655 10287 3661
rect 10229 3652 10241 3655
rect 10008 3624 10241 3652
rect 10008 3612 10014 3624
rect 10229 3621 10241 3624
rect 10275 3621 10287 3655
rect 11048 3652 11060 3661
rect 10967 3624 11060 3652
rect 10229 3615 10287 3621
rect 11048 3615 11060 3624
rect 11112 3652 11118 3664
rect 11974 3652 11980 3664
rect 11112 3624 11980 3652
rect 11054 3612 11060 3615
rect 11112 3612 11118 3624
rect 11974 3612 11980 3624
rect 12032 3612 12038 3664
rect 12250 3612 12256 3664
rect 12308 3652 12314 3664
rect 12308 3624 16896 3652
rect 12308 3612 12314 3624
rect 6917 3587 6975 3593
rect 6917 3584 6929 3587
rect 6604 3556 6929 3584
rect 6604 3544 6610 3556
rect 6917 3553 6929 3556
rect 6963 3584 6975 3587
rect 9677 3587 9735 3593
rect 6963 3556 7512 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 4065 3519 4123 3525
rect 4065 3516 4077 3519
rect 3936 3488 4077 3516
rect 3936 3476 3942 3488
rect 4065 3485 4077 3488
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 6730 3476 6736 3528
rect 6788 3516 6794 3528
rect 7009 3519 7067 3525
rect 7009 3516 7021 3519
rect 6788 3488 7021 3516
rect 6788 3476 6794 3488
rect 7009 3485 7021 3488
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 7101 3519 7159 3525
rect 7101 3485 7113 3519
rect 7147 3485 7159 3519
rect 7101 3479 7159 3485
rect 2041 3451 2099 3457
rect 2041 3417 2053 3451
rect 2087 3448 2099 3451
rect 2130 3448 2136 3460
rect 2087 3420 2136 3448
rect 2087 3417 2099 3420
rect 2041 3411 2099 3417
rect 2130 3408 2136 3420
rect 2188 3408 2194 3460
rect 7116 3448 7144 3479
rect 7374 3448 7380 3460
rect 6380 3420 7380 3448
rect 1673 3383 1731 3389
rect 1673 3349 1685 3383
rect 1719 3380 1731 3383
rect 1854 3380 1860 3392
rect 1719 3352 1860 3380
rect 1719 3349 1731 3352
rect 1673 3343 1731 3349
rect 1854 3340 1860 3352
rect 1912 3340 1918 3392
rect 3881 3383 3939 3389
rect 3881 3349 3893 3383
rect 3927 3380 3939 3383
rect 4338 3380 4344 3392
rect 3927 3352 4344 3380
rect 3927 3349 3939 3352
rect 3881 3343 3939 3349
rect 4338 3340 4344 3352
rect 4396 3340 4402 3392
rect 5534 3340 5540 3392
rect 5592 3380 5598 3392
rect 6380 3389 6408 3420
rect 7374 3408 7380 3420
rect 7432 3408 7438 3460
rect 7484 3448 7512 3556
rect 9677 3553 9689 3587
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 10781 3587 10839 3593
rect 10781 3553 10793 3587
rect 10827 3584 10839 3587
rect 10870 3584 10876 3596
rect 10827 3556 10876 3584
rect 10827 3553 10839 3556
rect 10781 3547 10839 3553
rect 10870 3544 10876 3556
rect 10928 3544 10934 3596
rect 13170 3584 13176 3596
rect 13131 3556 13176 3584
rect 13170 3544 13176 3556
rect 13228 3544 13234 3596
rect 13354 3544 13360 3596
rect 13412 3584 13418 3596
rect 13633 3587 13691 3593
rect 13633 3584 13645 3587
rect 13412 3556 13645 3584
rect 13412 3544 13418 3556
rect 13633 3553 13645 3556
rect 13679 3553 13691 3587
rect 13633 3547 13691 3553
rect 15286 3544 15292 3596
rect 15344 3584 15350 3596
rect 15657 3587 15715 3593
rect 15657 3584 15669 3587
rect 15344 3556 15669 3584
rect 15344 3544 15350 3556
rect 15657 3553 15669 3556
rect 15703 3584 15715 3587
rect 16206 3584 16212 3596
rect 15703 3556 16212 3584
rect 15703 3553 15715 3556
rect 15657 3547 15715 3553
rect 16206 3544 16212 3556
rect 16264 3544 16270 3596
rect 16390 3584 16396 3596
rect 16351 3556 16396 3584
rect 16390 3544 16396 3556
rect 16448 3544 16454 3596
rect 16868 3593 16896 3624
rect 17494 3612 17500 3664
rect 17552 3652 17558 3664
rect 18417 3655 18475 3661
rect 18417 3652 18429 3655
rect 17552 3624 18429 3652
rect 17552 3612 17558 3624
rect 18417 3621 18429 3624
rect 18463 3652 18475 3655
rect 18598 3652 18604 3664
rect 18463 3624 18604 3652
rect 18463 3621 18475 3624
rect 18417 3615 18475 3621
rect 18598 3612 18604 3624
rect 18656 3612 18662 3664
rect 20898 3612 20904 3664
rect 20956 3652 20962 3664
rect 21269 3655 21327 3661
rect 21269 3652 21281 3655
rect 20956 3624 21281 3652
rect 20956 3612 20962 3624
rect 21269 3621 21281 3624
rect 21315 3621 21327 3655
rect 21269 3615 21327 3621
rect 16853 3587 16911 3593
rect 16853 3553 16865 3587
rect 16899 3553 16911 3587
rect 16853 3547 16911 3553
rect 19705 3587 19763 3593
rect 19705 3553 19717 3587
rect 19751 3584 19763 3587
rect 20070 3584 20076 3596
rect 19751 3556 20076 3584
rect 19751 3553 19763 3556
rect 19705 3547 19763 3553
rect 20070 3544 20076 3556
rect 20128 3584 20134 3596
rect 20257 3587 20315 3593
rect 20257 3584 20269 3587
rect 20128 3556 20269 3584
rect 20128 3544 20134 3556
rect 20257 3553 20269 3556
rect 20303 3553 20315 3587
rect 20257 3547 20315 3553
rect 20717 3587 20775 3593
rect 20717 3553 20729 3587
rect 20763 3584 20775 3587
rect 20990 3584 20996 3596
rect 20763 3556 20996 3584
rect 20763 3553 20775 3556
rect 20717 3547 20775 3553
rect 20990 3544 20996 3556
rect 21048 3544 21054 3596
rect 22296 3584 22324 3683
rect 22462 3680 22468 3732
rect 22520 3720 22526 3732
rect 23017 3723 23075 3729
rect 23017 3720 23029 3723
rect 22520 3692 23029 3720
rect 22520 3680 22526 3692
rect 23017 3689 23029 3692
rect 23063 3689 23075 3723
rect 23017 3683 23075 3689
rect 23842 3661 23848 3664
rect 23836 3652 23848 3661
rect 23803 3624 23848 3652
rect 23836 3615 23848 3624
rect 23842 3612 23848 3615
rect 23900 3612 23906 3664
rect 22465 3587 22523 3593
rect 22465 3584 22477 3587
rect 22296 3556 22477 3584
rect 22465 3553 22477 3556
rect 22511 3553 22523 3587
rect 23566 3584 23572 3596
rect 23527 3556 23572 3584
rect 22465 3547 22523 3553
rect 23566 3544 23572 3556
rect 23624 3544 23630 3596
rect 7650 3516 7656 3528
rect 7611 3488 7656 3516
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 8570 3516 8576 3528
rect 8531 3488 8576 3516
rect 8570 3476 8576 3488
rect 8628 3476 8634 3528
rect 13722 3516 13728 3528
rect 13683 3488 13728 3516
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 15838 3516 15844 3528
rect 13872 3488 13917 3516
rect 15799 3488 15844 3516
rect 13872 3476 13878 3488
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 18506 3476 18512 3528
rect 18564 3516 18570 3528
rect 18601 3519 18659 3525
rect 18601 3516 18613 3519
rect 18564 3488 18613 3516
rect 18564 3476 18570 3488
rect 18601 3485 18613 3488
rect 18647 3485 18659 3519
rect 21450 3516 21456 3528
rect 21411 3488 21456 3516
rect 18601 3479 18659 3485
rect 21450 3476 21456 3488
rect 21508 3476 21514 3528
rect 15010 3448 15016 3460
rect 7484 3420 9996 3448
rect 5997 3383 6055 3389
rect 5997 3380 6009 3383
rect 5592 3352 6009 3380
rect 5592 3340 5598 3352
rect 5997 3349 6009 3352
rect 6043 3380 6055 3383
rect 6365 3383 6423 3389
rect 6365 3380 6377 3383
rect 6043 3352 6377 3380
rect 6043 3349 6055 3352
rect 5997 3343 6055 3349
rect 6365 3349 6377 3352
rect 6411 3349 6423 3383
rect 6365 3343 6423 3349
rect 8202 3340 8208 3392
rect 8260 3380 8266 3392
rect 8389 3383 8447 3389
rect 8389 3380 8401 3383
rect 8260 3352 8401 3380
rect 8260 3340 8266 3352
rect 8389 3349 8401 3352
rect 8435 3349 8447 3383
rect 8389 3343 8447 3349
rect 9125 3383 9183 3389
rect 9125 3349 9137 3383
rect 9171 3380 9183 3383
rect 9582 3380 9588 3392
rect 9171 3352 9588 3380
rect 9171 3349 9183 3352
rect 9125 3343 9183 3349
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 9858 3380 9864 3392
rect 9819 3352 9864 3380
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 9968 3380 9996 3420
rect 14660 3420 15016 3448
rect 11146 3380 11152 3392
rect 9968 3352 11152 3380
rect 11146 3340 11152 3352
rect 11204 3340 11210 3392
rect 14550 3340 14556 3392
rect 14608 3380 14614 3392
rect 14660 3389 14688 3420
rect 15010 3408 15016 3420
rect 15068 3408 15074 3460
rect 17957 3451 18015 3457
rect 17957 3417 17969 3451
rect 18003 3448 18015 3451
rect 18138 3448 18144 3460
rect 18003 3420 18144 3448
rect 18003 3417 18015 3420
rect 17957 3411 18015 3417
rect 18138 3408 18144 3420
rect 18196 3408 18202 3460
rect 20901 3451 20959 3457
rect 20901 3417 20913 3451
rect 20947 3448 20959 3451
rect 21266 3448 21272 3460
rect 20947 3420 21272 3448
rect 20947 3417 20959 3420
rect 20901 3411 20959 3417
rect 21266 3408 21272 3420
rect 21324 3408 21330 3460
rect 14645 3383 14703 3389
rect 14645 3380 14657 3383
rect 14608 3352 14657 3380
rect 14608 3340 14614 3352
rect 14645 3349 14657 3352
rect 14691 3349 14703 3383
rect 19886 3380 19892 3392
rect 19847 3352 19892 3380
rect 14645 3343 14703 3349
rect 19886 3340 19892 3352
rect 19944 3340 19950 3392
rect 22646 3380 22652 3392
rect 22607 3352 22652 3380
rect 22646 3340 22652 3352
rect 22704 3340 22710 3392
rect 23477 3383 23535 3389
rect 23477 3349 23489 3383
rect 23523 3380 23535 3383
rect 24762 3380 24768 3392
rect 23523 3352 24768 3380
rect 23523 3349 23535 3352
rect 23477 3343 23535 3349
rect 24762 3340 24768 3352
rect 24820 3380 24826 3392
rect 24949 3383 25007 3389
rect 24949 3380 24961 3383
rect 24820 3352 24961 3380
rect 24820 3340 24826 3352
rect 24949 3349 24961 3352
rect 24995 3349 25007 3383
rect 24949 3343 25007 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1946 3176 1952 3188
rect 1596 3148 1952 3176
rect 1596 3049 1624 3148
rect 1946 3136 1952 3148
rect 2004 3136 2010 3188
rect 2961 3179 3019 3185
rect 2961 3145 2973 3179
rect 3007 3176 3019 3179
rect 3234 3176 3240 3188
rect 3007 3148 3240 3176
rect 3007 3145 3019 3148
rect 2961 3139 3019 3145
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 4614 3136 4620 3188
rect 4672 3176 4678 3188
rect 6181 3179 6239 3185
rect 6181 3176 6193 3179
rect 4672 3148 6193 3176
rect 4672 3136 4678 3148
rect 6181 3145 6193 3148
rect 6227 3145 6239 3179
rect 6822 3176 6828 3188
rect 6783 3148 6828 3176
rect 6181 3139 6239 3145
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3040 1639 3043
rect 1627 3012 1716 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 1688 2984 1716 3012
rect 1670 2932 1676 2984
rect 1728 2932 1734 2984
rect 1854 2981 1860 2984
rect 1848 2972 1860 2981
rect 1815 2944 1860 2972
rect 1848 2935 1860 2944
rect 1854 2932 1860 2935
rect 1912 2932 1918 2984
rect 4249 2975 4307 2981
rect 4249 2941 4261 2975
rect 4295 2941 4307 2975
rect 4249 2935 4307 2941
rect 1688 2904 1716 2932
rect 3697 2907 3755 2913
rect 3697 2904 3709 2907
rect 1688 2876 3709 2904
rect 3697 2873 3709 2876
rect 3743 2904 3755 2907
rect 3878 2904 3884 2916
rect 3743 2876 3884 2904
rect 3743 2873 3755 2876
rect 3697 2867 3755 2873
rect 3878 2864 3884 2876
rect 3936 2904 3942 2916
rect 4065 2907 4123 2913
rect 4065 2904 4077 2907
rect 3936 2876 4077 2904
rect 3936 2864 3942 2876
rect 4065 2873 4077 2876
rect 4111 2904 4123 2907
rect 4264 2904 4292 2935
rect 4338 2932 4344 2984
rect 4396 2972 4402 2984
rect 4505 2975 4563 2981
rect 4505 2972 4517 2975
rect 4396 2944 4517 2972
rect 4396 2932 4402 2944
rect 4505 2941 4517 2944
rect 4551 2972 4563 2975
rect 5442 2972 5448 2984
rect 4551 2944 5448 2972
rect 4551 2941 4563 2944
rect 4505 2935 4563 2941
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 6196 2972 6224 3139
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7926 3176 7932 3188
rect 7887 3148 7932 3176
rect 7926 3136 7932 3148
rect 7984 3136 7990 3188
rect 8478 3136 8484 3188
rect 8536 3176 8542 3188
rect 8573 3179 8631 3185
rect 8573 3176 8585 3179
rect 8536 3148 8585 3176
rect 8536 3136 8542 3148
rect 8573 3145 8585 3148
rect 8619 3176 8631 3179
rect 10137 3179 10195 3185
rect 8619 3148 9904 3176
rect 8619 3145 8631 3148
rect 8573 3139 8631 3145
rect 7374 3040 7380 3052
rect 7335 3012 7380 3040
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3040 8355 3043
rect 9876 3040 9904 3148
rect 10137 3145 10149 3179
rect 10183 3176 10195 3179
rect 10226 3176 10232 3188
rect 10183 3148 10232 3176
rect 10183 3145 10195 3148
rect 10137 3139 10195 3145
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 10870 3176 10876 3188
rect 10831 3148 10876 3176
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 11790 3176 11796 3188
rect 11751 3148 11796 3176
rect 11790 3136 11796 3148
rect 11848 3176 11854 3188
rect 12894 3176 12900 3188
rect 11848 3148 12900 3176
rect 11848 3136 11854 3148
rect 12894 3136 12900 3148
rect 12952 3136 12958 3188
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 14185 3179 14243 3185
rect 14185 3176 14197 3179
rect 13872 3148 14197 3176
rect 13872 3136 13878 3148
rect 14185 3145 14197 3148
rect 14231 3145 14243 3179
rect 14185 3139 14243 3145
rect 15838 3136 15844 3188
rect 15896 3176 15902 3188
rect 16117 3179 16175 3185
rect 16117 3176 16129 3179
rect 15896 3148 16129 3176
rect 15896 3136 15902 3148
rect 16117 3145 16129 3148
rect 16163 3176 16175 3179
rect 17037 3179 17095 3185
rect 17037 3176 17049 3179
rect 16163 3148 17049 3176
rect 16163 3145 16175 3148
rect 16117 3139 16175 3145
rect 17037 3145 17049 3148
rect 17083 3145 17095 3179
rect 17494 3176 17500 3188
rect 17455 3148 17500 3176
rect 17037 3139 17095 3145
rect 17494 3136 17500 3148
rect 17552 3136 17558 3188
rect 17770 3176 17776 3188
rect 17731 3148 17776 3176
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 19426 3176 19432 3188
rect 19387 3148 19432 3176
rect 19426 3136 19432 3148
rect 19484 3136 19490 3188
rect 20073 3179 20131 3185
rect 20073 3145 20085 3179
rect 20119 3176 20131 3179
rect 20898 3176 20904 3188
rect 20119 3148 20904 3176
rect 20119 3145 20131 3148
rect 20073 3139 20131 3145
rect 20898 3136 20904 3148
rect 20956 3136 20962 3188
rect 21450 3136 21456 3188
rect 21508 3176 21514 3188
rect 22465 3179 22523 3185
rect 22465 3176 22477 3179
rect 21508 3148 22477 3176
rect 21508 3136 21514 3148
rect 22465 3145 22477 3148
rect 22511 3176 22523 3179
rect 22554 3176 22560 3188
rect 22511 3148 22560 3176
rect 22511 3145 22523 3148
rect 22465 3139 22523 3145
rect 22554 3136 22560 3148
rect 22612 3136 22618 3188
rect 23477 3179 23535 3185
rect 23477 3145 23489 3179
rect 23523 3176 23535 3179
rect 23566 3176 23572 3188
rect 23523 3148 23572 3176
rect 23523 3145 23535 3148
rect 23477 3139 23535 3145
rect 23566 3136 23572 3148
rect 23624 3176 23630 3188
rect 23937 3179 23995 3185
rect 23937 3176 23949 3179
rect 23624 3148 23949 3176
rect 23624 3136 23630 3148
rect 23937 3145 23949 3148
rect 23983 3145 23995 3179
rect 23937 3139 23995 3145
rect 9950 3068 9956 3120
rect 10008 3108 10014 3120
rect 12161 3111 12219 3117
rect 12161 3108 12173 3111
rect 10008 3080 12173 3108
rect 10008 3068 10014 3080
rect 12161 3077 12173 3080
rect 12207 3077 12219 3111
rect 12161 3071 12219 3077
rect 10870 3040 10876 3052
rect 8343 3012 8892 3040
rect 9876 3012 10876 3040
rect 8343 3009 8355 3012
rect 8297 3003 8355 3009
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 6196 2944 7297 2972
rect 7285 2941 7297 2944
rect 7331 2972 7343 2975
rect 7466 2972 7472 2984
rect 7331 2944 7472 2972
rect 7331 2941 7343 2944
rect 7285 2935 7343 2941
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 8478 2932 8484 2984
rect 8536 2972 8542 2984
rect 8757 2975 8815 2981
rect 8757 2972 8769 2975
rect 8536 2944 8769 2972
rect 8536 2932 8542 2944
rect 8757 2941 8769 2944
rect 8803 2941 8815 2975
rect 8864 2972 8892 3012
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 12176 3040 12204 3071
rect 12434 3068 12440 3120
rect 12492 3108 12498 3120
rect 12492 3080 12537 3108
rect 12492 3068 12498 3080
rect 13354 3068 13360 3120
rect 13412 3108 13418 3120
rect 13909 3111 13967 3117
rect 13909 3108 13921 3111
rect 13412 3080 13921 3108
rect 13412 3068 13418 3080
rect 13909 3077 13921 3080
rect 13955 3077 13967 3111
rect 13909 3071 13967 3077
rect 16206 3068 16212 3120
rect 16264 3108 16270 3120
rect 16669 3111 16727 3117
rect 16669 3108 16681 3111
rect 16264 3080 16681 3108
rect 16264 3068 16270 3080
rect 16669 3077 16681 3080
rect 16715 3077 16727 3111
rect 16669 3071 16727 3077
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12176 3012 13001 3040
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 17788 3040 17816 3136
rect 21910 3108 21916 3120
rect 21871 3080 21916 3108
rect 21910 3068 21916 3080
rect 21968 3068 21974 3120
rect 23109 3111 23167 3117
rect 23109 3077 23121 3111
rect 23155 3108 23167 3111
rect 23842 3108 23848 3120
rect 23155 3080 23848 3108
rect 23155 3077 23167 3080
rect 23109 3071 23167 3077
rect 23842 3068 23848 3080
rect 23900 3068 23906 3120
rect 18046 3040 18052 3052
rect 17788 3012 18052 3040
rect 12989 3003 13047 3009
rect 18046 3000 18052 3012
rect 18104 3000 18110 3052
rect 23952 3040 23980 3139
rect 24026 3136 24032 3188
rect 24084 3176 24090 3188
rect 25130 3176 25136 3188
rect 24084 3148 25136 3176
rect 24084 3136 24090 3148
rect 25130 3136 25136 3148
rect 25188 3176 25194 3188
rect 25501 3179 25559 3185
rect 25501 3176 25513 3179
rect 25188 3148 25513 3176
rect 25188 3136 25194 3148
rect 25501 3145 25513 3148
rect 25547 3145 25559 3179
rect 26050 3176 26056 3188
rect 26011 3148 26056 3176
rect 25501 3139 25559 3145
rect 26050 3136 26056 3148
rect 26108 3136 26114 3188
rect 24121 3043 24179 3049
rect 24121 3040 24133 3043
rect 23952 3012 24133 3040
rect 24121 3009 24133 3012
rect 24167 3009 24179 3043
rect 24121 3003 24179 3009
rect 9030 2981 9036 2984
rect 9024 2972 9036 2981
rect 8864 2944 9036 2972
rect 8757 2935 8815 2941
rect 9024 2935 9036 2944
rect 9030 2932 9036 2935
rect 9088 2932 9094 2984
rect 9306 2932 9312 2984
rect 9364 2972 9370 2984
rect 9582 2972 9588 2984
rect 9364 2944 9588 2972
rect 9364 2932 9370 2944
rect 9582 2932 9588 2944
rect 9640 2932 9646 2984
rect 11241 2975 11299 2981
rect 11241 2941 11253 2975
rect 11287 2972 11299 2975
rect 11330 2972 11336 2984
rect 11287 2944 11336 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 11330 2932 11336 2944
rect 11388 2932 11394 2984
rect 12894 2972 12900 2984
rect 12855 2944 12900 2972
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 14568 2944 14749 2972
rect 4111 2876 4292 2904
rect 4356 2876 5764 2904
rect 4111 2873 4123 2876
rect 4065 2867 4123 2873
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 4356 2836 4384 2876
rect 5626 2836 5632 2848
rect 2832 2808 4384 2836
rect 5587 2808 5632 2836
rect 2832 2796 2838 2808
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 5736 2836 5764 2876
rect 6086 2864 6092 2916
rect 6144 2904 6150 2916
rect 6454 2904 6460 2916
rect 6144 2876 6460 2904
rect 6144 2864 6150 2876
rect 6454 2864 6460 2876
rect 6512 2864 6518 2916
rect 6546 2864 6552 2916
rect 6604 2904 6610 2916
rect 6604 2876 6649 2904
rect 6604 2864 6610 2876
rect 12618 2864 12624 2916
rect 12676 2904 12682 2916
rect 12805 2907 12863 2913
rect 12805 2904 12817 2907
rect 12676 2876 12817 2904
rect 12676 2864 12682 2876
rect 12805 2873 12817 2876
rect 12851 2873 12863 2907
rect 12805 2867 12863 2873
rect 7193 2839 7251 2845
rect 7193 2836 7205 2839
rect 5736 2808 7205 2836
rect 7193 2805 7205 2808
rect 7239 2836 7251 2839
rect 7926 2836 7932 2848
rect 7239 2808 7932 2836
rect 7239 2805 7251 2808
rect 7193 2799 7251 2805
rect 7926 2796 7932 2808
rect 7984 2796 7990 2848
rect 11422 2836 11428 2848
rect 11383 2808 11428 2836
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 11514 2796 11520 2848
rect 11572 2836 11578 2848
rect 13449 2839 13507 2845
rect 13449 2836 13461 2839
rect 11572 2808 13461 2836
rect 11572 2796 11578 2808
rect 13449 2805 13461 2808
rect 13495 2836 13507 2839
rect 13722 2836 13728 2848
rect 13495 2808 13728 2836
rect 13495 2805 13507 2808
rect 13449 2799 13507 2805
rect 13722 2796 13728 2808
rect 13780 2796 13786 2848
rect 14458 2796 14464 2848
rect 14516 2836 14522 2848
rect 14568 2845 14596 2944
rect 14737 2941 14749 2944
rect 14783 2941 14795 2975
rect 14737 2935 14795 2941
rect 18138 2932 18144 2984
rect 18196 2972 18202 2984
rect 18305 2975 18363 2981
rect 18305 2972 18317 2975
rect 18196 2944 18317 2972
rect 18196 2932 18202 2944
rect 18305 2941 18317 2944
rect 18351 2941 18363 2975
rect 18305 2935 18363 2941
rect 20533 2975 20591 2981
rect 20533 2941 20545 2975
rect 20579 2941 20591 2975
rect 20533 2935 20591 2941
rect 24388 2975 24446 2981
rect 24388 2941 24400 2975
rect 24434 2972 24446 2975
rect 24762 2972 24768 2984
rect 24434 2944 24768 2972
rect 24434 2941 24446 2944
rect 24388 2935 24446 2941
rect 14826 2864 14832 2916
rect 14884 2904 14890 2916
rect 15010 2913 15016 2916
rect 14982 2907 15016 2913
rect 14982 2904 14994 2907
rect 14884 2876 14994 2904
rect 14884 2864 14890 2876
rect 14982 2873 14994 2876
rect 14982 2867 15016 2873
rect 15010 2864 15016 2867
rect 15068 2864 15074 2916
rect 18046 2864 18052 2916
rect 18104 2904 18110 2916
rect 20548 2904 20576 2935
rect 24762 2932 24768 2944
rect 24820 2932 24826 2984
rect 18104 2876 20576 2904
rect 18104 2864 18110 2876
rect 14553 2839 14611 2845
rect 14553 2836 14565 2839
rect 14516 2808 14565 2836
rect 14516 2796 14522 2808
rect 14553 2805 14565 2808
rect 14599 2805 14611 2839
rect 14553 2799 14611 2805
rect 20441 2839 20499 2845
rect 20441 2805 20453 2839
rect 20487 2836 20499 2839
rect 20548 2836 20576 2876
rect 20714 2864 20720 2916
rect 20772 2913 20778 2916
rect 20772 2907 20836 2913
rect 20772 2873 20790 2907
rect 20824 2873 20836 2907
rect 20772 2867 20836 2873
rect 20772 2864 20778 2867
rect 20898 2836 20904 2848
rect 20487 2808 20904 2836
rect 20487 2805 20499 2808
rect 20441 2799 20499 2805
rect 20898 2796 20904 2808
rect 20956 2796 20962 2848
rect 23474 2796 23480 2848
rect 23532 2836 23538 2848
rect 24026 2836 24032 2848
rect 23532 2808 24032 2836
rect 23532 2796 23538 2808
rect 24026 2796 24032 2808
rect 24084 2796 24090 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1670 2632 1676 2644
rect 1631 2604 1676 2632
rect 1670 2592 1676 2604
rect 1728 2592 1734 2644
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 2406 2632 2412 2644
rect 1903 2604 2412 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 2406 2592 2412 2604
rect 2464 2592 2470 2644
rect 2866 2632 2872 2644
rect 2827 2604 2872 2632
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 3878 2632 3884 2644
rect 3839 2604 3884 2632
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 5442 2592 5448 2644
rect 5500 2632 5506 2644
rect 5721 2635 5779 2641
rect 5721 2632 5733 2635
rect 5500 2604 5733 2632
rect 5500 2592 5506 2604
rect 5721 2601 5733 2604
rect 5767 2632 5779 2635
rect 6733 2635 6791 2641
rect 6733 2632 6745 2635
rect 5767 2604 6745 2632
rect 5767 2601 5779 2604
rect 5721 2595 5779 2601
rect 6733 2601 6745 2604
rect 6779 2601 6791 2635
rect 6733 2595 6791 2601
rect 8478 2592 8484 2644
rect 8536 2632 8542 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8536 2604 9137 2632
rect 8536 2592 8542 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9766 2632 9772 2644
rect 9727 2604 9772 2632
rect 9125 2595 9183 2601
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 10134 2632 10140 2644
rect 10095 2604 10140 2632
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 10873 2635 10931 2641
rect 10873 2601 10885 2635
rect 10919 2632 10931 2635
rect 11054 2632 11060 2644
rect 10919 2604 11060 2632
rect 10919 2601 10931 2604
rect 10873 2595 10931 2601
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 13998 2632 14004 2644
rect 13959 2604 14004 2632
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 16850 2632 16856 2644
rect 16811 2604 16856 2632
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 18046 2632 18052 2644
rect 18007 2604 18052 2632
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 18138 2592 18144 2644
rect 18196 2632 18202 2644
rect 18506 2632 18512 2644
rect 18196 2604 18512 2632
rect 18196 2592 18202 2604
rect 18506 2592 18512 2604
rect 18564 2632 18570 2644
rect 19705 2635 19763 2641
rect 19705 2632 19717 2635
rect 18564 2604 19717 2632
rect 18564 2592 18570 2604
rect 19705 2601 19717 2604
rect 19751 2601 19763 2635
rect 19705 2595 19763 2601
rect 20625 2635 20683 2641
rect 20625 2601 20637 2635
rect 20671 2632 20683 2635
rect 20714 2632 20720 2644
rect 20671 2604 20720 2632
rect 20671 2601 20683 2604
rect 20625 2595 20683 2601
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 20898 2632 20904 2644
rect 20811 2604 20904 2632
rect 20898 2592 20904 2604
rect 20956 2632 20962 2644
rect 22002 2632 22008 2644
rect 20956 2604 22008 2632
rect 20956 2592 20962 2604
rect 2314 2564 2320 2576
rect 2275 2536 2320 2564
rect 2314 2524 2320 2536
rect 2372 2524 2378 2576
rect 2222 2496 2228 2508
rect 2183 2468 2228 2496
rect 2222 2456 2228 2468
rect 2280 2456 2286 2508
rect 3896 2496 3924 2592
rect 7460 2567 7518 2573
rect 7460 2533 7472 2567
rect 7506 2564 7518 2567
rect 7650 2564 7656 2576
rect 7506 2536 7656 2564
rect 7506 2533 7518 2536
rect 7460 2527 7518 2533
rect 7650 2524 7656 2536
rect 7708 2524 7714 2576
rect 4614 2505 4620 2508
rect 4341 2499 4399 2505
rect 4341 2496 4353 2499
rect 3896 2468 4353 2496
rect 4341 2465 4353 2468
rect 4387 2465 4399 2499
rect 4608 2496 4620 2505
rect 4341 2459 4399 2465
rect 4448 2468 4620 2496
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2428 2559 2431
rect 3234 2428 3240 2440
rect 2547 2400 3240 2428
rect 2547 2397 2559 2400
rect 2501 2391 2559 2397
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2428 3571 2431
rect 4448 2428 4476 2468
rect 4608 2459 4620 2468
rect 4614 2456 4620 2459
rect 4672 2456 4678 2508
rect 6641 2499 6699 2505
rect 6641 2465 6653 2499
rect 6687 2496 6699 2499
rect 6730 2496 6736 2508
rect 6687 2468 6736 2496
rect 6687 2465 6699 2468
rect 6641 2459 6699 2465
rect 6730 2456 6736 2468
rect 6788 2456 6794 2508
rect 7193 2499 7251 2505
rect 7193 2465 7205 2499
rect 7239 2496 7251 2499
rect 8496 2496 8524 2592
rect 9674 2524 9680 2576
rect 9732 2564 9738 2576
rect 10229 2567 10287 2573
rect 10229 2564 10241 2567
rect 9732 2536 10241 2564
rect 9732 2524 9738 2536
rect 10229 2533 10241 2536
rect 10275 2533 10287 2567
rect 10229 2527 10287 2533
rect 12069 2567 12127 2573
rect 12069 2533 12081 2567
rect 12115 2564 12127 2567
rect 12802 2564 12808 2576
rect 12115 2536 12808 2564
rect 12115 2533 12127 2536
rect 12069 2527 12127 2533
rect 12802 2524 12808 2536
rect 12860 2573 12866 2576
rect 12860 2567 12924 2573
rect 12860 2533 12878 2567
rect 12912 2533 12924 2567
rect 12860 2527 12924 2533
rect 12860 2524 12866 2527
rect 9950 2496 9956 2508
rect 7239 2468 8524 2496
rect 8680 2468 9956 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 3559 2400 4476 2428
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 8294 2320 8300 2372
rect 8352 2360 8358 2372
rect 8573 2363 8631 2369
rect 8573 2360 8585 2363
rect 8352 2332 8585 2360
rect 8352 2320 8358 2332
rect 8573 2329 8585 2332
rect 8619 2360 8631 2363
rect 8680 2360 8708 2468
rect 9950 2456 9956 2468
rect 10008 2456 10014 2508
rect 11238 2496 11244 2508
rect 11199 2468 11244 2496
rect 11238 2456 11244 2468
rect 11296 2496 11302 2508
rect 11425 2499 11483 2505
rect 11425 2496 11437 2499
rect 11296 2468 11437 2496
rect 11296 2456 11302 2468
rect 11425 2465 11437 2468
rect 11471 2465 11483 2499
rect 14458 2496 14464 2508
rect 11425 2459 11483 2465
rect 12636 2468 14464 2496
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 8619 2332 8708 2360
rect 9508 2400 10333 2428
rect 8619 2329 8631 2332
rect 8573 2323 8631 2329
rect 290 2252 296 2304
rect 348 2292 354 2304
rect 1302 2292 1308 2304
rect 348 2264 1308 2292
rect 348 2252 354 2264
rect 1302 2252 1308 2264
rect 1360 2292 1366 2304
rect 6546 2292 6552 2304
rect 1360 2264 6552 2292
rect 1360 2252 1366 2264
rect 6546 2252 6552 2264
rect 6604 2252 6610 2304
rect 9508 2301 9536 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 10870 2388 10876 2440
rect 10928 2428 10934 2440
rect 12636 2437 12664 2468
rect 14458 2456 14464 2468
rect 14516 2496 14522 2508
rect 15197 2499 15255 2505
rect 15197 2496 15209 2499
rect 14516 2468 15209 2496
rect 14516 2456 14522 2468
rect 15197 2465 15209 2468
rect 15243 2496 15255 2499
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15243 2468 15485 2496
rect 15243 2465 15255 2468
rect 15197 2459 15255 2465
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 15729 2499 15787 2505
rect 15729 2496 15741 2499
rect 15473 2459 15531 2465
rect 15580 2468 15741 2496
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 10928 2400 12357 2428
rect 10928 2388 10934 2400
rect 12345 2397 12357 2400
rect 12391 2428 12403 2431
rect 12621 2431 12679 2437
rect 12621 2428 12633 2431
rect 12391 2400 12633 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 12621 2397 12633 2400
rect 12667 2397 12679 2431
rect 12621 2391 12679 2397
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 15580 2428 15608 2468
rect 15729 2465 15741 2468
rect 15775 2496 15787 2499
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 15775 2468 17693 2496
rect 15775 2465 15787 2468
rect 15729 2459 15787 2465
rect 17681 2465 17693 2468
rect 17727 2465 17739 2499
rect 18064 2496 18092 2592
rect 18592 2567 18650 2573
rect 18592 2533 18604 2567
rect 18638 2564 18650 2567
rect 18690 2564 18696 2576
rect 18638 2536 18696 2564
rect 18638 2533 18650 2536
rect 18592 2527 18650 2533
rect 18690 2524 18696 2536
rect 18748 2524 18754 2576
rect 21192 2505 21220 2604
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 22554 2632 22560 2644
rect 22515 2604 22560 2632
rect 22554 2592 22560 2604
rect 22612 2592 22618 2644
rect 23750 2632 23756 2644
rect 23711 2604 23756 2632
rect 23750 2592 23756 2604
rect 23808 2592 23814 2644
rect 24210 2632 24216 2644
rect 24171 2604 24216 2632
rect 24210 2592 24216 2604
rect 24268 2592 24274 2644
rect 21444 2567 21502 2573
rect 21444 2533 21456 2567
rect 21490 2564 21502 2567
rect 21910 2564 21916 2576
rect 21490 2536 21916 2564
rect 21490 2533 21502 2536
rect 21444 2527 21502 2533
rect 21910 2524 21916 2536
rect 21968 2524 21974 2576
rect 23768 2564 23796 2592
rect 24581 2567 24639 2573
rect 24581 2564 24593 2567
rect 23768 2536 24593 2564
rect 24581 2533 24593 2536
rect 24627 2533 24639 2567
rect 24581 2527 24639 2533
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 18064 2468 18337 2496
rect 17681 2459 17739 2465
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 18325 2459 18383 2465
rect 21177 2499 21235 2505
rect 21177 2465 21189 2499
rect 21223 2465 21235 2499
rect 21177 2459 21235 2465
rect 14967 2400 15608 2428
rect 17696 2428 17724 2459
rect 18138 2428 18144 2440
rect 17696 2400 18144 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 18138 2388 18144 2400
rect 18196 2388 18202 2440
rect 23477 2431 23535 2437
rect 23477 2397 23489 2431
rect 23523 2428 23535 2431
rect 24486 2428 24492 2440
rect 23523 2400 24492 2428
rect 23523 2397 23535 2400
rect 23477 2391 23535 2397
rect 24486 2388 24492 2400
rect 24544 2428 24550 2440
rect 24673 2431 24731 2437
rect 24673 2428 24685 2431
rect 24544 2400 24685 2428
rect 24544 2388 24550 2400
rect 24673 2397 24685 2400
rect 24719 2397 24731 2431
rect 24673 2391 24731 2397
rect 24762 2388 24768 2440
rect 24820 2428 24826 2440
rect 25225 2431 25283 2437
rect 25225 2428 25237 2431
rect 24820 2400 25237 2428
rect 24820 2388 24826 2400
rect 25225 2397 25237 2400
rect 25271 2397 25283 2431
rect 25225 2391 25283 2397
rect 9766 2320 9772 2372
rect 9824 2360 9830 2372
rect 11698 2360 11704 2372
rect 9824 2332 11704 2360
rect 9824 2320 9830 2332
rect 11698 2320 11704 2332
rect 11756 2320 11762 2372
rect 6733 2295 6791 2301
rect 6733 2261 6745 2295
rect 6779 2292 6791 2295
rect 9493 2295 9551 2301
rect 9493 2292 9505 2295
rect 6779 2264 9505 2292
rect 6779 2261 6791 2264
rect 6733 2255 6791 2261
rect 9493 2261 9505 2264
rect 9539 2261 9551 2295
rect 11606 2292 11612 2304
rect 11567 2264 11612 2292
rect 9493 2255 9551 2261
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 2038 2048 2044 2100
rect 2096 2088 2102 2100
rect 6362 2088 6368 2100
rect 2096 2060 6368 2088
rect 2096 2048 2102 2060
rect 6362 2048 6368 2060
rect 6420 2048 6426 2100
rect 11790 1640 11796 1692
rect 11848 1680 11854 1692
rect 18874 1680 18880 1692
rect 11848 1652 18880 1680
rect 11848 1640 11854 1652
rect 18874 1640 18880 1652
rect 18932 1640 18938 1692
rect 3786 552 3792 604
rect 3844 592 3850 604
rect 4522 592 4528 604
rect 3844 564 4528 592
rect 3844 552 3850 564
rect 4522 552 4528 564
rect 4580 552 4586 604
rect 7742 552 7748 604
rect 7800 592 7806 604
rect 9030 592 9036 604
rect 7800 564 9036 592
rect 7800 552 7806 564
rect 9030 552 9036 564
rect 9088 552 9094 604
rect 10686 552 10692 604
rect 10744 592 10750 604
rect 10778 592 10784 604
rect 10744 564 10784 592
rect 10744 552 10750 564
rect 10778 552 10784 564
rect 10836 552 10842 604
rect 11330 552 11336 604
rect 11388 592 11394 604
rect 12342 592 12348 604
rect 11388 564 12348 592
rect 11388 552 11394 564
rect 12342 552 12348 564
rect 12400 552 12406 604
rect 21266 552 21272 604
rect 21324 592 21330 604
rect 21542 592 21548 604
rect 21324 564 21548 592
rect 21324 552 21330 564
rect 21542 552 21548 564
rect 21600 552 21606 604
rect 4338 484 4344 536
rect 4396 524 4402 536
rect 5166 524 5172 536
rect 4396 496 5172 524
rect 4396 484 4402 496
rect 5166 484 5172 496
rect 5224 484 5230 536
<< via1 >>
rect 17224 26800 17276 26852
rect 23480 26800 23532 26852
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 24768 23307 24820 23316
rect 24768 23273 24777 23307
rect 24777 23273 24811 23307
rect 24811 23273 24820 23307
rect 24768 23264 24820 23273
rect 24676 23128 24728 23180
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1584 22763 1636 22772
rect 1584 22729 1593 22763
rect 1593 22729 1627 22763
rect 1627 22729 1636 22763
rect 1584 22720 1636 22729
rect 1768 22516 1820 22568
rect 24584 22423 24636 22432
rect 24584 22389 24593 22423
rect 24593 22389 24627 22423
rect 24627 22389 24636 22423
rect 24584 22380 24636 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 24584 22176 24636 22228
rect 23848 22040 23900 22092
rect 24124 22040 24176 22092
rect 24768 21947 24820 21956
rect 24768 21913 24777 21947
rect 24777 21913 24811 21947
rect 24811 21913 24820 21947
rect 24768 21904 24820 21913
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 24676 21632 24728 21684
rect 23848 21471 23900 21480
rect 23848 21437 23857 21471
rect 23857 21437 23891 21471
rect 23891 21437 23900 21471
rect 23848 21428 23900 21437
rect 23940 21428 23992 21480
rect 24124 21292 24176 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1768 21131 1820 21140
rect 1768 21097 1777 21131
rect 1777 21097 1811 21131
rect 1811 21097 1820 21131
rect 1768 21088 1820 21097
rect 2504 20952 2556 21004
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1584 20587 1636 20596
rect 1584 20553 1593 20587
rect 1593 20553 1627 20587
rect 1627 20553 1636 20587
rect 1584 20544 1636 20553
rect 13268 20408 13320 20460
rect 13728 20272 13780 20324
rect 1768 20204 1820 20256
rect 2504 20204 2556 20256
rect 14740 20247 14792 20256
rect 14740 20213 14749 20247
rect 14749 20213 14783 20247
rect 14783 20213 14792 20247
rect 14740 20204 14792 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1492 20000 1544 20052
rect 2136 19864 2188 19916
rect 13268 19660 13320 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 2412 19227 2464 19236
rect 2412 19193 2421 19227
rect 2421 19193 2455 19227
rect 2455 19193 2464 19227
rect 2412 19184 2464 19193
rect 1400 19116 1452 19168
rect 2136 19116 2188 19168
rect 13268 19116 13320 19168
rect 14096 19184 14148 19236
rect 14924 19159 14976 19168
rect 14924 19125 14933 19159
rect 14933 19125 14967 19159
rect 14967 19125 14976 19159
rect 14924 19116 14976 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1768 18955 1820 18964
rect 1768 18921 1777 18955
rect 1777 18921 1811 18955
rect 1811 18921 1820 18955
rect 1768 18912 1820 18921
rect 2412 18776 2464 18828
rect 12808 18819 12860 18828
rect 12808 18785 12817 18819
rect 12817 18785 12851 18819
rect 12851 18785 12860 18819
rect 12808 18776 12860 18785
rect 14924 18776 14976 18828
rect 13084 18751 13136 18760
rect 12440 18683 12492 18692
rect 12440 18649 12449 18683
rect 12449 18649 12483 18683
rect 12483 18649 12492 18683
rect 12440 18640 12492 18649
rect 12348 18615 12400 18624
rect 12348 18581 12357 18615
rect 12357 18581 12391 18615
rect 12391 18581 12400 18615
rect 13084 18717 13093 18751
rect 13093 18717 13127 18751
rect 13127 18717 13136 18751
rect 13084 18708 13136 18717
rect 14004 18751 14056 18760
rect 14004 18717 14013 18751
rect 14013 18717 14047 18751
rect 14047 18717 14056 18751
rect 14004 18708 14056 18717
rect 12348 18572 12400 18581
rect 14096 18572 14148 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1584 18411 1636 18420
rect 1584 18377 1593 18411
rect 1593 18377 1627 18411
rect 1627 18377 1636 18411
rect 1584 18368 1636 18377
rect 2412 18411 2464 18420
rect 2412 18377 2421 18411
rect 2421 18377 2455 18411
rect 2455 18377 2464 18411
rect 2412 18368 2464 18377
rect 12808 18368 12860 18420
rect 2044 18071 2096 18080
rect 2044 18037 2053 18071
rect 2053 18037 2087 18071
rect 2087 18037 2096 18071
rect 2044 18028 2096 18037
rect 11060 18028 11112 18080
rect 13268 18164 13320 18216
rect 12716 18139 12768 18148
rect 12716 18105 12750 18139
rect 12750 18105 12768 18139
rect 12716 18096 12768 18105
rect 13084 18028 13136 18080
rect 14096 18028 14148 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1676 17824 1728 17876
rect 12808 17824 12860 17876
rect 14004 17824 14056 17876
rect 14740 17824 14792 17876
rect 24768 17867 24820 17876
rect 24768 17833 24777 17867
rect 24777 17833 24811 17867
rect 24811 17833 24820 17867
rect 24768 17824 24820 17833
rect 2320 17688 2372 17740
rect 10784 17688 10836 17740
rect 24676 17688 24728 17740
rect 11060 17663 11112 17672
rect 11060 17629 11069 17663
rect 11069 17629 11103 17663
rect 11103 17629 11112 17663
rect 11060 17620 11112 17629
rect 13544 17620 13596 17672
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 15660 17620 15712 17672
rect 12716 17552 12768 17604
rect 13636 17552 13688 17604
rect 11336 17484 11388 17536
rect 13360 17527 13412 17536
rect 13360 17493 13369 17527
rect 13369 17493 13403 17527
rect 13403 17493 13412 17527
rect 13360 17484 13412 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1492 17280 1544 17332
rect 2320 17323 2372 17332
rect 2320 17289 2329 17323
rect 2329 17289 2363 17323
rect 2363 17289 2372 17323
rect 2320 17280 2372 17289
rect 12440 17323 12492 17332
rect 12440 17289 12449 17323
rect 12449 17289 12483 17323
rect 12483 17289 12492 17323
rect 12440 17280 12492 17289
rect 24216 17280 24268 17332
rect 10140 17144 10192 17196
rect 11336 17187 11388 17196
rect 11336 17153 11345 17187
rect 11345 17153 11379 17187
rect 11379 17153 11388 17187
rect 11336 17144 11388 17153
rect 11796 17144 11848 17196
rect 10784 17076 10836 17128
rect 3332 16940 3384 16992
rect 10140 16983 10192 16992
rect 10140 16949 10149 16983
rect 10149 16949 10183 16983
rect 10183 16949 10192 16983
rect 10140 16940 10192 16949
rect 10692 16983 10744 16992
rect 10692 16949 10701 16983
rect 10701 16949 10735 16983
rect 10735 16949 10744 16983
rect 10692 16940 10744 16949
rect 11060 16983 11112 16992
rect 11060 16949 11069 16983
rect 11069 16949 11103 16983
rect 11103 16949 11112 16983
rect 11060 16940 11112 16949
rect 11244 16940 11296 16992
rect 12532 17144 12584 17196
rect 14372 17187 14424 17196
rect 14372 17153 14381 17187
rect 14381 17153 14415 17187
rect 14415 17153 14424 17187
rect 14372 17144 14424 17153
rect 13360 17076 13412 17128
rect 23664 17076 23716 17128
rect 13912 17008 13964 17060
rect 14740 17008 14792 17060
rect 12256 16983 12308 16992
rect 12256 16949 12265 16983
rect 12265 16949 12299 16983
rect 12299 16949 12308 16983
rect 12256 16940 12308 16949
rect 13544 16983 13596 16992
rect 13544 16949 13553 16983
rect 13553 16949 13587 16983
rect 13587 16949 13596 16983
rect 13544 16940 13596 16949
rect 15384 16940 15436 16992
rect 24400 16983 24452 16992
rect 24400 16949 24409 16983
rect 24409 16949 24443 16983
rect 24443 16949 24452 16983
rect 24400 16940 24452 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1584 16779 1636 16788
rect 1584 16745 1593 16779
rect 1593 16745 1627 16779
rect 1627 16745 1636 16779
rect 1584 16736 1636 16745
rect 10784 16736 10836 16788
rect 12532 16779 12584 16788
rect 12532 16745 12541 16779
rect 12541 16745 12575 16779
rect 12575 16745 12584 16779
rect 12532 16736 12584 16745
rect 13360 16736 13412 16788
rect 14004 16779 14056 16788
rect 14004 16745 14013 16779
rect 14013 16745 14047 16779
rect 14047 16745 14056 16779
rect 14004 16736 14056 16745
rect 14740 16736 14792 16788
rect 17040 16779 17092 16788
rect 14096 16668 14148 16720
rect 17040 16745 17049 16779
rect 17049 16745 17083 16779
rect 17083 16745 17092 16779
rect 17040 16736 17092 16745
rect 24400 16736 24452 16788
rect 24768 16779 24820 16788
rect 24768 16745 24777 16779
rect 24777 16745 24811 16779
rect 24811 16745 24820 16779
rect 24768 16736 24820 16745
rect 2412 16600 2464 16652
rect 9772 16600 9824 16652
rect 9220 16396 9272 16448
rect 10324 16439 10376 16448
rect 10324 16405 10333 16439
rect 10333 16405 10367 16439
rect 10367 16405 10376 16439
rect 10324 16396 10376 16405
rect 12164 16532 12216 16584
rect 13268 16532 13320 16584
rect 13636 16575 13688 16584
rect 13636 16541 13645 16575
rect 13645 16541 13679 16575
rect 13679 16541 13688 16575
rect 13636 16532 13688 16541
rect 14740 16532 14792 16584
rect 17132 16600 17184 16652
rect 23848 16600 23900 16652
rect 24124 16600 24176 16652
rect 13728 16464 13780 16516
rect 14096 16464 14148 16516
rect 11244 16396 11296 16448
rect 13084 16396 13136 16448
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 16764 16396 16816 16448
rect 17224 16396 17276 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2320 16192 2372 16244
rect 9680 16192 9732 16244
rect 13636 16192 13688 16244
rect 14740 16235 14792 16244
rect 14740 16201 14749 16235
rect 14749 16201 14783 16235
rect 14783 16201 14792 16235
rect 14740 16192 14792 16201
rect 16764 16235 16816 16244
rect 16764 16201 16773 16235
rect 16773 16201 16807 16235
rect 16807 16201 16816 16235
rect 16764 16192 16816 16201
rect 24124 16192 24176 16244
rect 3056 16124 3108 16176
rect 9772 16167 9824 16176
rect 9772 16133 9781 16167
rect 9781 16133 9815 16167
rect 9815 16133 9824 16167
rect 9772 16124 9824 16133
rect 11336 16124 11388 16176
rect 14004 16124 14056 16176
rect 18236 16167 18288 16176
rect 18236 16133 18245 16167
rect 18245 16133 18279 16167
rect 18279 16133 18288 16167
rect 18236 16124 18288 16133
rect 8392 16056 8444 16108
rect 10324 16056 10376 16108
rect 10692 16099 10744 16108
rect 10692 16065 10701 16099
rect 10701 16065 10735 16099
rect 10735 16065 10744 16099
rect 10692 16056 10744 16065
rect 10784 16099 10836 16108
rect 10784 16065 10793 16099
rect 10793 16065 10827 16099
rect 10827 16065 10836 16099
rect 13912 16099 13964 16108
rect 10784 16056 10836 16065
rect 13912 16065 13921 16099
rect 13921 16065 13955 16099
rect 13955 16065 13964 16099
rect 13912 16056 13964 16065
rect 14372 16056 14424 16108
rect 15384 15988 15436 16040
rect 17684 15988 17736 16040
rect 23848 16031 23900 16040
rect 23848 15997 23857 16031
rect 23857 15997 23891 16031
rect 23891 15997 23900 16031
rect 23848 15988 23900 15997
rect 7564 15920 7616 15972
rect 10784 15920 10836 15972
rect 13544 15920 13596 15972
rect 15568 15920 15620 15972
rect 2044 15895 2096 15904
rect 2044 15861 2053 15895
rect 2053 15861 2087 15895
rect 2087 15861 2096 15895
rect 2044 15852 2096 15861
rect 2412 15895 2464 15904
rect 2412 15861 2421 15895
rect 2421 15861 2455 15895
rect 2455 15861 2464 15895
rect 2412 15852 2464 15861
rect 8392 15852 8444 15904
rect 8668 15895 8720 15904
rect 8668 15861 8677 15895
rect 8677 15861 8711 15895
rect 8711 15861 8720 15895
rect 8668 15852 8720 15861
rect 9036 15895 9088 15904
rect 9036 15861 9045 15895
rect 9045 15861 9079 15895
rect 9079 15861 9088 15895
rect 9036 15852 9088 15861
rect 9220 15852 9272 15904
rect 11244 15895 11296 15904
rect 11244 15861 11253 15895
rect 11253 15861 11287 15895
rect 11287 15861 11296 15895
rect 11244 15852 11296 15861
rect 12164 15895 12216 15904
rect 12164 15861 12173 15895
rect 12173 15861 12207 15895
rect 12207 15861 12216 15895
rect 12164 15852 12216 15861
rect 13268 15852 13320 15904
rect 13360 15852 13412 15904
rect 16580 15852 16632 15904
rect 17132 15895 17184 15904
rect 17132 15861 17141 15895
rect 17141 15861 17175 15895
rect 17175 15861 17184 15895
rect 17132 15852 17184 15861
rect 23848 15852 23900 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1400 15648 1452 15700
rect 8668 15648 8720 15700
rect 13820 15648 13872 15700
rect 14096 15691 14148 15700
rect 14096 15657 14105 15691
rect 14105 15657 14139 15691
rect 14139 15657 14148 15691
rect 14096 15648 14148 15657
rect 14372 15648 14424 15700
rect 15384 15648 15436 15700
rect 19432 15648 19484 15700
rect 24676 15648 24728 15700
rect 11060 15580 11112 15632
rect 16028 15580 16080 15632
rect 1860 15512 1912 15564
rect 8668 15512 8720 15564
rect 8300 15444 8352 15496
rect 9680 15487 9732 15496
rect 9680 15453 9689 15487
rect 9689 15453 9723 15487
rect 9723 15453 9732 15487
rect 9680 15444 9732 15453
rect 10232 15444 10284 15496
rect 11244 15512 11296 15564
rect 14004 15555 14056 15564
rect 14004 15521 14013 15555
rect 14013 15521 14047 15555
rect 14047 15521 14056 15555
rect 14004 15512 14056 15521
rect 16396 15512 16448 15564
rect 17592 15512 17644 15564
rect 18420 15555 18472 15564
rect 18420 15521 18429 15555
rect 18429 15521 18463 15555
rect 18463 15521 18472 15555
rect 18420 15512 18472 15521
rect 19340 15512 19392 15564
rect 23940 15512 23992 15564
rect 24860 15512 24912 15564
rect 11888 15444 11940 15496
rect 12256 15444 12308 15496
rect 13360 15444 13412 15496
rect 13544 15444 13596 15496
rect 15384 15444 15436 15496
rect 15844 15487 15896 15496
rect 15844 15453 15853 15487
rect 15853 15453 15887 15487
rect 15887 15453 15896 15487
rect 17316 15487 17368 15496
rect 15844 15444 15896 15453
rect 17316 15453 17325 15487
rect 17325 15453 17359 15487
rect 17359 15453 17368 15487
rect 17316 15444 17368 15453
rect 8024 15419 8076 15428
rect 8024 15385 8033 15419
rect 8033 15385 8067 15419
rect 8067 15385 8076 15419
rect 8024 15376 8076 15385
rect 13636 15419 13688 15428
rect 13636 15385 13645 15419
rect 13645 15385 13679 15419
rect 13679 15385 13688 15419
rect 13636 15376 13688 15385
rect 16580 15376 16632 15428
rect 22284 15444 22336 15496
rect 4252 15351 4304 15360
rect 4252 15317 4261 15351
rect 4261 15317 4295 15351
rect 4295 15317 4304 15351
rect 4252 15308 4304 15317
rect 11336 15308 11388 15360
rect 15292 15351 15344 15360
rect 15292 15317 15301 15351
rect 15301 15317 15335 15351
rect 15335 15317 15344 15351
rect 15292 15308 15344 15317
rect 16488 15308 16540 15360
rect 18236 15308 18288 15360
rect 22468 15308 22520 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1952 15104 2004 15156
rect 8300 15104 8352 15156
rect 9680 15104 9732 15156
rect 13544 15147 13596 15156
rect 10784 15079 10836 15088
rect 10784 15045 10793 15079
rect 10793 15045 10827 15079
rect 10827 15045 10836 15079
rect 10784 15036 10836 15045
rect 5724 14968 5776 15020
rect 4252 14943 4304 14952
rect 4252 14909 4261 14943
rect 4261 14909 4295 14943
rect 4295 14909 4304 14943
rect 4252 14900 4304 14909
rect 13544 15113 13553 15147
rect 13553 15113 13587 15147
rect 13587 15113 13596 15147
rect 13544 15104 13596 15113
rect 12808 15036 12860 15088
rect 14372 15104 14424 15156
rect 16028 15147 16080 15156
rect 16028 15113 16037 15147
rect 16037 15113 16071 15147
rect 16071 15113 16080 15147
rect 16028 15104 16080 15113
rect 16120 15104 16172 15156
rect 16396 15147 16448 15156
rect 16396 15113 16405 15147
rect 16405 15113 16439 15147
rect 16439 15113 16448 15147
rect 16396 15104 16448 15113
rect 17316 15147 17368 15156
rect 17316 15113 17325 15147
rect 17325 15113 17359 15147
rect 17359 15113 17368 15147
rect 17316 15104 17368 15113
rect 24768 15147 24820 15156
rect 24768 15113 24777 15147
rect 24777 15113 24811 15147
rect 24811 15113 24820 15147
rect 24768 15104 24820 15113
rect 11336 15011 11388 15020
rect 11336 14977 11345 15011
rect 11345 14977 11379 15011
rect 11379 14977 11388 15011
rect 11336 14968 11388 14977
rect 11704 14968 11756 15020
rect 12624 14968 12676 15020
rect 12992 15011 13044 15020
rect 12992 14977 13001 15011
rect 13001 14977 13035 15011
rect 13035 14977 13044 15011
rect 12992 14968 13044 14977
rect 20444 15036 20496 15088
rect 1860 14764 1912 14816
rect 2504 14807 2556 14816
rect 2504 14773 2513 14807
rect 2513 14773 2547 14807
rect 2547 14773 2556 14807
rect 2504 14764 2556 14773
rect 3056 14764 3108 14816
rect 3884 14807 3936 14816
rect 3884 14773 3893 14807
rect 3893 14773 3927 14807
rect 3927 14773 3936 14807
rect 3884 14764 3936 14773
rect 6920 14807 6972 14816
rect 6920 14773 6929 14807
rect 6929 14773 6963 14807
rect 6963 14773 6972 14807
rect 6920 14764 6972 14773
rect 7104 14764 7156 14816
rect 8576 14832 8628 14884
rect 9680 14832 9732 14884
rect 10232 14875 10284 14884
rect 10232 14841 10241 14875
rect 10241 14841 10275 14875
rect 10275 14841 10284 14875
rect 10232 14832 10284 14841
rect 12348 14832 12400 14884
rect 16304 14900 16356 14952
rect 16488 14943 16540 14952
rect 16488 14909 16497 14943
rect 16497 14909 16531 14943
rect 16531 14909 16540 14943
rect 16488 14900 16540 14909
rect 18880 14900 18932 14952
rect 9956 14764 10008 14816
rect 11244 14807 11296 14816
rect 11244 14773 11253 14807
rect 11253 14773 11287 14807
rect 11287 14773 11296 14807
rect 11244 14764 11296 14773
rect 12440 14807 12492 14816
rect 12440 14773 12449 14807
rect 12449 14773 12483 14807
rect 12483 14773 12492 14807
rect 12440 14764 12492 14773
rect 12624 14764 12676 14816
rect 14096 14832 14148 14884
rect 16580 14832 16632 14884
rect 17960 14832 18012 14884
rect 18420 14832 18472 14884
rect 19340 14900 19392 14952
rect 20352 14943 20404 14952
rect 20352 14909 20361 14943
rect 20361 14909 20395 14943
rect 20395 14909 20404 14943
rect 20352 14900 20404 14909
rect 15200 14764 15252 14816
rect 16856 14764 16908 14816
rect 17592 14764 17644 14816
rect 18696 14764 18748 14816
rect 20536 14807 20588 14816
rect 20536 14773 20545 14807
rect 20545 14773 20579 14807
rect 20579 14773 20588 14807
rect 20536 14764 20588 14773
rect 21548 14807 21600 14816
rect 21548 14773 21557 14807
rect 21557 14773 21591 14807
rect 21591 14773 21600 14807
rect 21548 14764 21600 14773
rect 22744 14807 22796 14816
rect 22744 14773 22753 14807
rect 22753 14773 22787 14807
rect 22787 14773 22796 14807
rect 22744 14764 22796 14773
rect 24124 14900 24176 14952
rect 23572 14832 23624 14884
rect 24952 14832 25004 14884
rect 23204 14764 23256 14816
rect 23940 14807 23992 14816
rect 23940 14773 23949 14807
rect 23949 14773 23983 14807
rect 23983 14773 23992 14807
rect 23940 14764 23992 14773
rect 24124 14764 24176 14816
rect 24860 14764 24912 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 2504 14560 2556 14612
rect 4252 14560 4304 14612
rect 11060 14603 11112 14612
rect 11060 14569 11069 14603
rect 11069 14569 11103 14603
rect 11103 14569 11112 14603
rect 11060 14560 11112 14569
rect 11336 14560 11388 14612
rect 13728 14603 13780 14612
rect 13728 14569 13737 14603
rect 13737 14569 13771 14603
rect 13771 14569 13780 14603
rect 13728 14560 13780 14569
rect 14004 14560 14056 14612
rect 14832 14560 14884 14612
rect 15292 14560 15344 14612
rect 15844 14560 15896 14612
rect 17316 14603 17368 14612
rect 17316 14569 17325 14603
rect 17325 14569 17359 14603
rect 17359 14569 17368 14603
rect 17316 14560 17368 14569
rect 17776 14560 17828 14612
rect 18604 14603 18656 14612
rect 18604 14569 18613 14603
rect 18613 14569 18647 14603
rect 18647 14569 18656 14603
rect 18604 14560 18656 14569
rect 24216 14560 24268 14612
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 3884 14492 3936 14544
rect 4160 14492 4212 14544
rect 2780 14424 2832 14476
rect 3516 14424 3568 14476
rect 4436 14467 4488 14476
rect 4436 14433 4445 14467
rect 4445 14433 4479 14467
rect 4479 14433 4488 14467
rect 4436 14424 4488 14433
rect 5724 14492 5776 14544
rect 14096 14535 14148 14544
rect 14096 14501 14105 14535
rect 14105 14501 14139 14535
rect 14139 14501 14148 14535
rect 14096 14492 14148 14501
rect 15660 14535 15712 14544
rect 15660 14501 15669 14535
rect 15669 14501 15703 14535
rect 15703 14501 15712 14535
rect 15660 14492 15712 14501
rect 16580 14492 16632 14544
rect 9956 14467 10008 14476
rect 9956 14433 9990 14467
rect 9990 14433 10008 14467
rect 9956 14424 10008 14433
rect 12256 14424 12308 14476
rect 14188 14467 14240 14476
rect 14188 14433 14197 14467
rect 14197 14433 14231 14467
rect 14231 14433 14240 14467
rect 14188 14424 14240 14433
rect 17224 14467 17276 14476
rect 17224 14433 17233 14467
rect 17233 14433 17267 14467
rect 17267 14433 17276 14467
rect 17224 14424 17276 14433
rect 2780 14288 2832 14340
rect 8208 14399 8260 14408
rect 4528 14288 4580 14340
rect 8208 14365 8217 14399
rect 8217 14365 8251 14399
rect 8251 14365 8260 14399
rect 8208 14356 8260 14365
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 12624 14399 12676 14408
rect 12624 14365 12633 14399
rect 12633 14365 12667 14399
rect 12667 14365 12676 14399
rect 12624 14356 12676 14365
rect 8576 14288 8628 14340
rect 11060 14288 11112 14340
rect 12992 14356 13044 14408
rect 13360 14356 13412 14408
rect 15200 14356 15252 14408
rect 15384 14356 15436 14408
rect 15752 14356 15804 14408
rect 17776 14424 17828 14476
rect 19432 14424 19484 14476
rect 20168 14424 20220 14476
rect 20628 14424 20680 14476
rect 22560 14467 22612 14476
rect 22560 14433 22569 14467
rect 22569 14433 22603 14467
rect 22603 14433 22612 14467
rect 22560 14424 22612 14433
rect 23572 14467 23624 14476
rect 23572 14433 23581 14467
rect 23581 14433 23615 14467
rect 23615 14433 23624 14467
rect 23572 14424 23624 14433
rect 24676 14424 24728 14476
rect 17592 14288 17644 14340
rect 1952 14263 2004 14272
rect 1952 14229 1961 14263
rect 1961 14229 1995 14263
rect 1995 14229 2004 14263
rect 1952 14220 2004 14229
rect 3148 14263 3200 14272
rect 3148 14229 3157 14263
rect 3157 14229 3191 14263
rect 3191 14229 3200 14263
rect 3148 14220 3200 14229
rect 3424 14263 3476 14272
rect 3424 14229 3433 14263
rect 3433 14229 3467 14263
rect 3467 14229 3476 14263
rect 3424 14220 3476 14229
rect 7288 14220 7340 14272
rect 8668 14263 8720 14272
rect 8668 14229 8677 14263
rect 8677 14229 8711 14263
rect 8711 14229 8720 14263
rect 8668 14220 8720 14229
rect 11980 14263 12032 14272
rect 11980 14229 11989 14263
rect 11989 14229 12023 14263
rect 12023 14229 12032 14263
rect 11980 14220 12032 14229
rect 14372 14263 14424 14272
rect 14372 14229 14381 14263
rect 14381 14229 14415 14263
rect 14415 14229 14424 14263
rect 14372 14220 14424 14229
rect 16396 14263 16448 14272
rect 16396 14229 16405 14263
rect 16405 14229 16439 14263
rect 16439 14229 16448 14263
rect 16396 14220 16448 14229
rect 16580 14220 16632 14272
rect 16764 14220 16816 14272
rect 18420 14220 18472 14272
rect 19248 14220 19300 14272
rect 19984 14220 20036 14272
rect 20260 14220 20312 14272
rect 22928 14220 22980 14272
rect 23756 14263 23808 14272
rect 23756 14229 23765 14263
rect 23765 14229 23799 14263
rect 23799 14229 23808 14263
rect 23756 14220 23808 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1400 14016 1452 14068
rect 2228 14016 2280 14068
rect 4436 14016 4488 14068
rect 5540 14016 5592 14068
rect 9680 14059 9732 14068
rect 9680 14025 9689 14059
rect 9689 14025 9723 14059
rect 9723 14025 9732 14059
rect 9680 14016 9732 14025
rect 10692 14016 10744 14068
rect 11060 14016 11112 14068
rect 12256 14059 12308 14068
rect 12256 14025 12265 14059
rect 12265 14025 12299 14059
rect 12299 14025 12308 14059
rect 12256 14016 12308 14025
rect 15660 14016 15712 14068
rect 15752 14059 15804 14068
rect 15752 14025 15761 14059
rect 15761 14025 15795 14059
rect 15795 14025 15804 14059
rect 15752 14016 15804 14025
rect 17316 14016 17368 14068
rect 18052 14059 18104 14068
rect 18052 14025 18061 14059
rect 18061 14025 18095 14059
rect 18095 14025 18104 14059
rect 18052 14016 18104 14025
rect 19432 14059 19484 14068
rect 19432 14025 19441 14059
rect 19441 14025 19475 14059
rect 19475 14025 19484 14059
rect 19432 14016 19484 14025
rect 22192 14016 22244 14068
rect 22560 14016 22612 14068
rect 2136 13948 2188 14000
rect 4160 13991 4212 14000
rect 4160 13957 4169 13991
rect 4169 13957 4203 13991
rect 4203 13957 4212 13991
rect 12624 13991 12676 14000
rect 4160 13948 4212 13957
rect 10968 13923 11020 13932
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 10968 13880 11020 13889
rect 11060 13880 11112 13932
rect 11336 13880 11388 13932
rect 12624 13957 12633 13991
rect 12633 13957 12667 13991
rect 12667 13957 12676 13991
rect 12624 13948 12676 13957
rect 16488 13948 16540 14000
rect 24768 13991 24820 14000
rect 24768 13957 24777 13991
rect 24777 13957 24811 13991
rect 24811 13957 24820 13991
rect 24768 13948 24820 13957
rect 12532 13880 12584 13932
rect 2044 13855 2096 13864
rect 2044 13821 2053 13855
rect 2053 13821 2087 13855
rect 2087 13821 2096 13855
rect 2044 13812 2096 13821
rect 2136 13812 2188 13864
rect 4528 13855 4580 13864
rect 4528 13821 4551 13855
rect 4551 13821 4580 13855
rect 4528 13812 4580 13821
rect 5540 13812 5592 13864
rect 7104 13855 7156 13864
rect 7104 13821 7113 13855
rect 7113 13821 7147 13855
rect 7147 13821 7156 13855
rect 7104 13812 7156 13821
rect 7288 13812 7340 13864
rect 8116 13744 8168 13796
rect 9956 13812 10008 13864
rect 11980 13812 12032 13864
rect 12808 13812 12860 13864
rect 16396 13880 16448 13932
rect 16672 13923 16724 13932
rect 16672 13889 16681 13923
rect 16681 13889 16715 13923
rect 16715 13889 16724 13923
rect 16672 13880 16724 13889
rect 18604 13923 18656 13932
rect 18604 13889 18613 13923
rect 18613 13889 18647 13923
rect 18647 13889 18656 13923
rect 18604 13880 18656 13889
rect 13360 13855 13412 13864
rect 13360 13821 13394 13855
rect 13394 13821 13412 13855
rect 13360 13812 13412 13821
rect 15200 13812 15252 13864
rect 17224 13812 17276 13864
rect 14648 13744 14700 13796
rect 15936 13744 15988 13796
rect 16764 13744 16816 13796
rect 19248 13812 19300 13864
rect 20168 13855 20220 13864
rect 20168 13821 20177 13855
rect 20177 13821 20211 13855
rect 20211 13821 20220 13855
rect 20168 13812 20220 13821
rect 21640 13812 21692 13864
rect 23020 13855 23072 13864
rect 23020 13821 23029 13855
rect 23029 13821 23063 13855
rect 23063 13821 23072 13855
rect 23020 13812 23072 13821
rect 23572 13812 23624 13864
rect 24584 13855 24636 13864
rect 24584 13821 24593 13855
rect 24593 13821 24627 13855
rect 24627 13821 24636 13855
rect 24584 13812 24636 13821
rect 2688 13719 2740 13728
rect 2688 13685 2697 13719
rect 2697 13685 2731 13719
rect 2731 13685 2740 13719
rect 2688 13676 2740 13685
rect 3608 13676 3660 13728
rect 8576 13719 8628 13728
rect 8576 13685 8585 13719
rect 8585 13685 8619 13719
rect 8619 13685 8628 13719
rect 8576 13676 8628 13685
rect 14280 13676 14332 13728
rect 18420 13719 18472 13728
rect 18420 13685 18429 13719
rect 18429 13685 18463 13719
rect 18463 13685 18472 13719
rect 18420 13676 18472 13685
rect 20628 13676 20680 13728
rect 22652 13676 22704 13728
rect 24400 13719 24452 13728
rect 24400 13685 24409 13719
rect 24409 13685 24443 13719
rect 24443 13685 24452 13719
rect 24400 13676 24452 13685
rect 24676 13676 24728 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1400 13472 1452 13524
rect 2688 13472 2740 13524
rect 5540 13472 5592 13524
rect 7288 13515 7340 13524
rect 7288 13481 7297 13515
rect 7297 13481 7331 13515
rect 7331 13481 7340 13515
rect 7288 13472 7340 13481
rect 7564 13515 7616 13524
rect 7564 13481 7573 13515
rect 7573 13481 7607 13515
rect 7607 13481 7616 13515
rect 7564 13472 7616 13481
rect 9128 13472 9180 13524
rect 6644 13404 6696 13456
rect 7748 13404 7800 13456
rect 10968 13472 11020 13524
rect 12256 13515 12308 13524
rect 12256 13481 12265 13515
rect 12265 13481 12299 13515
rect 12299 13481 12308 13515
rect 12256 13472 12308 13481
rect 12808 13472 12860 13524
rect 11152 13404 11204 13456
rect 2044 13336 2096 13388
rect 2504 13379 2556 13388
rect 2504 13345 2513 13379
rect 2513 13345 2547 13379
rect 2547 13345 2556 13379
rect 2504 13336 2556 13345
rect 4160 13336 4212 13388
rect 5080 13336 5132 13388
rect 7564 13336 7616 13388
rect 9312 13336 9364 13388
rect 10692 13336 10744 13388
rect 10968 13336 11020 13388
rect 12624 13336 12676 13388
rect 14188 13472 14240 13524
rect 14372 13472 14424 13524
rect 15108 13515 15160 13524
rect 15108 13481 15117 13515
rect 15117 13481 15151 13515
rect 15151 13481 15160 13515
rect 15108 13472 15160 13481
rect 15844 13515 15896 13524
rect 15844 13481 15853 13515
rect 15853 13481 15887 13515
rect 15887 13481 15896 13515
rect 15844 13472 15896 13481
rect 16672 13472 16724 13524
rect 17316 13472 17368 13524
rect 24400 13472 24452 13524
rect 24768 13515 24820 13524
rect 24768 13481 24777 13515
rect 24777 13481 24811 13515
rect 24811 13481 24820 13515
rect 24768 13472 24820 13481
rect 19432 13404 19484 13456
rect 19800 13404 19852 13456
rect 13636 13336 13688 13388
rect 13912 13379 13964 13388
rect 13912 13345 13921 13379
rect 13921 13345 13955 13379
rect 13955 13345 13964 13379
rect 13912 13336 13964 13345
rect 2872 13268 2924 13320
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 12532 13311 12584 13320
rect 10232 13268 10284 13277
rect 12532 13277 12541 13311
rect 12541 13277 12575 13311
rect 12575 13277 12584 13311
rect 12532 13268 12584 13277
rect 2596 13200 2648 13252
rect 14464 13336 14516 13388
rect 14188 13311 14240 13320
rect 14188 13277 14197 13311
rect 14197 13277 14231 13311
rect 14231 13277 14240 13311
rect 16580 13336 16632 13388
rect 18788 13336 18840 13388
rect 23480 13336 23532 13388
rect 24216 13336 24268 13388
rect 16028 13311 16080 13320
rect 14188 13268 14240 13277
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 18972 13311 19024 13320
rect 18972 13277 18981 13311
rect 18981 13277 19015 13311
rect 19015 13277 19024 13311
rect 18972 13268 19024 13277
rect 19064 13311 19116 13320
rect 19064 13277 19073 13311
rect 19073 13277 19107 13311
rect 19107 13277 19116 13311
rect 19064 13268 19116 13277
rect 19432 13268 19484 13320
rect 20076 13268 20128 13320
rect 21088 13268 21140 13320
rect 23112 13268 23164 13320
rect 23848 13268 23900 13320
rect 24768 13268 24820 13320
rect 14280 13200 14332 13252
rect 14556 13200 14608 13252
rect 20352 13200 20404 13252
rect 1676 13132 1728 13184
rect 2780 13132 2832 13184
rect 3884 13175 3936 13184
rect 3884 13141 3893 13175
rect 3893 13141 3927 13175
rect 3927 13141 3936 13175
rect 3884 13132 3936 13141
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 9404 13175 9456 13184
rect 9404 13141 9413 13175
rect 9413 13141 9447 13175
rect 9447 13141 9456 13175
rect 9404 13132 9456 13141
rect 9772 13132 9824 13184
rect 11336 13175 11388 13184
rect 11336 13141 11345 13175
rect 11345 13141 11379 13175
rect 11379 13141 11388 13175
rect 11336 13132 11388 13141
rect 12808 13132 12860 13184
rect 15568 13175 15620 13184
rect 15568 13141 15577 13175
rect 15577 13141 15611 13175
rect 15611 13141 15620 13175
rect 15568 13132 15620 13141
rect 18328 13132 18380 13184
rect 18512 13175 18564 13184
rect 18512 13141 18521 13175
rect 18521 13141 18555 13175
rect 18555 13141 18564 13175
rect 18512 13132 18564 13141
rect 19616 13175 19668 13184
rect 19616 13141 19625 13175
rect 19625 13141 19659 13175
rect 19659 13141 19668 13175
rect 19616 13132 19668 13141
rect 20076 13175 20128 13184
rect 20076 13141 20085 13175
rect 20085 13141 20119 13175
rect 20119 13141 20128 13175
rect 20076 13132 20128 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1492 12928 1544 12980
rect 1676 12928 1728 12980
rect 1860 12928 1912 12980
rect 3056 12971 3108 12980
rect 3056 12937 3065 12971
rect 3065 12937 3099 12971
rect 3099 12937 3108 12971
rect 3056 12928 3108 12937
rect 6644 12971 6696 12980
rect 6644 12937 6653 12971
rect 6653 12937 6687 12971
rect 6687 12937 6696 12971
rect 6644 12928 6696 12937
rect 7564 12928 7616 12980
rect 9128 12971 9180 12980
rect 9128 12937 9137 12971
rect 9137 12937 9171 12971
rect 9171 12937 9180 12971
rect 9128 12928 9180 12937
rect 9312 12928 9364 12980
rect 11152 12971 11204 12980
rect 11152 12937 11161 12971
rect 11161 12937 11195 12971
rect 11195 12937 11204 12971
rect 11152 12928 11204 12937
rect 12256 12928 12308 12980
rect 13912 12928 13964 12980
rect 14648 12971 14700 12980
rect 14648 12937 14657 12971
rect 14657 12937 14691 12971
rect 14691 12937 14700 12971
rect 14648 12928 14700 12937
rect 15936 12928 15988 12980
rect 16028 12928 16080 12980
rect 16580 12971 16632 12980
rect 16580 12937 16589 12971
rect 16589 12937 16623 12971
rect 16623 12937 16632 12971
rect 16580 12928 16632 12937
rect 17776 12928 17828 12980
rect 19340 12928 19392 12980
rect 20720 12971 20772 12980
rect 20720 12937 20729 12971
rect 20729 12937 20763 12971
rect 20763 12937 20772 12971
rect 20720 12928 20772 12937
rect 20904 12928 20956 12980
rect 23480 12928 23532 12980
rect 24952 12928 25004 12980
rect 2320 12792 2372 12844
rect 2596 12792 2648 12844
rect 3148 12792 3200 12844
rect 3608 12835 3660 12844
rect 3608 12801 3617 12835
rect 3617 12801 3651 12835
rect 3651 12801 3660 12835
rect 3608 12792 3660 12801
rect 5080 12792 5132 12844
rect 8576 12792 8628 12844
rect 10232 12835 10284 12844
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10232 12792 10284 12801
rect 15568 12792 15620 12844
rect 15936 12792 15988 12844
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 2044 12767 2096 12776
rect 2044 12733 2053 12767
rect 2053 12733 2087 12767
rect 2087 12733 2096 12767
rect 2044 12724 2096 12733
rect 3424 12767 3476 12776
rect 3424 12733 3433 12767
rect 3433 12733 3467 12767
rect 3467 12733 3476 12767
rect 3424 12724 3476 12733
rect 4160 12724 4212 12776
rect 7380 12724 7432 12776
rect 8208 12724 8260 12776
rect 11336 12767 11388 12776
rect 11336 12733 11345 12767
rect 11345 12733 11379 12767
rect 11379 12733 11388 12767
rect 11336 12724 11388 12733
rect 12808 12724 12860 12776
rect 13360 12724 13412 12776
rect 14004 12767 14056 12776
rect 14004 12733 14013 12767
rect 14013 12733 14047 12767
rect 14047 12733 14056 12767
rect 14004 12724 14056 12733
rect 16580 12724 16632 12776
rect 17960 12860 18012 12912
rect 24216 12860 24268 12912
rect 17132 12792 17184 12844
rect 20076 12792 20128 12844
rect 3608 12656 3660 12708
rect 4988 12699 5040 12708
rect 4988 12665 4997 12699
rect 4997 12665 5031 12699
rect 5031 12665 5040 12699
rect 4988 12656 5040 12665
rect 1400 12588 1452 12640
rect 2044 12588 2096 12640
rect 2228 12588 2280 12640
rect 3332 12588 3384 12640
rect 7472 12656 7524 12708
rect 9864 12656 9916 12708
rect 7932 12588 7984 12640
rect 8576 12631 8628 12640
rect 8576 12597 8585 12631
rect 8585 12597 8619 12631
rect 8619 12597 8628 12631
rect 8576 12588 8628 12597
rect 9680 12631 9732 12640
rect 9680 12597 9689 12631
rect 9689 12597 9723 12631
rect 9723 12597 9732 12631
rect 9680 12588 9732 12597
rect 10048 12631 10100 12640
rect 10048 12597 10057 12631
rect 10057 12597 10091 12631
rect 10091 12597 10100 12631
rect 10048 12588 10100 12597
rect 11244 12656 11296 12708
rect 11336 12588 11388 12640
rect 12532 12588 12584 12640
rect 15292 12656 15344 12708
rect 16672 12656 16724 12708
rect 18144 12656 18196 12708
rect 19064 12699 19116 12708
rect 19064 12665 19073 12699
rect 19073 12665 19107 12699
rect 19107 12665 19116 12699
rect 19064 12656 19116 12665
rect 15476 12588 15528 12640
rect 15660 12631 15712 12640
rect 15660 12597 15669 12631
rect 15669 12597 15703 12631
rect 15703 12597 15712 12631
rect 15660 12588 15712 12597
rect 18052 12631 18104 12640
rect 18052 12597 18061 12631
rect 18061 12597 18095 12631
rect 18095 12597 18104 12631
rect 18052 12588 18104 12597
rect 18328 12588 18380 12640
rect 19248 12588 19300 12640
rect 19616 12724 19668 12776
rect 22560 12767 22612 12776
rect 22560 12733 22569 12767
rect 22569 12733 22603 12767
rect 22603 12733 22612 12767
rect 22560 12724 22612 12733
rect 24124 12724 24176 12776
rect 20352 12656 20404 12708
rect 21180 12631 21232 12640
rect 21180 12597 21189 12631
rect 21189 12597 21223 12631
rect 21223 12597 21232 12631
rect 21180 12588 21232 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1492 12384 1544 12436
rect 1768 12384 1820 12436
rect 2688 12384 2740 12436
rect 3148 12384 3200 12436
rect 3516 12384 3568 12436
rect 4436 12384 4488 12436
rect 7748 12427 7800 12436
rect 7748 12393 7757 12427
rect 7757 12393 7791 12427
rect 7791 12393 7800 12427
rect 7748 12384 7800 12393
rect 8116 12384 8168 12436
rect 7104 12316 7156 12368
rect 1952 12248 2004 12300
rect 2044 12248 2096 12300
rect 3332 12248 3384 12300
rect 4252 12248 4304 12300
rect 6184 12248 6236 12300
rect 9588 12384 9640 12436
rect 11796 12427 11848 12436
rect 11796 12393 11805 12427
rect 11805 12393 11839 12427
rect 11839 12393 11848 12427
rect 11796 12384 11848 12393
rect 12440 12427 12492 12436
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 14188 12427 14240 12436
rect 12440 12384 12492 12393
rect 14188 12393 14197 12427
rect 14197 12393 14231 12427
rect 14231 12393 14240 12427
rect 14188 12384 14240 12393
rect 14464 12384 14516 12436
rect 15292 12427 15344 12436
rect 15292 12393 15301 12427
rect 15301 12393 15335 12427
rect 15335 12393 15344 12427
rect 15292 12384 15344 12393
rect 15844 12427 15896 12436
rect 15844 12393 15853 12427
rect 15853 12393 15887 12427
rect 15887 12393 15896 12427
rect 15844 12384 15896 12393
rect 17960 12384 18012 12436
rect 19064 12427 19116 12436
rect 19064 12393 19073 12427
rect 19073 12393 19107 12427
rect 19107 12393 19116 12427
rect 19064 12384 19116 12393
rect 21824 12427 21876 12436
rect 21824 12393 21833 12427
rect 21833 12393 21867 12427
rect 21867 12393 21876 12427
rect 21824 12384 21876 12393
rect 24032 12384 24084 12436
rect 10876 12316 10928 12368
rect 12164 12316 12216 12368
rect 12992 12316 13044 12368
rect 13912 12316 13964 12368
rect 9864 12248 9916 12300
rect 10968 12248 11020 12300
rect 13176 12248 13228 12300
rect 17316 12248 17368 12300
rect 19340 12248 19392 12300
rect 22100 12316 22152 12368
rect 22284 12291 22336 12300
rect 22284 12257 22318 12291
rect 22318 12257 22336 12291
rect 22284 12248 22336 12257
rect 24676 12248 24728 12300
rect 1860 12180 1912 12232
rect 5172 12180 5224 12232
rect 5540 12180 5592 12232
rect 6460 12180 6512 12232
rect 7012 12180 7064 12232
rect 7748 12180 7800 12232
rect 2504 12112 2556 12164
rect 4160 12112 4212 12164
rect 6000 12112 6052 12164
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 3240 12044 3292 12096
rect 3976 12044 4028 12096
rect 5172 12087 5224 12096
rect 5172 12053 5181 12087
rect 5181 12053 5215 12087
rect 5215 12053 5224 12087
rect 5172 12044 5224 12053
rect 6276 12087 6328 12096
rect 6276 12053 6285 12087
rect 6285 12053 6319 12087
rect 6319 12053 6328 12087
rect 6276 12044 6328 12053
rect 6644 12087 6696 12096
rect 6644 12053 6653 12087
rect 6653 12053 6687 12087
rect 6687 12053 6696 12087
rect 6644 12044 6696 12053
rect 7380 12044 7432 12096
rect 8116 12112 8168 12164
rect 8484 12180 8536 12232
rect 9496 12223 9548 12232
rect 9496 12189 9505 12223
rect 9505 12189 9539 12223
rect 9539 12189 9548 12223
rect 9496 12180 9548 12189
rect 10416 12223 10468 12232
rect 10416 12189 10425 12223
rect 10425 12189 10459 12223
rect 10459 12189 10468 12223
rect 10416 12180 10468 12189
rect 13912 12180 13964 12232
rect 16028 12180 16080 12232
rect 16580 12223 16632 12232
rect 16580 12189 16589 12223
rect 16589 12189 16623 12223
rect 16623 12189 16632 12223
rect 16580 12180 16632 12189
rect 19524 12223 19576 12232
rect 19524 12189 19533 12223
rect 19533 12189 19567 12223
rect 19567 12189 19576 12223
rect 19524 12180 19576 12189
rect 19616 12223 19668 12232
rect 19616 12189 19625 12223
rect 19625 12189 19659 12223
rect 19659 12189 19668 12223
rect 19616 12180 19668 12189
rect 21272 12180 21324 12232
rect 13452 12112 13504 12164
rect 8392 12044 8444 12096
rect 9496 12044 9548 12096
rect 10048 12044 10100 12096
rect 15568 12044 15620 12096
rect 17960 12087 18012 12096
rect 17960 12053 17969 12087
rect 17969 12053 18003 12087
rect 18003 12053 18012 12087
rect 17960 12044 18012 12053
rect 18972 12087 19024 12096
rect 18972 12053 18981 12087
rect 18981 12053 19015 12087
rect 19015 12053 19024 12087
rect 18972 12044 19024 12053
rect 19616 12044 19668 12096
rect 20996 12044 21048 12096
rect 24032 12087 24084 12096
rect 24032 12053 24041 12087
rect 24041 12053 24075 12087
rect 24075 12053 24084 12087
rect 24032 12044 24084 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2228 11883 2280 11892
rect 2228 11849 2237 11883
rect 2237 11849 2271 11883
rect 2271 11849 2280 11883
rect 2228 11840 2280 11849
rect 2320 11840 2372 11892
rect 2504 11840 2556 11892
rect 3332 11883 3384 11892
rect 3332 11849 3341 11883
rect 3341 11849 3375 11883
rect 3375 11849 3384 11883
rect 5172 11883 5224 11892
rect 3332 11840 3384 11849
rect 3148 11772 3200 11824
rect 5172 11849 5181 11883
rect 5181 11849 5215 11883
rect 5215 11849 5224 11883
rect 6460 11883 6512 11892
rect 5172 11840 5224 11849
rect 6460 11849 6469 11883
rect 6469 11849 6503 11883
rect 6503 11849 6512 11883
rect 6460 11840 6512 11849
rect 9036 11840 9088 11892
rect 9588 11840 9640 11892
rect 9772 11840 9824 11892
rect 13176 11883 13228 11892
rect 13176 11849 13185 11883
rect 13185 11849 13219 11883
rect 13219 11849 13228 11883
rect 13176 11840 13228 11849
rect 15660 11840 15712 11892
rect 17224 11840 17276 11892
rect 17316 11840 17368 11892
rect 22100 11840 22152 11892
rect 1952 11704 2004 11756
rect 2320 11568 2372 11620
rect 2688 11611 2740 11620
rect 2688 11577 2697 11611
rect 2697 11577 2731 11611
rect 2731 11577 2740 11611
rect 2688 11568 2740 11577
rect 2596 11543 2648 11552
rect 2596 11509 2605 11543
rect 2605 11509 2639 11543
rect 2639 11509 2648 11543
rect 2596 11500 2648 11509
rect 7104 11636 7156 11688
rect 7288 11679 7340 11688
rect 7288 11645 7297 11679
rect 7297 11645 7331 11679
rect 7331 11645 7340 11679
rect 7288 11636 7340 11645
rect 7564 11679 7616 11688
rect 7564 11645 7598 11679
rect 7598 11645 7616 11679
rect 10048 11772 10100 11824
rect 10968 11772 11020 11824
rect 15108 11772 15160 11824
rect 15936 11772 15988 11824
rect 18972 11772 19024 11824
rect 19248 11772 19300 11824
rect 21456 11772 21508 11824
rect 21640 11772 21692 11824
rect 8392 11704 8444 11756
rect 9588 11704 9640 11756
rect 7564 11636 7616 11645
rect 9036 11636 9088 11688
rect 10048 11636 10100 11688
rect 11428 11704 11480 11756
rect 14648 11704 14700 11756
rect 17960 11704 18012 11756
rect 20996 11704 21048 11756
rect 12624 11636 12676 11688
rect 13636 11679 13688 11688
rect 13636 11645 13645 11679
rect 13645 11645 13679 11679
rect 13679 11645 13688 11679
rect 13636 11636 13688 11645
rect 13912 11679 13964 11688
rect 13912 11645 13946 11679
rect 13946 11645 13964 11679
rect 13912 11636 13964 11645
rect 15568 11636 15620 11688
rect 19248 11636 19300 11688
rect 21364 11679 21416 11688
rect 21364 11645 21373 11679
rect 21373 11645 21407 11679
rect 21407 11645 21416 11679
rect 21364 11636 21416 11645
rect 22284 11636 22336 11688
rect 4068 11611 4120 11620
rect 4068 11577 4102 11611
rect 4102 11577 4120 11611
rect 4068 11568 4120 11577
rect 4252 11568 4304 11620
rect 5540 11568 5592 11620
rect 6552 11568 6604 11620
rect 7932 11568 7984 11620
rect 8852 11568 8904 11620
rect 10416 11568 10468 11620
rect 11152 11568 11204 11620
rect 14004 11568 14056 11620
rect 21088 11568 21140 11620
rect 24032 11568 24084 11620
rect 6000 11500 6052 11552
rect 6184 11543 6236 11552
rect 6184 11509 6193 11543
rect 6193 11509 6227 11543
rect 6227 11509 6236 11543
rect 6184 11500 6236 11509
rect 8300 11500 8352 11552
rect 9312 11543 9364 11552
rect 9312 11509 9321 11543
rect 9321 11509 9355 11543
rect 9355 11509 9364 11543
rect 9312 11500 9364 11509
rect 9496 11543 9548 11552
rect 9496 11509 9505 11543
rect 9505 11509 9539 11543
rect 9539 11509 9548 11543
rect 9496 11500 9548 11509
rect 9772 11543 9824 11552
rect 9772 11509 9781 11543
rect 9781 11509 9815 11543
rect 9815 11509 9824 11543
rect 9772 11500 9824 11509
rect 10876 11500 10928 11552
rect 11244 11543 11296 11552
rect 11244 11509 11253 11543
rect 11253 11509 11287 11543
rect 11287 11509 11296 11543
rect 11244 11500 11296 11509
rect 11796 11543 11848 11552
rect 11796 11509 11805 11543
rect 11805 11509 11839 11543
rect 11839 11509 11848 11543
rect 11796 11500 11848 11509
rect 12072 11500 12124 11552
rect 13452 11500 13504 11552
rect 15936 11543 15988 11552
rect 15936 11509 15945 11543
rect 15945 11509 15979 11543
rect 15979 11509 15988 11543
rect 15936 11500 15988 11509
rect 16580 11500 16632 11552
rect 17500 11500 17552 11552
rect 18052 11500 18104 11552
rect 18788 11543 18840 11552
rect 18788 11509 18797 11543
rect 18797 11509 18831 11543
rect 18831 11509 18840 11543
rect 18788 11500 18840 11509
rect 19248 11543 19300 11552
rect 19248 11509 19257 11543
rect 19257 11509 19291 11543
rect 19291 11509 19300 11543
rect 19248 11500 19300 11509
rect 20996 11500 21048 11552
rect 21732 11500 21784 11552
rect 21916 11500 21968 11552
rect 24860 11500 24912 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1492 11296 1544 11348
rect 2320 11339 2372 11348
rect 2320 11305 2329 11339
rect 2329 11305 2363 11339
rect 2363 11305 2372 11339
rect 2320 11296 2372 11305
rect 2412 11296 2464 11348
rect 2044 11228 2096 11280
rect 4344 11296 4396 11348
rect 6644 11296 6696 11348
rect 7012 11339 7064 11348
rect 7012 11305 7021 11339
rect 7021 11305 7055 11339
rect 7055 11305 7064 11339
rect 7012 11296 7064 11305
rect 7564 11296 7616 11348
rect 7656 11296 7708 11348
rect 9312 11296 9364 11348
rect 11244 11296 11296 11348
rect 12992 11339 13044 11348
rect 12992 11305 13001 11339
rect 13001 11305 13035 11339
rect 13035 11305 13044 11339
rect 12992 11296 13044 11305
rect 13176 11339 13228 11348
rect 13176 11305 13185 11339
rect 13185 11305 13219 11339
rect 13219 11305 13228 11339
rect 13176 11296 13228 11305
rect 14648 11339 14700 11348
rect 14648 11305 14657 11339
rect 14657 11305 14691 11339
rect 14691 11305 14700 11339
rect 14648 11296 14700 11305
rect 15108 11339 15160 11348
rect 15108 11305 15117 11339
rect 15117 11305 15151 11339
rect 15151 11305 15160 11339
rect 15108 11296 15160 11305
rect 17224 11339 17276 11348
rect 4528 11271 4580 11280
rect 4528 11237 4537 11271
rect 4537 11237 4571 11271
rect 4571 11237 4580 11271
rect 4528 11228 4580 11237
rect 6276 11228 6328 11280
rect 8116 11228 8168 11280
rect 9772 11228 9824 11280
rect 10692 11228 10744 11280
rect 11060 11228 11112 11280
rect 13084 11228 13136 11280
rect 13728 11228 13780 11280
rect 16580 11228 16632 11280
rect 17224 11305 17233 11339
rect 17233 11305 17267 11339
rect 17267 11305 17276 11339
rect 17224 11296 17276 11305
rect 18144 11296 18196 11348
rect 18788 11296 18840 11348
rect 21088 11296 21140 11348
rect 21732 11296 21784 11348
rect 22284 11339 22336 11348
rect 22284 11305 22293 11339
rect 22293 11305 22327 11339
rect 22327 11305 22336 11339
rect 22284 11296 22336 11305
rect 23848 11339 23900 11348
rect 23848 11305 23857 11339
rect 23857 11305 23891 11339
rect 23891 11305 23900 11339
rect 23848 11296 23900 11305
rect 25228 11339 25280 11348
rect 25228 11305 25237 11339
rect 25237 11305 25271 11339
rect 25271 11305 25280 11339
rect 25228 11296 25280 11305
rect 2320 11160 2372 11212
rect 2872 11160 2924 11212
rect 3056 11160 3108 11212
rect 3148 11160 3200 11212
rect 6460 11160 6512 11212
rect 9496 11160 9548 11212
rect 4620 11135 4672 11144
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 6092 11135 6144 11144
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6092 11092 6144 11101
rect 8668 11135 8720 11144
rect 2872 11024 2924 11076
rect 4068 11024 4120 11076
rect 6000 11024 6052 11076
rect 8668 11101 8677 11135
rect 8677 11101 8711 11135
rect 8711 11101 8720 11135
rect 8668 11092 8720 11101
rect 11244 11160 11296 11212
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 13912 11092 13964 11144
rect 14004 11092 14056 11144
rect 15292 11135 15344 11144
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 17500 11092 17552 11144
rect 19248 11228 19300 11280
rect 19064 11160 19116 11212
rect 22100 11228 22152 11280
rect 22836 11228 22888 11280
rect 24676 11228 24728 11280
rect 24952 11228 25004 11280
rect 20996 11160 21048 11212
rect 22284 11160 22336 11212
rect 25044 11203 25096 11212
rect 25044 11169 25053 11203
rect 25053 11169 25087 11203
rect 25087 11169 25096 11203
rect 25044 11160 25096 11169
rect 24032 11135 24084 11144
rect 24032 11101 24041 11135
rect 24041 11101 24075 11135
rect 24075 11101 24084 11135
rect 24584 11135 24636 11144
rect 24032 11092 24084 11101
rect 24584 11101 24593 11135
rect 24593 11101 24627 11135
rect 24627 11101 24636 11135
rect 24584 11092 24636 11101
rect 9588 11024 9640 11076
rect 3608 10956 3660 11008
rect 5172 10999 5224 11008
rect 5172 10965 5181 10999
rect 5181 10965 5215 10999
rect 5215 10965 5224 10999
rect 5172 10956 5224 10965
rect 5448 10956 5500 11008
rect 6092 10956 6144 11008
rect 8944 10956 8996 11008
rect 10048 11024 10100 11076
rect 10232 11067 10284 11076
rect 10232 11033 10241 11067
rect 10241 11033 10275 11067
rect 10275 11033 10284 11067
rect 10232 11024 10284 11033
rect 20720 11024 20772 11076
rect 10692 10956 10744 11008
rect 17960 10999 18012 11008
rect 17960 10965 17969 10999
rect 17969 10965 18003 10999
rect 18003 10965 18012 10999
rect 17960 10956 18012 10965
rect 20076 10956 20128 11008
rect 22468 11024 22520 11076
rect 22100 10956 22152 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2964 10752 3016 10804
rect 4620 10795 4672 10804
rect 4620 10761 4629 10795
rect 4629 10761 4663 10795
rect 4663 10761 4672 10795
rect 4620 10752 4672 10761
rect 6460 10795 6512 10804
rect 6460 10761 6469 10795
rect 6469 10761 6503 10795
rect 6503 10761 6512 10795
rect 6460 10752 6512 10761
rect 8484 10752 8536 10804
rect 8944 10795 8996 10804
rect 8944 10761 8953 10795
rect 8953 10761 8987 10795
rect 8987 10761 8996 10795
rect 8944 10752 8996 10761
rect 13636 10752 13688 10804
rect 13912 10752 13964 10804
rect 16856 10795 16908 10804
rect 16856 10761 16865 10795
rect 16865 10761 16899 10795
rect 16899 10761 16908 10795
rect 16856 10752 16908 10761
rect 18880 10752 18932 10804
rect 20628 10795 20680 10804
rect 20628 10761 20637 10795
rect 20637 10761 20671 10795
rect 20671 10761 20680 10795
rect 20628 10752 20680 10761
rect 23296 10752 23348 10804
rect 24676 10795 24728 10804
rect 24676 10761 24685 10795
rect 24685 10761 24719 10795
rect 24719 10761 24728 10795
rect 24676 10752 24728 10761
rect 25044 10795 25096 10804
rect 25044 10761 25053 10795
rect 25053 10761 25087 10795
rect 25087 10761 25096 10795
rect 25044 10752 25096 10761
rect 25504 10752 25556 10804
rect 11796 10684 11848 10736
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 6000 10616 6052 10668
rect 3332 10548 3384 10600
rect 3608 10548 3660 10600
rect 5540 10548 5592 10600
rect 7288 10548 7340 10600
rect 7656 10548 7708 10600
rect 2872 10523 2924 10532
rect 2872 10489 2906 10523
rect 2906 10489 2924 10523
rect 2872 10480 2924 10489
rect 2964 10480 3016 10532
rect 3884 10480 3936 10532
rect 2320 10455 2372 10464
rect 2320 10421 2329 10455
rect 2329 10421 2363 10455
rect 2363 10421 2372 10455
rect 2320 10412 2372 10421
rect 8208 10548 8260 10600
rect 9680 10548 9732 10600
rect 11704 10616 11756 10668
rect 12072 10616 12124 10668
rect 18788 10659 18840 10668
rect 18788 10625 18797 10659
rect 18797 10625 18831 10659
rect 18831 10625 18840 10659
rect 18788 10616 18840 10625
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 21364 10616 21416 10668
rect 24308 10659 24360 10668
rect 24308 10625 24317 10659
rect 24317 10625 24351 10659
rect 24351 10625 24360 10659
rect 24308 10616 24360 10625
rect 24860 10616 24912 10668
rect 10968 10548 11020 10600
rect 12624 10548 12676 10600
rect 13084 10548 13136 10600
rect 15292 10548 15344 10600
rect 13728 10480 13780 10532
rect 14556 10480 14608 10532
rect 5172 10412 5224 10464
rect 6184 10455 6236 10464
rect 6184 10421 6193 10455
rect 6193 10421 6227 10455
rect 6227 10421 6236 10455
rect 6184 10412 6236 10421
rect 7656 10412 7708 10464
rect 9588 10455 9640 10464
rect 9588 10421 9597 10455
rect 9597 10421 9631 10455
rect 9631 10421 9640 10455
rect 9588 10412 9640 10421
rect 9772 10412 9824 10464
rect 10692 10412 10744 10464
rect 11244 10412 11296 10464
rect 13636 10412 13688 10464
rect 14464 10455 14516 10464
rect 14464 10421 14473 10455
rect 14473 10421 14507 10455
rect 14507 10421 14516 10455
rect 14464 10412 14516 10421
rect 15568 10548 15620 10600
rect 16488 10548 16540 10600
rect 20720 10548 20772 10600
rect 22468 10591 22520 10600
rect 22468 10557 22477 10591
rect 22477 10557 22511 10591
rect 22511 10557 22520 10591
rect 22468 10548 22520 10557
rect 23112 10548 23164 10600
rect 25228 10591 25280 10600
rect 25228 10557 25237 10591
rect 25237 10557 25271 10591
rect 25271 10557 25280 10591
rect 25228 10548 25280 10557
rect 17960 10480 18012 10532
rect 22284 10480 22336 10532
rect 23756 10480 23808 10532
rect 24124 10523 24176 10532
rect 24124 10489 24133 10523
rect 24133 10489 24167 10523
rect 24167 10489 24176 10523
rect 24124 10480 24176 10489
rect 17500 10412 17552 10464
rect 18696 10455 18748 10464
rect 18696 10421 18705 10455
rect 18705 10421 18739 10455
rect 18739 10421 18748 10455
rect 18696 10412 18748 10421
rect 19064 10412 19116 10464
rect 19432 10412 19484 10464
rect 20352 10412 20404 10464
rect 22560 10412 22612 10464
rect 23664 10455 23716 10464
rect 23664 10421 23673 10455
rect 23673 10421 23707 10455
rect 23707 10421 23716 10455
rect 23664 10412 23716 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2412 10251 2464 10260
rect 2412 10217 2421 10251
rect 2421 10217 2455 10251
rect 2455 10217 2464 10251
rect 2412 10208 2464 10217
rect 7564 10251 7616 10260
rect 7564 10217 7573 10251
rect 7573 10217 7607 10251
rect 7607 10217 7616 10251
rect 7564 10208 7616 10217
rect 8668 10251 8720 10260
rect 8668 10217 8677 10251
rect 8677 10217 8711 10251
rect 8711 10217 8720 10251
rect 8668 10208 8720 10217
rect 9312 10251 9364 10260
rect 9312 10217 9321 10251
rect 9321 10217 9355 10251
rect 9355 10217 9364 10251
rect 9312 10208 9364 10217
rect 11152 10251 11204 10260
rect 11152 10217 11161 10251
rect 11161 10217 11195 10251
rect 11195 10217 11204 10251
rect 11152 10208 11204 10217
rect 11796 10208 11848 10260
rect 14464 10251 14516 10260
rect 14464 10217 14473 10251
rect 14473 10217 14507 10251
rect 14507 10217 14516 10251
rect 14464 10208 14516 10217
rect 15568 10208 15620 10260
rect 17960 10208 18012 10260
rect 20444 10208 20496 10260
rect 20720 10208 20772 10260
rect 21272 10251 21324 10260
rect 21272 10217 21281 10251
rect 21281 10217 21315 10251
rect 21315 10217 21324 10251
rect 21272 10208 21324 10217
rect 21364 10251 21416 10260
rect 21364 10217 21373 10251
rect 21373 10217 21407 10251
rect 21407 10217 21416 10251
rect 21364 10208 21416 10217
rect 21916 10208 21968 10260
rect 22100 10251 22152 10260
rect 22100 10217 22109 10251
rect 22109 10217 22143 10251
rect 22143 10217 22152 10251
rect 23112 10251 23164 10260
rect 22100 10208 22152 10217
rect 23112 10217 23121 10251
rect 23121 10217 23155 10251
rect 23155 10217 23164 10251
rect 23112 10208 23164 10217
rect 2872 10140 2924 10192
rect 2780 10115 2832 10124
rect 2780 10081 2789 10115
rect 2789 10081 2823 10115
rect 2823 10081 2832 10115
rect 2780 10072 2832 10081
rect 2964 10004 3016 10056
rect 3332 10072 3384 10124
rect 5356 10140 5408 10192
rect 6184 10140 6236 10192
rect 8944 10183 8996 10192
rect 6000 10072 6052 10124
rect 7564 10072 7616 10124
rect 8944 10149 8953 10183
rect 8953 10149 8987 10183
rect 8987 10149 8996 10183
rect 8944 10140 8996 10149
rect 9864 10140 9916 10192
rect 15292 10140 15344 10192
rect 18052 10183 18104 10192
rect 18052 10149 18061 10183
rect 18061 10149 18095 10183
rect 18095 10149 18104 10183
rect 18052 10140 18104 10149
rect 23664 10140 23716 10192
rect 8392 10072 8444 10124
rect 11060 10115 11112 10124
rect 11060 10081 11069 10115
rect 11069 10081 11103 10115
rect 11103 10081 11112 10115
rect 11060 10072 11112 10081
rect 12348 10072 12400 10124
rect 8208 10047 8260 10056
rect 1492 9936 1544 9988
rect 2596 9936 2648 9988
rect 1768 9868 1820 9920
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 11612 10004 11664 10056
rect 7748 9936 7800 9988
rect 12900 10072 12952 10124
rect 13084 10115 13136 10124
rect 13084 10081 13093 10115
rect 13093 10081 13127 10115
rect 13127 10081 13136 10115
rect 13084 10072 13136 10081
rect 15936 10072 15988 10124
rect 17776 10072 17828 10124
rect 19340 10072 19392 10124
rect 19892 10072 19944 10124
rect 22560 10072 22612 10124
rect 23112 10072 23164 10124
rect 24308 10072 24360 10124
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 15384 10004 15436 10056
rect 16672 10047 16724 10056
rect 16672 10013 16681 10047
rect 16681 10013 16715 10047
rect 16715 10013 16724 10047
rect 16672 10004 16724 10013
rect 18144 10004 18196 10056
rect 14832 9936 14884 9988
rect 19432 9936 19484 9988
rect 19984 9979 20036 9988
rect 19984 9945 19993 9979
rect 19993 9945 20027 9979
rect 20027 9945 20036 9979
rect 19984 9936 20036 9945
rect 20352 9936 20404 9988
rect 20996 9936 21048 9988
rect 22284 10004 22336 10056
rect 22836 10004 22888 10056
rect 5172 9868 5224 9920
rect 6000 9868 6052 9920
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 6920 9868 6972 9877
rect 9864 9868 9916 9920
rect 10692 9911 10744 9920
rect 10692 9877 10701 9911
rect 10701 9877 10735 9911
rect 10735 9877 10744 9911
rect 10692 9868 10744 9877
rect 12624 9868 12676 9920
rect 12992 9868 13044 9920
rect 13912 9868 13964 9920
rect 14004 9868 14056 9920
rect 16396 9911 16448 9920
rect 16396 9877 16405 9911
rect 16405 9877 16439 9911
rect 16439 9877 16448 9911
rect 16396 9868 16448 9877
rect 17592 9911 17644 9920
rect 17592 9877 17601 9911
rect 17601 9877 17635 9911
rect 17635 9877 17644 9911
rect 17592 9868 17644 9877
rect 24768 9868 24820 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 8668 9664 8720 9716
rect 10600 9664 10652 9716
rect 10876 9664 10928 9716
rect 13268 9664 13320 9716
rect 19432 9707 19484 9716
rect 19432 9673 19441 9707
rect 19441 9673 19475 9707
rect 19475 9673 19484 9707
rect 19432 9664 19484 9673
rect 19892 9664 19944 9716
rect 20352 9707 20404 9716
rect 20352 9673 20361 9707
rect 20361 9673 20395 9707
rect 20395 9673 20404 9707
rect 20352 9664 20404 9673
rect 21272 9664 21324 9716
rect 22008 9664 22060 9716
rect 22652 9664 22704 9716
rect 22836 9664 22888 9716
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 2596 9596 2648 9648
rect 4068 9596 4120 9648
rect 4344 9639 4396 9648
rect 4344 9605 4353 9639
rect 4353 9605 4387 9639
rect 4387 9605 4396 9639
rect 4344 9596 4396 9605
rect 11152 9596 11204 9648
rect 12164 9639 12216 9648
rect 12164 9605 12173 9639
rect 12173 9605 12207 9639
rect 12207 9605 12216 9639
rect 12164 9596 12216 9605
rect 12440 9639 12492 9648
rect 12440 9605 12449 9639
rect 12449 9605 12483 9639
rect 12483 9605 12492 9639
rect 12440 9596 12492 9605
rect 12900 9596 12952 9648
rect 14280 9639 14332 9648
rect 14280 9605 14289 9639
rect 14289 9605 14323 9639
rect 14323 9605 14332 9639
rect 14280 9596 14332 9605
rect 17132 9639 17184 9648
rect 1584 9460 1636 9512
rect 1860 9392 1912 9444
rect 1308 9324 1360 9376
rect 2964 9392 3016 9444
rect 5172 9528 5224 9580
rect 5448 9460 5500 9512
rect 7656 9460 7708 9512
rect 10692 9528 10744 9580
rect 10876 9528 10928 9580
rect 17132 9605 17141 9639
rect 17141 9605 17175 9639
rect 17175 9605 17184 9639
rect 17132 9596 17184 9605
rect 17500 9639 17552 9648
rect 17500 9605 17509 9639
rect 17509 9605 17543 9639
rect 17543 9605 17552 9639
rect 17500 9596 17552 9605
rect 17776 9639 17828 9648
rect 17776 9605 17785 9639
rect 17785 9605 17819 9639
rect 17819 9605 17828 9639
rect 17776 9596 17828 9605
rect 21824 9596 21876 9648
rect 22100 9596 22152 9648
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 13268 9528 13320 9580
rect 15016 9571 15068 9580
rect 15016 9537 15025 9571
rect 15025 9537 15059 9571
rect 15059 9537 15068 9571
rect 15016 9528 15068 9537
rect 16672 9571 16724 9580
rect 16672 9537 16681 9571
rect 16681 9537 16715 9571
rect 16715 9537 16724 9571
rect 16672 9528 16724 9537
rect 8484 9460 8536 9512
rect 12440 9460 12492 9512
rect 12900 9503 12952 9512
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 21364 9528 21416 9580
rect 23480 9596 23532 9648
rect 25412 9639 25464 9648
rect 25412 9605 25421 9639
rect 25421 9605 25455 9639
rect 25455 9605 25464 9639
rect 25412 9596 25464 9605
rect 23112 9528 23164 9580
rect 14464 9460 14516 9512
rect 15936 9460 15988 9512
rect 17776 9460 17828 9512
rect 20444 9460 20496 9512
rect 21916 9503 21968 9512
rect 21916 9469 21925 9503
rect 21925 9469 21959 9503
rect 21959 9469 21968 9503
rect 21916 9460 21968 9469
rect 23664 9460 23716 9512
rect 24768 9460 24820 9512
rect 25228 9503 25280 9512
rect 25228 9469 25237 9503
rect 25237 9469 25271 9503
rect 25271 9469 25280 9503
rect 25228 9460 25280 9469
rect 8576 9392 8628 9444
rect 3424 9324 3476 9376
rect 5356 9367 5408 9376
rect 5356 9333 5365 9367
rect 5365 9333 5399 9367
rect 5399 9333 5408 9367
rect 5356 9324 5408 9333
rect 5448 9324 5500 9376
rect 6000 9324 6052 9376
rect 6276 9324 6328 9376
rect 7564 9367 7616 9376
rect 7564 9333 7573 9367
rect 7573 9333 7607 9367
rect 7607 9333 7616 9367
rect 7564 9324 7616 9333
rect 9220 9324 9272 9376
rect 13268 9392 13320 9444
rect 14280 9392 14332 9444
rect 16120 9392 16172 9444
rect 17960 9392 18012 9444
rect 10140 9324 10192 9376
rect 11612 9367 11664 9376
rect 11612 9333 11621 9367
rect 11621 9333 11655 9367
rect 11655 9333 11664 9367
rect 11612 9324 11664 9333
rect 14464 9367 14516 9376
rect 14464 9333 14473 9367
rect 14473 9333 14507 9367
rect 14507 9333 14516 9367
rect 14464 9324 14516 9333
rect 15844 9367 15896 9376
rect 15844 9333 15853 9367
rect 15853 9333 15887 9367
rect 15887 9333 15896 9367
rect 15844 9324 15896 9333
rect 16028 9367 16080 9376
rect 16028 9333 16037 9367
rect 16037 9333 16071 9367
rect 16071 9333 16080 9367
rect 16028 9324 16080 9333
rect 16396 9367 16448 9376
rect 16396 9333 16405 9367
rect 16405 9333 16439 9367
rect 16439 9333 16448 9367
rect 16396 9324 16448 9333
rect 24860 9324 24912 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 2228 9120 2280 9172
rect 4068 9120 4120 9172
rect 7196 9163 7248 9172
rect 7196 9129 7205 9163
rect 7205 9129 7239 9163
rect 7239 9129 7248 9163
rect 7196 9120 7248 9129
rect 8668 9120 8720 9172
rect 11060 9120 11112 9172
rect 12440 9163 12492 9172
rect 12440 9129 12449 9163
rect 12449 9129 12483 9163
rect 12483 9129 12492 9163
rect 15016 9163 15068 9172
rect 12440 9120 12492 9129
rect 15016 9129 15025 9163
rect 15025 9129 15059 9163
rect 15059 9129 15068 9163
rect 15016 9120 15068 9129
rect 15384 9120 15436 9172
rect 17592 9163 17644 9172
rect 17592 9129 17601 9163
rect 17601 9129 17635 9163
rect 17635 9129 17644 9163
rect 17592 9120 17644 9129
rect 18696 9120 18748 9172
rect 20260 9163 20312 9172
rect 20260 9129 20269 9163
rect 20269 9129 20303 9163
rect 20303 9129 20312 9163
rect 20260 9120 20312 9129
rect 20352 9120 20404 9172
rect 21180 9120 21232 9172
rect 21364 9163 21416 9172
rect 21364 9129 21373 9163
rect 21373 9129 21407 9163
rect 21407 9129 21416 9163
rect 21364 9120 21416 9129
rect 23112 9120 23164 9172
rect 2872 9052 2924 9104
rect 6184 9052 6236 9104
rect 15660 9052 15712 9104
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 1860 8984 1912 9036
rect 4344 9027 4396 9036
rect 4344 8993 4378 9027
rect 4378 8993 4396 9027
rect 4344 8984 4396 8993
rect 8024 8984 8076 9036
rect 8392 8984 8444 9036
rect 2596 8916 2648 8968
rect 2964 8959 3016 8968
rect 2964 8925 2973 8959
rect 2973 8925 3007 8959
rect 3007 8925 3016 8959
rect 4068 8959 4120 8968
rect 2964 8916 3016 8925
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 7748 8959 7800 8968
rect 7748 8925 7757 8959
rect 7757 8925 7791 8959
rect 7791 8925 7800 8959
rect 7748 8916 7800 8925
rect 9588 8984 9640 9036
rect 10508 9027 10560 9036
rect 10508 8993 10542 9027
rect 10542 8993 10560 9027
rect 10508 8984 10560 8993
rect 12992 9027 13044 9036
rect 12992 8993 13026 9027
rect 13026 8993 13044 9027
rect 12992 8984 13044 8993
rect 14740 8984 14792 9036
rect 18052 8984 18104 9036
rect 18236 8984 18288 9036
rect 8576 8916 8628 8968
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 12440 8916 12492 8968
rect 20628 9052 20680 9104
rect 24768 9052 24820 9104
rect 20536 8984 20588 9036
rect 22836 8984 22888 9036
rect 23756 9027 23808 9036
rect 23756 8993 23765 9027
rect 23765 8993 23799 9027
rect 23799 8993 23808 9027
rect 23756 8984 23808 8993
rect 1952 8823 2004 8832
rect 1952 8789 1961 8823
rect 1961 8789 1995 8823
rect 1995 8789 2004 8823
rect 1952 8780 2004 8789
rect 3332 8780 3384 8832
rect 3884 8823 3936 8832
rect 3884 8789 3893 8823
rect 3893 8789 3927 8823
rect 3927 8789 3936 8823
rect 3884 8780 3936 8789
rect 8300 8848 8352 8900
rect 15108 8848 15160 8900
rect 17500 8848 17552 8900
rect 20904 8916 20956 8968
rect 5448 8823 5500 8832
rect 5448 8789 5457 8823
rect 5457 8789 5491 8823
rect 5491 8789 5500 8823
rect 5448 8780 5500 8789
rect 6000 8823 6052 8832
rect 6000 8789 6009 8823
rect 6009 8789 6043 8823
rect 6043 8789 6052 8823
rect 6000 8780 6052 8789
rect 6368 8823 6420 8832
rect 6368 8789 6377 8823
rect 6377 8789 6411 8823
rect 6411 8789 6420 8823
rect 6368 8780 6420 8789
rect 7104 8823 7156 8832
rect 7104 8789 7113 8823
rect 7113 8789 7147 8823
rect 7147 8789 7156 8823
rect 7104 8780 7156 8789
rect 7196 8780 7248 8832
rect 9404 8780 9456 8832
rect 9864 8823 9916 8832
rect 9864 8789 9873 8823
rect 9873 8789 9907 8823
rect 9907 8789 9916 8823
rect 9864 8780 9916 8789
rect 10416 8780 10468 8832
rect 10968 8780 11020 8832
rect 14096 8823 14148 8832
rect 14096 8789 14105 8823
rect 14105 8789 14139 8823
rect 14139 8789 14148 8823
rect 14096 8780 14148 8789
rect 17960 8823 18012 8832
rect 17960 8789 17969 8823
rect 17969 8789 18003 8823
rect 18003 8789 18012 8823
rect 17960 8780 18012 8789
rect 21272 8848 21324 8900
rect 23204 8916 23256 8968
rect 18604 8780 18656 8832
rect 19064 8823 19116 8832
rect 19064 8789 19073 8823
rect 19073 8789 19107 8823
rect 19107 8789 19116 8823
rect 19064 8780 19116 8789
rect 19432 8823 19484 8832
rect 19432 8789 19441 8823
rect 19441 8789 19475 8823
rect 19475 8789 19484 8823
rect 19432 8780 19484 8789
rect 20444 8780 20496 8832
rect 20720 8780 20772 8832
rect 21364 8780 21416 8832
rect 21732 8780 21784 8832
rect 25136 8823 25188 8832
rect 25136 8789 25145 8823
rect 25145 8789 25179 8823
rect 25179 8789 25188 8823
rect 25136 8780 25188 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2596 8576 2648 8628
rect 4620 8576 4672 8628
rect 5264 8576 5316 8628
rect 7196 8619 7248 8628
rect 7196 8585 7205 8619
rect 7205 8585 7239 8619
rect 7239 8585 7248 8619
rect 7196 8576 7248 8585
rect 4068 8508 4120 8560
rect 5356 8508 5408 8560
rect 5540 8508 5592 8560
rect 7288 8508 7340 8560
rect 7472 8508 7524 8560
rect 2228 8415 2280 8424
rect 2228 8381 2237 8415
rect 2237 8381 2271 8415
rect 2271 8381 2280 8415
rect 2228 8372 2280 8381
rect 5448 8440 5500 8492
rect 7104 8440 7156 8492
rect 10508 8576 10560 8628
rect 10692 8576 10744 8628
rect 14188 8576 14240 8628
rect 16672 8576 16724 8628
rect 17500 8619 17552 8628
rect 17500 8585 17509 8619
rect 17509 8585 17543 8619
rect 17543 8585 17552 8619
rect 17500 8576 17552 8585
rect 17960 8576 18012 8628
rect 20352 8576 20404 8628
rect 20628 8576 20680 8628
rect 24860 8619 24912 8628
rect 24860 8585 24869 8619
rect 24869 8585 24903 8619
rect 24903 8585 24912 8619
rect 24860 8576 24912 8585
rect 25136 8576 25188 8628
rect 25596 8619 25648 8628
rect 25596 8585 25605 8619
rect 25605 8585 25639 8619
rect 25639 8585 25648 8619
rect 25596 8576 25648 8585
rect 8576 8551 8628 8560
rect 8576 8517 8585 8551
rect 8585 8517 8619 8551
rect 8619 8517 8628 8551
rect 8576 8508 8628 8517
rect 8024 8440 8076 8492
rect 2872 8372 2924 8424
rect 3056 8372 3108 8424
rect 5356 8372 5408 8424
rect 8576 8372 8628 8424
rect 10232 8440 10284 8492
rect 11060 8440 11112 8492
rect 11244 8440 11296 8492
rect 11612 8440 11664 8492
rect 9312 8372 9364 8424
rect 12440 8415 12492 8424
rect 12440 8381 12449 8415
rect 12449 8381 12483 8415
rect 12483 8381 12492 8415
rect 12440 8372 12492 8381
rect 14096 8372 14148 8424
rect 1952 8304 2004 8356
rect 2504 8347 2556 8356
rect 2504 8313 2516 8347
rect 2516 8313 2556 8347
rect 2504 8304 2556 8313
rect 2596 8236 2648 8288
rect 4344 8304 4396 8356
rect 6184 8304 6236 8356
rect 5448 8236 5500 8288
rect 8668 8304 8720 8356
rect 12900 8304 12952 8356
rect 14740 8372 14792 8424
rect 15016 8415 15068 8424
rect 15016 8381 15025 8415
rect 15025 8381 15059 8415
rect 15059 8381 15068 8415
rect 15016 8372 15068 8381
rect 15108 8372 15160 8424
rect 15568 8372 15620 8424
rect 16304 8508 16356 8560
rect 18052 8508 18104 8560
rect 21732 8508 21784 8560
rect 24492 8483 24544 8492
rect 24492 8449 24501 8483
rect 24501 8449 24535 8483
rect 24535 8449 24544 8483
rect 24492 8440 24544 8449
rect 17776 8372 17828 8424
rect 20628 8415 20680 8424
rect 20628 8381 20637 8415
rect 20637 8381 20671 8415
rect 20671 8381 20680 8415
rect 20628 8372 20680 8381
rect 24676 8372 24728 8424
rect 25412 8415 25464 8424
rect 25412 8381 25421 8415
rect 25421 8381 25455 8415
rect 25455 8381 25464 8415
rect 25412 8372 25464 8381
rect 7564 8279 7616 8288
rect 7564 8245 7573 8279
rect 7573 8245 7607 8279
rect 7607 8245 7616 8279
rect 7564 8236 7616 8245
rect 11244 8279 11296 8288
rect 11244 8245 11253 8279
rect 11253 8245 11287 8279
rect 11287 8245 11296 8279
rect 11244 8236 11296 8245
rect 12716 8236 12768 8288
rect 15384 8304 15436 8356
rect 16764 8304 16816 8356
rect 19248 8304 19300 8356
rect 20904 8347 20956 8356
rect 20904 8313 20916 8347
rect 20916 8313 20956 8347
rect 23480 8347 23532 8356
rect 20904 8304 20956 8313
rect 15660 8236 15712 8288
rect 20352 8236 20404 8288
rect 23480 8313 23489 8347
rect 23489 8313 23523 8347
rect 23523 8313 23532 8347
rect 23480 8304 23532 8313
rect 22284 8236 22336 8288
rect 22560 8279 22612 8288
rect 22560 8245 22569 8279
rect 22569 8245 22603 8279
rect 22603 8245 22612 8279
rect 22560 8236 22612 8245
rect 23848 8279 23900 8288
rect 23848 8245 23857 8279
rect 23857 8245 23891 8279
rect 23891 8245 23900 8279
rect 23848 8236 23900 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2136 8032 2188 8084
rect 2504 8032 2556 8084
rect 5356 8032 5408 8084
rect 7748 8032 7800 8084
rect 9220 8032 9272 8084
rect 9588 8032 9640 8084
rect 9680 8032 9732 8084
rect 11244 8032 11296 8084
rect 12164 8032 12216 8084
rect 12900 8032 12952 8084
rect 12992 8032 13044 8084
rect 13544 8032 13596 8084
rect 14464 8032 14516 8084
rect 1676 7964 1728 8016
rect 2228 8007 2280 8016
rect 2228 7973 2237 8007
rect 2237 7973 2271 8007
rect 2271 7973 2280 8007
rect 2228 7964 2280 7973
rect 2412 7964 2464 8016
rect 2688 8007 2740 8016
rect 2688 7973 2697 8007
rect 2697 7973 2731 8007
rect 2731 7973 2740 8007
rect 2688 7964 2740 7973
rect 8668 7964 8720 8016
rect 11612 8007 11664 8016
rect 11612 7973 11621 8007
rect 11621 7973 11655 8007
rect 11655 7973 11664 8007
rect 11612 7964 11664 7973
rect 12348 7964 12400 8016
rect 14832 8032 14884 8084
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 17408 8032 17460 8084
rect 17868 8032 17920 8084
rect 18052 8075 18104 8084
rect 18052 8041 18061 8075
rect 18061 8041 18095 8075
rect 18095 8041 18104 8075
rect 18052 8032 18104 8041
rect 19064 8032 19116 8084
rect 19248 8032 19300 8084
rect 20628 8032 20680 8084
rect 22284 8075 22336 8084
rect 22284 8041 22293 8075
rect 22293 8041 22327 8075
rect 22327 8041 22336 8075
rect 22284 8032 22336 8041
rect 22744 8032 22796 8084
rect 23756 8075 23808 8084
rect 23756 8041 23765 8075
rect 23765 8041 23799 8075
rect 23799 8041 23808 8075
rect 23756 8032 23808 8041
rect 15016 7964 15068 8016
rect 17776 7964 17828 8016
rect 20536 7964 20588 8016
rect 21272 7964 21324 8016
rect 3608 7896 3660 7948
rect 6092 7896 6144 7948
rect 8944 7896 8996 7948
rect 10508 7939 10560 7948
rect 10508 7905 10517 7939
rect 10517 7905 10551 7939
rect 10551 7905 10560 7939
rect 10508 7896 10560 7905
rect 1676 7828 1728 7880
rect 2596 7828 2648 7880
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 5540 7871 5592 7880
rect 5540 7837 5549 7871
rect 5549 7837 5583 7871
rect 5583 7837 5592 7871
rect 5540 7828 5592 7837
rect 8852 7828 8904 7880
rect 9128 7828 9180 7880
rect 9496 7828 9548 7880
rect 10600 7871 10652 7880
rect 10600 7837 10609 7871
rect 10609 7837 10643 7871
rect 10643 7837 10652 7871
rect 10600 7828 10652 7837
rect 10692 7871 10744 7880
rect 10692 7837 10701 7871
rect 10701 7837 10735 7871
rect 10735 7837 10744 7871
rect 10692 7828 10744 7837
rect 11796 7828 11848 7880
rect 15568 7896 15620 7948
rect 15844 7896 15896 7948
rect 17960 7896 18012 7948
rect 16764 7871 16816 7880
rect 2964 7760 3016 7812
rect 7288 7760 7340 7812
rect 7932 7760 7984 7812
rect 10876 7760 10928 7812
rect 16764 7837 16773 7871
rect 16773 7837 16807 7871
rect 16807 7837 16816 7871
rect 16764 7828 16816 7837
rect 19984 7896 20036 7948
rect 24492 7964 24544 8016
rect 19800 7871 19852 7880
rect 12716 7760 12768 7812
rect 15568 7760 15620 7812
rect 19800 7837 19809 7871
rect 19809 7837 19843 7871
rect 19843 7837 19852 7871
rect 19800 7828 19852 7837
rect 20352 7828 20404 7880
rect 20904 7871 20956 7880
rect 20904 7837 20913 7871
rect 20913 7837 20947 7871
rect 20947 7837 20956 7871
rect 20904 7828 20956 7837
rect 18512 7760 18564 7812
rect 1400 7692 1452 7744
rect 2872 7692 2924 7744
rect 4528 7735 4580 7744
rect 4528 7701 4537 7735
rect 4537 7701 4571 7735
rect 4571 7701 4580 7735
rect 4528 7692 4580 7701
rect 6920 7735 6972 7744
rect 6920 7701 6929 7735
rect 6929 7701 6963 7735
rect 6963 7701 6972 7735
rect 6920 7692 6972 7701
rect 7564 7735 7616 7744
rect 7564 7701 7573 7735
rect 7573 7701 7607 7735
rect 7607 7701 7616 7735
rect 7564 7692 7616 7701
rect 8024 7735 8076 7744
rect 8024 7701 8033 7735
rect 8033 7701 8067 7735
rect 8067 7701 8076 7735
rect 8024 7692 8076 7701
rect 9036 7735 9088 7744
rect 9036 7701 9045 7735
rect 9045 7701 9079 7735
rect 9079 7701 9088 7735
rect 9036 7692 9088 7701
rect 9128 7692 9180 7744
rect 10048 7735 10100 7744
rect 10048 7701 10057 7735
rect 10057 7701 10091 7735
rect 10091 7701 10100 7735
rect 10048 7692 10100 7701
rect 11244 7735 11296 7744
rect 11244 7701 11253 7735
rect 11253 7701 11287 7735
rect 11287 7701 11296 7735
rect 11244 7692 11296 7701
rect 11704 7735 11756 7744
rect 11704 7701 11713 7735
rect 11713 7701 11747 7735
rect 11747 7701 11756 7735
rect 11704 7692 11756 7701
rect 15660 7692 15712 7744
rect 16856 7692 16908 7744
rect 16948 7692 17000 7744
rect 24676 7692 24728 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1676 7531 1728 7540
rect 1676 7497 1685 7531
rect 1685 7497 1719 7531
rect 1719 7497 1728 7531
rect 1676 7488 1728 7497
rect 3516 7531 3568 7540
rect 3516 7497 3525 7531
rect 3525 7497 3559 7531
rect 3559 7497 3568 7531
rect 3516 7488 3568 7497
rect 5172 7531 5224 7540
rect 5172 7497 5181 7531
rect 5181 7497 5215 7531
rect 5215 7497 5224 7531
rect 5172 7488 5224 7497
rect 6092 7488 6144 7540
rect 10784 7531 10836 7540
rect 10784 7497 10793 7531
rect 10793 7497 10827 7531
rect 10827 7497 10836 7531
rect 10784 7488 10836 7497
rect 11796 7531 11848 7540
rect 11796 7497 11805 7531
rect 11805 7497 11839 7531
rect 11839 7497 11848 7531
rect 11796 7488 11848 7497
rect 12164 7531 12216 7540
rect 12164 7497 12173 7531
rect 12173 7497 12207 7531
rect 12207 7497 12216 7531
rect 12164 7488 12216 7497
rect 12716 7531 12768 7540
rect 12716 7497 12725 7531
rect 12725 7497 12759 7531
rect 12759 7497 12768 7531
rect 12716 7488 12768 7497
rect 12900 7488 12952 7540
rect 4436 7395 4488 7404
rect 4436 7361 4445 7395
rect 4445 7361 4479 7395
rect 4479 7361 4488 7395
rect 4436 7352 4488 7361
rect 5632 7352 5684 7404
rect 10692 7420 10744 7472
rect 15660 7488 15712 7540
rect 15844 7531 15896 7540
rect 15844 7497 15853 7531
rect 15853 7497 15887 7531
rect 15887 7497 15896 7531
rect 15844 7488 15896 7497
rect 16212 7488 16264 7540
rect 17408 7531 17460 7540
rect 17408 7497 17417 7531
rect 17417 7497 17451 7531
rect 17451 7497 17460 7531
rect 17408 7488 17460 7497
rect 18052 7531 18104 7540
rect 18052 7497 18061 7531
rect 18061 7497 18095 7531
rect 18095 7497 18104 7531
rect 18052 7488 18104 7497
rect 19800 7488 19852 7540
rect 15292 7420 15344 7472
rect 17316 7420 17368 7472
rect 9772 7352 9824 7404
rect 10508 7352 10560 7404
rect 11244 7352 11296 7404
rect 13636 7352 13688 7404
rect 16856 7395 16908 7404
rect 16856 7361 16865 7395
rect 16865 7361 16899 7395
rect 16899 7361 16908 7395
rect 16856 7352 16908 7361
rect 19984 7420 20036 7472
rect 19248 7352 19300 7404
rect 21272 7395 21324 7404
rect 21272 7361 21281 7395
rect 21281 7361 21315 7395
rect 21315 7361 21324 7395
rect 22560 7488 22612 7540
rect 23664 7531 23716 7540
rect 23664 7497 23673 7531
rect 23673 7497 23707 7531
rect 23707 7497 23716 7531
rect 23664 7488 23716 7497
rect 23756 7488 23808 7540
rect 25136 7531 25188 7540
rect 25136 7497 25145 7531
rect 25145 7497 25179 7531
rect 25179 7497 25188 7531
rect 25136 7488 25188 7497
rect 25320 7488 25372 7540
rect 21272 7352 21324 7361
rect 23848 7352 23900 7404
rect 1952 7284 2004 7336
rect 5724 7284 5776 7336
rect 7656 7284 7708 7336
rect 9680 7284 9732 7336
rect 10600 7327 10652 7336
rect 10600 7293 10609 7327
rect 10609 7293 10643 7327
rect 10643 7293 10652 7327
rect 10600 7284 10652 7293
rect 11152 7284 11204 7336
rect 2228 7216 2280 7268
rect 5908 7216 5960 7268
rect 2136 7148 2188 7200
rect 4804 7148 4856 7200
rect 6276 7216 6328 7268
rect 6920 7216 6972 7268
rect 7104 7259 7156 7268
rect 7104 7225 7138 7259
rect 7138 7225 7156 7259
rect 7104 7216 7156 7225
rect 8668 7216 8720 7268
rect 9220 7216 9272 7268
rect 10968 7216 11020 7268
rect 12900 7284 12952 7336
rect 13452 7284 13504 7336
rect 18144 7284 18196 7336
rect 20260 7284 20312 7336
rect 22744 7284 22796 7336
rect 23112 7327 23164 7336
rect 23112 7293 23121 7327
rect 23121 7293 23155 7327
rect 23155 7293 23164 7327
rect 24676 7352 24728 7404
rect 25228 7327 25280 7336
rect 23112 7284 23164 7293
rect 25228 7293 25237 7327
rect 25237 7293 25271 7327
rect 25271 7293 25280 7327
rect 25228 7284 25280 7293
rect 14372 7216 14424 7268
rect 8944 7148 8996 7200
rect 11704 7148 11756 7200
rect 13544 7148 13596 7200
rect 16120 7191 16172 7200
rect 16120 7157 16129 7191
rect 16129 7157 16163 7191
rect 16163 7157 16172 7191
rect 18972 7216 19024 7268
rect 19892 7216 19944 7268
rect 21180 7259 21232 7268
rect 21180 7225 21189 7259
rect 21189 7225 21223 7259
rect 21223 7225 21232 7259
rect 21180 7216 21232 7225
rect 23480 7259 23532 7268
rect 23480 7225 23489 7259
rect 23489 7225 23523 7259
rect 23523 7225 23532 7259
rect 23480 7216 23532 7225
rect 16120 7148 16172 7157
rect 16856 7148 16908 7200
rect 20352 7148 20404 7200
rect 20720 7148 20772 7200
rect 21548 7148 21600 7200
rect 23296 7148 23348 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 2412 6987 2464 6996
rect 2412 6953 2421 6987
rect 2421 6953 2455 6987
rect 2455 6953 2464 6987
rect 2412 6944 2464 6953
rect 2596 6944 2648 6996
rect 4068 6944 4120 6996
rect 5632 6987 5684 6996
rect 5632 6953 5641 6987
rect 5641 6953 5675 6987
rect 5675 6953 5684 6987
rect 5632 6944 5684 6953
rect 5908 6987 5960 6996
rect 5908 6953 5917 6987
rect 5917 6953 5951 6987
rect 5951 6953 5960 6987
rect 5908 6944 5960 6953
rect 6828 6944 6880 6996
rect 8300 6987 8352 6996
rect 8300 6953 8309 6987
rect 8309 6953 8343 6987
rect 8343 6953 8352 6987
rect 8300 6944 8352 6953
rect 3516 6919 3568 6928
rect 3516 6885 3525 6919
rect 3525 6885 3559 6919
rect 3559 6885 3568 6919
rect 3516 6876 3568 6885
rect 5172 6876 5224 6928
rect 8116 6876 8168 6928
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 6276 6851 6328 6860
rect 6276 6817 6285 6851
rect 6285 6817 6319 6851
rect 6319 6817 6328 6851
rect 6276 6808 6328 6817
rect 9956 6808 10008 6860
rect 11060 6944 11112 6996
rect 11244 6944 11296 6996
rect 13176 6987 13228 6996
rect 13176 6953 13185 6987
rect 13185 6953 13219 6987
rect 13219 6953 13228 6987
rect 13176 6944 13228 6953
rect 14464 6944 14516 6996
rect 15568 6987 15620 6996
rect 15568 6953 15577 6987
rect 15577 6953 15611 6987
rect 15611 6953 15620 6987
rect 15568 6944 15620 6953
rect 16764 6944 16816 6996
rect 18144 6987 18196 6996
rect 18144 6953 18153 6987
rect 18153 6953 18187 6987
rect 18187 6953 18196 6987
rect 18144 6944 18196 6953
rect 19984 6987 20036 6996
rect 19984 6953 19993 6987
rect 19993 6953 20027 6987
rect 20027 6953 20036 6987
rect 19984 6944 20036 6953
rect 20628 6944 20680 6996
rect 21272 6944 21324 6996
rect 22560 6944 22612 6996
rect 23848 6944 23900 6996
rect 13636 6876 13688 6928
rect 18052 6876 18104 6928
rect 19432 6876 19484 6928
rect 24676 6876 24728 6928
rect 10876 6808 10928 6860
rect 16304 6851 16356 6860
rect 16304 6817 16338 6851
rect 16338 6817 16356 6851
rect 16304 6808 16356 6817
rect 18880 6851 18932 6860
rect 18880 6817 18889 6851
rect 18889 6817 18923 6851
rect 18923 6817 18932 6851
rect 18880 6808 18932 6817
rect 20628 6808 20680 6860
rect 23756 6851 23808 6860
rect 23756 6817 23765 6851
rect 23765 6817 23799 6851
rect 23799 6817 23808 6851
rect 23756 6808 23808 6817
rect 4804 6783 4856 6792
rect 1584 6715 1636 6724
rect 1584 6681 1593 6715
rect 1593 6681 1627 6715
rect 1627 6681 1636 6715
rect 1584 6672 1636 6681
rect 2504 6672 2556 6724
rect 4804 6749 4813 6783
rect 4813 6749 4847 6783
rect 4847 6749 4856 6783
rect 4804 6740 4856 6749
rect 4896 6783 4948 6792
rect 4896 6749 4905 6783
rect 4905 6749 4939 6783
rect 4939 6749 4948 6783
rect 4896 6740 4948 6749
rect 6092 6740 6144 6792
rect 6460 6740 6512 6792
rect 8484 6783 8536 6792
rect 3700 6672 3752 6724
rect 3976 6672 4028 6724
rect 8484 6749 8493 6783
rect 8493 6749 8527 6783
rect 8527 6749 8536 6783
rect 8484 6740 8536 6749
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 13360 6740 13412 6792
rect 7104 6672 7156 6724
rect 2228 6647 2280 6656
rect 2228 6613 2237 6647
rect 2237 6613 2271 6647
rect 2271 6613 2280 6647
rect 2228 6604 2280 6613
rect 3792 6647 3844 6656
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 6920 6604 6972 6656
rect 8116 6604 8168 6656
rect 8760 6672 8812 6724
rect 15844 6740 15896 6792
rect 18696 6740 18748 6792
rect 19064 6783 19116 6792
rect 19064 6749 19073 6783
rect 19073 6749 19107 6783
rect 19107 6749 19116 6783
rect 20904 6783 20956 6792
rect 19064 6740 19116 6749
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 20904 6740 20956 6749
rect 14096 6672 14148 6724
rect 8852 6647 8904 6656
rect 8852 6613 8861 6647
rect 8861 6613 8895 6647
rect 8895 6613 8904 6647
rect 8852 6604 8904 6613
rect 9220 6647 9272 6656
rect 9220 6613 9229 6647
rect 9229 6613 9263 6647
rect 9263 6613 9272 6647
rect 9220 6604 9272 6613
rect 11060 6604 11112 6656
rect 13176 6604 13228 6656
rect 13820 6604 13872 6656
rect 17408 6647 17460 6656
rect 17408 6613 17417 6647
rect 17417 6613 17451 6647
rect 17451 6613 17460 6647
rect 17408 6604 17460 6613
rect 18512 6647 18564 6656
rect 18512 6613 18521 6647
rect 18521 6613 18555 6647
rect 18555 6613 18564 6647
rect 18512 6604 18564 6613
rect 19616 6647 19668 6656
rect 19616 6613 19625 6647
rect 19625 6613 19659 6647
rect 19659 6613 19668 6647
rect 19616 6604 19668 6613
rect 21548 6604 21600 6656
rect 22744 6604 22796 6656
rect 25136 6647 25188 6656
rect 25136 6613 25145 6647
rect 25145 6613 25179 6647
rect 25179 6613 25188 6647
rect 25136 6604 25188 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2504 6443 2556 6452
rect 2504 6409 2513 6443
rect 2513 6409 2547 6443
rect 2547 6409 2556 6443
rect 2504 6400 2556 6409
rect 2780 6443 2832 6452
rect 2780 6409 2789 6443
rect 2789 6409 2823 6443
rect 2823 6409 2832 6443
rect 2780 6400 2832 6409
rect 3608 6400 3660 6452
rect 6092 6400 6144 6452
rect 6276 6443 6328 6452
rect 6276 6409 6285 6443
rect 6285 6409 6319 6443
rect 6319 6409 6328 6443
rect 6276 6400 6328 6409
rect 8484 6400 8536 6452
rect 10692 6400 10744 6452
rect 13084 6400 13136 6452
rect 13360 6443 13412 6452
rect 13360 6409 13369 6443
rect 13369 6409 13403 6443
rect 13403 6409 13412 6443
rect 13360 6400 13412 6409
rect 14372 6400 14424 6452
rect 17408 6400 17460 6452
rect 19064 6400 19116 6452
rect 23112 6443 23164 6452
rect 23112 6409 23121 6443
rect 23121 6409 23155 6443
rect 23155 6409 23164 6443
rect 23112 6400 23164 6409
rect 23756 6400 23808 6452
rect 2596 6332 2648 6384
rect 4804 6332 4856 6384
rect 5448 6332 5500 6384
rect 3240 6307 3292 6316
rect 3240 6273 3249 6307
rect 3249 6273 3283 6307
rect 3283 6273 3292 6307
rect 3240 6264 3292 6273
rect 3516 6264 3568 6316
rect 4896 6307 4948 6316
rect 4896 6273 4905 6307
rect 4905 6273 4939 6307
rect 4939 6273 4948 6307
rect 4896 6264 4948 6273
rect 9772 6332 9824 6384
rect 10968 6332 11020 6384
rect 12716 6332 12768 6384
rect 3976 6196 4028 6248
rect 4712 6239 4764 6248
rect 4712 6205 4721 6239
rect 4721 6205 4755 6239
rect 4755 6205 4764 6239
rect 4712 6196 4764 6205
rect 8024 6196 8076 6248
rect 7564 6128 7616 6180
rect 8392 6171 8444 6180
rect 8392 6137 8426 6171
rect 8426 6137 8444 6171
rect 8392 6128 8444 6137
rect 1584 6060 1636 6112
rect 8024 6103 8076 6112
rect 8024 6069 8033 6103
rect 8033 6069 8067 6103
rect 8067 6069 8076 6103
rect 8024 6060 8076 6069
rect 8852 6060 8904 6112
rect 10784 6196 10836 6248
rect 12532 6196 12584 6248
rect 16488 6264 16540 6316
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 18696 6375 18748 6384
rect 18696 6341 18705 6375
rect 18705 6341 18739 6375
rect 18739 6341 18748 6375
rect 18696 6332 18748 6341
rect 17040 6264 17092 6273
rect 22744 6264 22796 6316
rect 15844 6239 15896 6248
rect 15844 6205 15853 6239
rect 15853 6205 15887 6239
rect 15887 6205 15896 6239
rect 15844 6196 15896 6205
rect 18328 6196 18380 6248
rect 14096 6128 14148 6180
rect 10692 6060 10744 6112
rect 11060 6060 11112 6112
rect 13544 6060 13596 6112
rect 16580 6060 16632 6112
rect 17776 6128 17828 6180
rect 21732 6196 21784 6248
rect 19616 6128 19668 6180
rect 19984 6128 20036 6180
rect 23388 6196 23440 6248
rect 24400 6239 24452 6248
rect 24400 6205 24434 6239
rect 24434 6205 24452 6239
rect 24400 6196 24452 6205
rect 25136 6196 25188 6248
rect 16856 6060 16908 6112
rect 18420 6060 18472 6112
rect 20628 6103 20680 6112
rect 20628 6069 20637 6103
rect 20637 6069 20671 6103
rect 20671 6069 20680 6103
rect 20628 6060 20680 6069
rect 21732 6060 21784 6112
rect 21916 6060 21968 6112
rect 25136 6060 25188 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 2412 5856 2464 5908
rect 2688 5856 2740 5908
rect 3516 5856 3568 5908
rect 3884 5856 3936 5908
rect 4252 5856 4304 5908
rect 5540 5856 5592 5908
rect 6368 5856 6420 5908
rect 8208 5856 8260 5908
rect 9864 5856 9916 5908
rect 10876 5899 10928 5908
rect 10876 5865 10885 5899
rect 10885 5865 10919 5899
rect 10919 5865 10928 5899
rect 10876 5856 10928 5865
rect 11336 5899 11388 5908
rect 11336 5865 11345 5899
rect 11345 5865 11379 5899
rect 11379 5865 11388 5899
rect 11336 5856 11388 5865
rect 12440 5856 12492 5908
rect 13728 5856 13780 5908
rect 14096 5899 14148 5908
rect 14096 5865 14105 5899
rect 14105 5865 14139 5899
rect 14139 5865 14148 5899
rect 14096 5856 14148 5865
rect 14740 5856 14792 5908
rect 2228 5788 2280 5840
rect 4896 5788 4948 5840
rect 6276 5788 6328 5840
rect 6736 5788 6788 5840
rect 8116 5788 8168 5840
rect 13176 5788 13228 5840
rect 2688 5763 2740 5772
rect 2688 5729 2697 5763
rect 2697 5729 2731 5763
rect 2731 5729 2740 5763
rect 2688 5720 2740 5729
rect 4068 5720 4120 5772
rect 5172 5763 5224 5772
rect 5172 5729 5181 5763
rect 5181 5729 5215 5763
rect 5215 5729 5224 5763
rect 5172 5720 5224 5729
rect 7748 5720 7800 5772
rect 10048 5763 10100 5772
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 10048 5720 10100 5729
rect 2504 5652 2556 5704
rect 6092 5695 6144 5704
rect 1860 5584 1912 5636
rect 6092 5661 6101 5695
rect 6101 5661 6135 5695
rect 6135 5661 6144 5695
rect 6092 5652 6144 5661
rect 5264 5584 5316 5636
rect 6736 5652 6788 5704
rect 7104 5652 7156 5704
rect 8576 5652 8628 5704
rect 3424 5516 3476 5568
rect 8392 5584 8444 5636
rect 8760 5652 8812 5704
rect 9680 5652 9732 5704
rect 10876 5720 10928 5772
rect 11612 5763 11664 5772
rect 11612 5729 11621 5763
rect 11621 5729 11655 5763
rect 11655 5729 11664 5763
rect 11612 5720 11664 5729
rect 11980 5720 12032 5772
rect 14188 5720 14240 5772
rect 16304 5856 16356 5908
rect 16488 5899 16540 5908
rect 16488 5865 16497 5899
rect 16497 5865 16531 5899
rect 16531 5865 16540 5899
rect 16488 5856 16540 5865
rect 18880 5856 18932 5908
rect 18972 5856 19024 5908
rect 17040 5831 17092 5840
rect 17040 5797 17074 5831
rect 17074 5797 17092 5831
rect 17040 5788 17092 5797
rect 19524 5856 19576 5908
rect 21548 5899 21600 5908
rect 21548 5865 21557 5899
rect 21557 5865 21591 5899
rect 21591 5865 21600 5899
rect 21548 5856 21600 5865
rect 15844 5720 15896 5772
rect 16856 5720 16908 5772
rect 18328 5720 18380 5772
rect 22100 5856 22152 5908
rect 24400 5899 24452 5908
rect 24400 5865 24409 5899
rect 24409 5865 24443 5899
rect 24443 5865 24452 5899
rect 24400 5856 24452 5865
rect 24676 5856 24728 5908
rect 24952 5899 25004 5908
rect 24952 5865 24961 5899
rect 24961 5865 24995 5899
rect 24995 5865 25004 5899
rect 24952 5856 25004 5865
rect 23756 5788 23808 5840
rect 22376 5763 22428 5772
rect 22376 5729 22410 5763
rect 22410 5729 22428 5763
rect 10784 5652 10836 5704
rect 12716 5695 12768 5704
rect 12716 5661 12725 5695
rect 12725 5661 12759 5695
rect 12759 5661 12768 5695
rect 12716 5652 12768 5661
rect 19892 5695 19944 5704
rect 19892 5661 19901 5695
rect 19901 5661 19935 5695
rect 19935 5661 19944 5695
rect 19892 5652 19944 5661
rect 22008 5584 22060 5636
rect 22376 5720 22428 5729
rect 24768 5652 24820 5704
rect 25136 5695 25188 5704
rect 25136 5661 25145 5695
rect 25145 5661 25179 5695
rect 25179 5661 25188 5695
rect 25136 5652 25188 5661
rect 23940 5584 23992 5636
rect 6920 5516 6972 5568
rect 9404 5559 9456 5568
rect 9404 5525 9413 5559
rect 9413 5525 9447 5559
rect 9447 5525 9456 5559
rect 9404 5516 9456 5525
rect 11704 5516 11756 5568
rect 12900 5516 12952 5568
rect 13728 5516 13780 5568
rect 15936 5516 15988 5568
rect 18144 5559 18196 5568
rect 18144 5525 18153 5559
rect 18153 5525 18187 5559
rect 18187 5525 18196 5559
rect 18144 5516 18196 5525
rect 19340 5516 19392 5568
rect 20628 5559 20680 5568
rect 20628 5525 20637 5559
rect 20637 5525 20671 5559
rect 20671 5525 20680 5559
rect 20628 5516 20680 5525
rect 21456 5516 21508 5568
rect 22744 5516 22796 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 2228 5312 2280 5364
rect 2964 5312 3016 5364
rect 1860 5176 1912 5228
rect 4068 5312 4120 5364
rect 4252 5312 4304 5364
rect 5356 5312 5408 5364
rect 7104 5312 7156 5364
rect 10876 5312 10928 5364
rect 12808 5312 12860 5364
rect 8300 5244 8352 5296
rect 9220 5244 9272 5296
rect 13176 5244 13228 5296
rect 12716 5176 12768 5228
rect 14004 5219 14056 5228
rect 1584 5108 1636 5160
rect 4252 5151 4304 5160
rect 4252 5117 4261 5151
rect 4261 5117 4295 5151
rect 4295 5117 4304 5151
rect 4252 5108 4304 5117
rect 7104 5151 7156 5160
rect 7104 5117 7138 5151
rect 7138 5117 7156 5151
rect 1400 5040 1452 5092
rect 2504 5040 2556 5092
rect 5264 5040 5316 5092
rect 7104 5108 7156 5117
rect 8024 5040 8076 5092
rect 8484 5108 8536 5160
rect 9220 5108 9272 5160
rect 12440 5151 12492 5160
rect 12440 5117 12449 5151
rect 12449 5117 12483 5151
rect 12483 5117 12492 5151
rect 14004 5185 14013 5219
rect 14013 5185 14047 5219
rect 14047 5185 14056 5219
rect 14004 5176 14056 5185
rect 14372 5312 14424 5364
rect 16856 5312 16908 5364
rect 17776 5355 17828 5364
rect 17776 5321 17785 5355
rect 17785 5321 17819 5355
rect 17819 5321 17828 5355
rect 17776 5312 17828 5321
rect 19524 5312 19576 5364
rect 20444 5312 20496 5364
rect 21548 5312 21600 5364
rect 22928 5312 22980 5364
rect 24768 5312 24820 5364
rect 24952 5312 25004 5364
rect 19064 5244 19116 5296
rect 24216 5287 24268 5296
rect 24216 5253 24225 5287
rect 24225 5253 24259 5287
rect 24259 5253 24268 5287
rect 24216 5244 24268 5253
rect 19892 5176 19944 5228
rect 24676 5176 24728 5228
rect 12440 5108 12492 5117
rect 18144 5108 18196 5160
rect 9404 5040 9456 5092
rect 13820 5040 13872 5092
rect 15844 5040 15896 5092
rect 17500 5083 17552 5092
rect 17500 5049 17509 5083
rect 17509 5049 17543 5083
rect 17543 5049 17552 5083
rect 17500 5040 17552 5049
rect 1492 4972 1544 5024
rect 2688 4972 2740 5024
rect 2780 4972 2832 5024
rect 4068 4972 4120 5024
rect 5172 4972 5224 5024
rect 6092 4972 6144 5024
rect 8208 5015 8260 5024
rect 8208 4981 8217 5015
rect 8217 4981 8251 5015
rect 8251 4981 8260 5015
rect 8208 4972 8260 4981
rect 8576 4972 8628 5024
rect 9036 4972 9088 5024
rect 12440 4972 12492 5024
rect 12992 4972 13044 5024
rect 16488 5015 16540 5024
rect 16488 4981 16497 5015
rect 16497 4981 16531 5015
rect 16531 4981 16540 5015
rect 16488 4972 16540 4981
rect 20260 4972 20312 5024
rect 21732 5108 21784 5160
rect 22928 5108 22980 5160
rect 24860 5151 24912 5160
rect 24860 5117 24869 5151
rect 24869 5117 24903 5151
rect 24903 5117 24912 5151
rect 24860 5108 24912 5117
rect 20444 5040 20496 5092
rect 24216 5040 24268 5092
rect 20536 5015 20588 5024
rect 20536 4981 20545 5015
rect 20545 4981 20579 5015
rect 20579 4981 20588 5015
rect 20536 4972 20588 4981
rect 22008 4972 22060 5024
rect 22652 5015 22704 5024
rect 22652 4981 22661 5015
rect 22661 4981 22695 5015
rect 22695 4981 22704 5015
rect 22652 4972 22704 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1492 4768 1544 4820
rect 2044 4811 2096 4820
rect 2044 4777 2053 4811
rect 2053 4777 2087 4811
rect 2087 4777 2096 4811
rect 2044 4768 2096 4777
rect 2412 4811 2464 4820
rect 2412 4777 2421 4811
rect 2421 4777 2455 4811
rect 2455 4777 2464 4811
rect 2412 4768 2464 4777
rect 4160 4768 4212 4820
rect 5448 4768 5500 4820
rect 6368 4811 6420 4820
rect 6368 4777 6377 4811
rect 6377 4777 6411 4811
rect 6411 4777 6420 4811
rect 6368 4768 6420 4777
rect 6644 4768 6696 4820
rect 7932 4811 7984 4820
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 9220 4768 9272 4820
rect 10784 4768 10836 4820
rect 12532 4811 12584 4820
rect 12532 4777 12541 4811
rect 12541 4777 12575 4811
rect 12575 4777 12584 4811
rect 12532 4768 12584 4777
rect 12808 4768 12860 4820
rect 14004 4768 14056 4820
rect 14648 4768 14700 4820
rect 16028 4768 16080 4820
rect 16488 4768 16540 4820
rect 17040 4768 17092 4820
rect 18512 4768 18564 4820
rect 19156 4811 19208 4820
rect 19156 4777 19165 4811
rect 19165 4777 19199 4811
rect 19199 4777 19208 4811
rect 19156 4768 19208 4777
rect 19340 4768 19392 4820
rect 20444 4768 20496 4820
rect 20812 4768 20864 4820
rect 21640 4768 21692 4820
rect 22376 4768 22428 4820
rect 24768 4768 24820 4820
rect 3792 4700 3844 4752
rect 6552 4700 6604 4752
rect 7196 4700 7248 4752
rect 8024 4700 8076 4752
rect 11244 4700 11296 4752
rect 11520 4700 11572 4752
rect 13912 4700 13964 4752
rect 16580 4700 16632 4752
rect 17408 4700 17460 4752
rect 19064 4743 19116 4752
rect 19064 4709 19073 4743
rect 19073 4709 19107 4743
rect 19107 4709 19116 4743
rect 19064 4700 19116 4709
rect 5264 4632 5316 4684
rect 5540 4632 5592 4684
rect 8300 4675 8352 4684
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 9956 4632 10008 4684
rect 10876 4632 10928 4684
rect 14004 4675 14056 4684
rect 14004 4641 14013 4675
rect 14013 4641 14047 4675
rect 14047 4641 14056 4675
rect 14004 4632 14056 4641
rect 16212 4632 16264 4684
rect 19524 4632 19576 4684
rect 20536 4700 20588 4752
rect 20996 4700 21048 4752
rect 21916 4700 21968 4752
rect 25136 4700 25188 4752
rect 22008 4632 22060 4684
rect 22744 4675 22796 4684
rect 22744 4641 22778 4675
rect 22778 4641 22796 4675
rect 22744 4632 22796 4641
rect 24952 4675 25004 4684
rect 24952 4641 24961 4675
rect 24961 4641 24995 4675
rect 24995 4641 25004 4675
rect 24952 4632 25004 4641
rect 3240 4564 3292 4616
rect 5356 4607 5408 4616
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 6644 4564 6696 4616
rect 8208 4564 8260 4616
rect 7472 4539 7524 4548
rect 7472 4505 7481 4539
rect 7481 4505 7515 4539
rect 7515 4505 7524 4539
rect 7472 4496 7524 4505
rect 14096 4564 14148 4616
rect 17500 4607 17552 4616
rect 10784 4496 10836 4548
rect 3056 4471 3108 4480
rect 3056 4437 3065 4471
rect 3065 4437 3099 4471
rect 3099 4437 3108 4471
rect 3056 4428 3108 4437
rect 4160 4428 4212 4480
rect 5448 4428 5500 4480
rect 6368 4428 6420 4480
rect 6644 4428 6696 4480
rect 7012 4428 7064 4480
rect 8852 4428 8904 4480
rect 9128 4428 9180 4480
rect 10048 4428 10100 4480
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 15660 4496 15712 4548
rect 17500 4573 17509 4607
rect 17509 4573 17543 4607
rect 17543 4573 17552 4607
rect 17500 4564 17552 4573
rect 19708 4607 19760 4616
rect 19708 4573 19717 4607
rect 19717 4573 19751 4607
rect 19751 4573 19760 4607
rect 19708 4564 19760 4573
rect 20628 4564 20680 4616
rect 22284 4564 22336 4616
rect 17684 4496 17736 4548
rect 12532 4428 12584 4480
rect 13176 4471 13228 4480
rect 13176 4437 13185 4471
rect 13185 4437 13219 4471
rect 13219 4437 13228 4471
rect 13176 4428 13228 4437
rect 13544 4471 13596 4480
rect 13544 4437 13553 4471
rect 13553 4437 13587 4471
rect 13587 4437 13596 4471
rect 13544 4428 13596 4437
rect 14740 4471 14792 4480
rect 14740 4437 14749 4471
rect 14749 4437 14783 4471
rect 14783 4437 14792 4471
rect 14740 4428 14792 4437
rect 15292 4471 15344 4480
rect 15292 4437 15301 4471
rect 15301 4437 15335 4471
rect 15335 4437 15344 4471
rect 15292 4428 15344 4437
rect 18328 4471 18380 4480
rect 18328 4437 18337 4471
rect 18337 4437 18371 4471
rect 18371 4437 18380 4471
rect 18328 4428 18380 4437
rect 18880 4428 18932 4480
rect 23848 4471 23900 4480
rect 23848 4437 23857 4471
rect 23857 4437 23891 4471
rect 23891 4437 23900 4471
rect 23848 4428 23900 4437
rect 27068 4428 27120 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 6552 4224 6604 4276
rect 10232 4224 10284 4276
rect 11060 4224 11112 4276
rect 13912 4224 13964 4276
rect 14004 4224 14056 4276
rect 16212 4267 16264 4276
rect 16212 4233 16221 4267
rect 16221 4233 16255 4267
rect 16255 4233 16264 4267
rect 16212 4224 16264 4233
rect 17500 4224 17552 4276
rect 19708 4224 19760 4276
rect 21640 4224 21692 4276
rect 22744 4224 22796 4276
rect 24952 4224 25004 4276
rect 5356 4156 5408 4208
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 6736 4156 6788 4208
rect 7472 4156 7524 4208
rect 1952 4088 2004 4097
rect 7564 4088 7616 4140
rect 9128 4156 9180 4208
rect 10876 4156 10928 4208
rect 11244 4156 11296 4208
rect 13176 4156 13228 4208
rect 9864 4131 9916 4140
rect 6000 4020 6052 4072
rect 6368 4020 6420 4072
rect 7932 4020 7984 4072
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 13360 4088 13412 4140
rect 14556 4131 14608 4140
rect 14556 4097 14565 4131
rect 14565 4097 14599 4131
rect 14599 4097 14608 4131
rect 14556 4088 14608 4097
rect 14740 4088 14792 4140
rect 9404 4063 9456 4072
rect 9404 4029 9413 4063
rect 9413 4029 9447 4063
rect 9447 4029 9456 4063
rect 9404 4020 9456 4029
rect 10692 4020 10744 4072
rect 3240 3952 3292 4004
rect 2872 3884 2924 3936
rect 4068 3927 4120 3936
rect 4068 3893 4077 3927
rect 4077 3893 4111 3927
rect 4111 3893 4120 3927
rect 4068 3884 4120 3893
rect 6092 3884 6144 3936
rect 6368 3884 6420 3936
rect 6828 3927 6880 3936
rect 6828 3893 6837 3927
rect 6837 3893 6871 3927
rect 6871 3893 6880 3927
rect 6828 3884 6880 3893
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 8208 3884 8260 3936
rect 8392 3927 8444 3936
rect 8392 3893 8401 3927
rect 8401 3893 8435 3927
rect 8435 3893 8444 3927
rect 8392 3884 8444 3893
rect 10048 3884 10100 3936
rect 11428 4020 11480 4072
rect 12164 4063 12216 4072
rect 12164 4029 12173 4063
rect 12173 4029 12207 4063
rect 12207 4029 12216 4063
rect 12164 4020 12216 4029
rect 12716 4020 12768 4072
rect 13176 4020 13228 4072
rect 15016 3995 15068 4004
rect 15016 3961 15025 3995
rect 15025 3961 15059 3995
rect 15059 3961 15068 3995
rect 15016 3952 15068 3961
rect 12440 3884 12492 3936
rect 15568 3952 15620 4004
rect 17684 4088 17736 4140
rect 18236 4088 18288 4140
rect 18328 4088 18380 4140
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 18880 4131 18932 4140
rect 18880 4097 18889 4131
rect 18889 4097 18923 4131
rect 18923 4097 18932 4131
rect 18880 4088 18932 4097
rect 21916 4088 21968 4140
rect 22100 4088 22152 4140
rect 23572 4088 23624 4140
rect 25136 4088 25188 4140
rect 16580 4063 16632 4072
rect 16580 4029 16589 4063
rect 16589 4029 16623 4063
rect 16623 4029 16632 4063
rect 16580 4020 16632 4029
rect 20536 4020 20588 4072
rect 22468 4063 22520 4072
rect 22468 4029 22477 4063
rect 22477 4029 22511 4063
rect 22511 4029 22520 4063
rect 22468 4020 22520 4029
rect 23664 4020 23716 4072
rect 16396 3952 16448 4004
rect 22284 3952 22336 4004
rect 23848 3952 23900 4004
rect 24032 4020 24084 4072
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 15660 3884 15712 3893
rect 15936 3927 15988 3936
rect 15936 3893 15945 3927
rect 15945 3893 15979 3927
rect 15979 3893 15988 3927
rect 15936 3884 15988 3893
rect 18236 3927 18288 3936
rect 18236 3893 18245 3927
rect 18245 3893 18279 3927
rect 18279 3893 18288 3927
rect 18236 3884 18288 3893
rect 20536 3927 20588 3936
rect 20536 3893 20545 3927
rect 20545 3893 20579 3927
rect 20579 3893 20588 3927
rect 20536 3884 20588 3893
rect 20720 3927 20772 3936
rect 20720 3893 20729 3927
rect 20729 3893 20763 3927
rect 20763 3893 20772 3927
rect 20720 3884 20772 3893
rect 21180 3927 21232 3936
rect 21180 3893 21189 3927
rect 21189 3893 21223 3927
rect 21223 3893 21232 3927
rect 22652 3927 22704 3936
rect 21180 3884 21232 3893
rect 22652 3893 22661 3927
rect 22661 3893 22695 3927
rect 22695 3893 22704 3927
rect 22652 3884 22704 3893
rect 23204 3884 23256 3936
rect 24032 3884 24084 3936
rect 24216 3952 24268 4004
rect 25136 3927 25188 3936
rect 25136 3893 25145 3927
rect 25145 3893 25179 3927
rect 25179 3893 25188 3927
rect 25136 3884 25188 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 2044 3680 2096 3732
rect 3240 3680 3292 3732
rect 5264 3680 5316 3732
rect 5540 3680 5592 3732
rect 8024 3723 8076 3732
rect 8024 3689 8033 3723
rect 8033 3689 8067 3723
rect 8067 3689 8076 3723
rect 8024 3680 8076 3689
rect 10048 3680 10100 3732
rect 10692 3723 10744 3732
rect 10692 3689 10701 3723
rect 10701 3689 10735 3723
rect 10735 3689 10744 3723
rect 10692 3680 10744 3689
rect 12164 3723 12216 3732
rect 12164 3689 12173 3723
rect 12173 3689 12207 3723
rect 12207 3689 12216 3723
rect 12164 3680 12216 3689
rect 12624 3680 12676 3732
rect 13268 3723 13320 3732
rect 13268 3689 13277 3723
rect 13277 3689 13311 3723
rect 13311 3689 13320 3723
rect 13268 3680 13320 3689
rect 14096 3680 14148 3732
rect 14740 3680 14792 3732
rect 15384 3680 15436 3732
rect 15936 3680 15988 3732
rect 16212 3680 16264 3732
rect 17224 3680 17276 3732
rect 17408 3723 17460 3732
rect 17408 3689 17417 3723
rect 17417 3689 17451 3723
rect 17451 3689 17460 3723
rect 17408 3680 17460 3689
rect 18052 3723 18104 3732
rect 18052 3689 18061 3723
rect 18061 3689 18095 3723
rect 18095 3689 18104 3723
rect 18052 3680 18104 3689
rect 18236 3680 18288 3732
rect 18696 3680 18748 3732
rect 18880 3680 18932 3732
rect 19432 3680 19484 3732
rect 19524 3723 19576 3732
rect 19524 3689 19533 3723
rect 19533 3689 19567 3723
rect 19567 3689 19576 3723
rect 19524 3680 19576 3689
rect 20720 3680 20772 3732
rect 21364 3723 21416 3732
rect 21364 3689 21373 3723
rect 21373 3689 21407 3723
rect 21407 3689 21416 3723
rect 21364 3680 21416 3689
rect 21916 3723 21968 3732
rect 21916 3689 21925 3723
rect 21925 3689 21959 3723
rect 21959 3689 21968 3723
rect 21916 3680 21968 3689
rect 22192 3680 22244 3732
rect 2412 3655 2464 3664
rect 2412 3621 2421 3655
rect 2421 3621 2455 3655
rect 2455 3621 2464 3655
rect 2412 3612 2464 3621
rect 3332 3612 3384 3664
rect 4068 3612 4120 3664
rect 2872 3476 2924 3528
rect 3884 3476 3936 3528
rect 4160 3544 4212 3596
rect 6552 3544 6604 3596
rect 9956 3612 10008 3664
rect 11060 3655 11112 3664
rect 11060 3621 11094 3655
rect 11094 3621 11112 3655
rect 11060 3612 11112 3621
rect 11980 3612 12032 3664
rect 12256 3612 12308 3664
rect 6736 3476 6788 3528
rect 2136 3408 2188 3460
rect 1860 3340 1912 3392
rect 4344 3340 4396 3392
rect 5540 3340 5592 3392
rect 7380 3408 7432 3460
rect 10876 3544 10928 3596
rect 13176 3587 13228 3596
rect 13176 3553 13185 3587
rect 13185 3553 13219 3587
rect 13219 3553 13228 3587
rect 13176 3544 13228 3553
rect 13360 3544 13412 3596
rect 15292 3544 15344 3596
rect 16212 3544 16264 3596
rect 16396 3587 16448 3596
rect 16396 3553 16405 3587
rect 16405 3553 16439 3587
rect 16439 3553 16448 3587
rect 16396 3544 16448 3553
rect 17500 3612 17552 3664
rect 18604 3612 18656 3664
rect 20904 3612 20956 3664
rect 20076 3544 20128 3596
rect 20996 3544 21048 3596
rect 22468 3680 22520 3732
rect 23848 3655 23900 3664
rect 23848 3621 23882 3655
rect 23882 3621 23900 3655
rect 23848 3612 23900 3621
rect 23572 3587 23624 3596
rect 23572 3553 23581 3587
rect 23581 3553 23615 3587
rect 23615 3553 23624 3587
rect 23572 3544 23624 3553
rect 7656 3519 7708 3528
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 8576 3519 8628 3528
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 8576 3476 8628 3485
rect 13728 3519 13780 3528
rect 13728 3485 13737 3519
rect 13737 3485 13771 3519
rect 13771 3485 13780 3519
rect 13728 3476 13780 3485
rect 13820 3519 13872 3528
rect 13820 3485 13829 3519
rect 13829 3485 13863 3519
rect 13863 3485 13872 3519
rect 15844 3519 15896 3528
rect 13820 3476 13872 3485
rect 15844 3485 15853 3519
rect 15853 3485 15887 3519
rect 15887 3485 15896 3519
rect 15844 3476 15896 3485
rect 18512 3476 18564 3528
rect 21456 3519 21508 3528
rect 21456 3485 21465 3519
rect 21465 3485 21499 3519
rect 21499 3485 21508 3519
rect 21456 3476 21508 3485
rect 8208 3340 8260 3392
rect 9588 3340 9640 3392
rect 9864 3383 9916 3392
rect 9864 3349 9873 3383
rect 9873 3349 9907 3383
rect 9907 3349 9916 3383
rect 9864 3340 9916 3349
rect 11152 3340 11204 3392
rect 14556 3340 14608 3392
rect 15016 3408 15068 3460
rect 18144 3408 18196 3460
rect 21272 3408 21324 3460
rect 19892 3383 19944 3392
rect 19892 3349 19901 3383
rect 19901 3349 19935 3383
rect 19935 3349 19944 3383
rect 19892 3340 19944 3349
rect 22652 3383 22704 3392
rect 22652 3349 22661 3383
rect 22661 3349 22695 3383
rect 22695 3349 22704 3383
rect 22652 3340 22704 3349
rect 24768 3340 24820 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1952 3136 2004 3188
rect 3240 3136 3292 3188
rect 4620 3136 4672 3188
rect 6828 3179 6880 3188
rect 1676 2932 1728 2984
rect 1860 2975 1912 2984
rect 1860 2941 1894 2975
rect 1894 2941 1912 2975
rect 1860 2932 1912 2941
rect 3884 2864 3936 2916
rect 4344 2932 4396 2984
rect 5448 2932 5500 2984
rect 6828 3145 6837 3179
rect 6837 3145 6871 3179
rect 6871 3145 6880 3179
rect 6828 3136 6880 3145
rect 7932 3179 7984 3188
rect 7932 3145 7941 3179
rect 7941 3145 7975 3179
rect 7975 3145 7984 3179
rect 7932 3136 7984 3145
rect 8484 3136 8536 3188
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 10232 3136 10284 3188
rect 10876 3179 10928 3188
rect 10876 3145 10885 3179
rect 10885 3145 10919 3179
rect 10919 3145 10928 3179
rect 10876 3136 10928 3145
rect 11796 3179 11848 3188
rect 11796 3145 11805 3179
rect 11805 3145 11839 3179
rect 11839 3145 11848 3179
rect 11796 3136 11848 3145
rect 12900 3136 12952 3188
rect 13820 3136 13872 3188
rect 15844 3136 15896 3188
rect 17500 3179 17552 3188
rect 17500 3145 17509 3179
rect 17509 3145 17543 3179
rect 17543 3145 17552 3179
rect 17500 3136 17552 3145
rect 17776 3179 17828 3188
rect 17776 3145 17785 3179
rect 17785 3145 17819 3179
rect 17819 3145 17828 3179
rect 17776 3136 17828 3145
rect 19432 3179 19484 3188
rect 19432 3145 19441 3179
rect 19441 3145 19475 3179
rect 19475 3145 19484 3179
rect 19432 3136 19484 3145
rect 20904 3136 20956 3188
rect 21456 3136 21508 3188
rect 22560 3136 22612 3188
rect 23572 3136 23624 3188
rect 9956 3068 10008 3120
rect 7472 2932 7524 2984
rect 8484 2932 8536 2984
rect 10876 3000 10928 3052
rect 12440 3111 12492 3120
rect 12440 3077 12449 3111
rect 12449 3077 12483 3111
rect 12483 3077 12492 3111
rect 12440 3068 12492 3077
rect 13360 3068 13412 3120
rect 16212 3068 16264 3120
rect 21916 3111 21968 3120
rect 21916 3077 21925 3111
rect 21925 3077 21959 3111
rect 21959 3077 21968 3111
rect 21916 3068 21968 3077
rect 23848 3068 23900 3120
rect 18052 3043 18104 3052
rect 18052 3009 18061 3043
rect 18061 3009 18095 3043
rect 18095 3009 18104 3043
rect 18052 3000 18104 3009
rect 24032 3136 24084 3188
rect 25136 3136 25188 3188
rect 26056 3179 26108 3188
rect 26056 3145 26065 3179
rect 26065 3145 26099 3179
rect 26099 3145 26108 3179
rect 26056 3136 26108 3145
rect 9036 2975 9088 2984
rect 9036 2941 9070 2975
rect 9070 2941 9088 2975
rect 9036 2932 9088 2941
rect 9312 2932 9364 2984
rect 9588 2932 9640 2984
rect 11336 2932 11388 2984
rect 12900 2975 12952 2984
rect 12900 2941 12909 2975
rect 12909 2941 12943 2975
rect 12943 2941 12952 2975
rect 12900 2932 12952 2941
rect 2780 2796 2832 2848
rect 5632 2839 5684 2848
rect 5632 2805 5641 2839
rect 5641 2805 5675 2839
rect 5675 2805 5684 2839
rect 5632 2796 5684 2805
rect 6092 2864 6144 2916
rect 6460 2864 6512 2916
rect 6552 2907 6604 2916
rect 6552 2873 6561 2907
rect 6561 2873 6595 2907
rect 6595 2873 6604 2907
rect 6552 2864 6604 2873
rect 12624 2864 12676 2916
rect 7932 2796 7984 2848
rect 11428 2839 11480 2848
rect 11428 2805 11437 2839
rect 11437 2805 11471 2839
rect 11471 2805 11480 2839
rect 11428 2796 11480 2805
rect 11520 2796 11572 2848
rect 13728 2796 13780 2848
rect 14464 2796 14516 2848
rect 18144 2932 18196 2984
rect 14832 2864 14884 2916
rect 15016 2907 15068 2916
rect 15016 2873 15028 2907
rect 15028 2873 15068 2907
rect 15016 2864 15068 2873
rect 18052 2864 18104 2916
rect 24768 2932 24820 2984
rect 20720 2864 20772 2916
rect 20904 2796 20956 2848
rect 23480 2796 23532 2848
rect 24032 2796 24084 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1676 2635 1728 2644
rect 1676 2601 1685 2635
rect 1685 2601 1719 2635
rect 1719 2601 1728 2635
rect 1676 2592 1728 2601
rect 2412 2592 2464 2644
rect 2872 2635 2924 2644
rect 2872 2601 2881 2635
rect 2881 2601 2915 2635
rect 2915 2601 2924 2635
rect 2872 2592 2924 2601
rect 3884 2635 3936 2644
rect 3884 2601 3893 2635
rect 3893 2601 3927 2635
rect 3927 2601 3936 2635
rect 3884 2592 3936 2601
rect 5448 2592 5500 2644
rect 8484 2592 8536 2644
rect 9772 2635 9824 2644
rect 9772 2601 9781 2635
rect 9781 2601 9815 2635
rect 9815 2601 9824 2635
rect 9772 2592 9824 2601
rect 10140 2635 10192 2644
rect 10140 2601 10149 2635
rect 10149 2601 10183 2635
rect 10183 2601 10192 2635
rect 10140 2592 10192 2601
rect 11060 2592 11112 2644
rect 14004 2635 14056 2644
rect 14004 2601 14013 2635
rect 14013 2601 14047 2635
rect 14047 2601 14056 2635
rect 14004 2592 14056 2601
rect 16856 2635 16908 2644
rect 16856 2601 16865 2635
rect 16865 2601 16899 2635
rect 16899 2601 16908 2635
rect 16856 2592 16908 2601
rect 18052 2635 18104 2644
rect 18052 2601 18061 2635
rect 18061 2601 18095 2635
rect 18095 2601 18104 2635
rect 18052 2592 18104 2601
rect 18144 2592 18196 2644
rect 18512 2592 18564 2644
rect 20720 2592 20772 2644
rect 20904 2635 20956 2644
rect 20904 2601 20913 2635
rect 20913 2601 20947 2635
rect 20947 2601 20956 2635
rect 20904 2592 20956 2601
rect 2320 2567 2372 2576
rect 2320 2533 2329 2567
rect 2329 2533 2363 2567
rect 2363 2533 2372 2567
rect 2320 2524 2372 2533
rect 2228 2499 2280 2508
rect 2228 2465 2237 2499
rect 2237 2465 2271 2499
rect 2271 2465 2280 2499
rect 2228 2456 2280 2465
rect 7656 2524 7708 2576
rect 4620 2499 4672 2508
rect 3240 2388 3292 2440
rect 4620 2465 4654 2499
rect 4654 2465 4672 2499
rect 4620 2456 4672 2465
rect 6736 2456 6788 2508
rect 9680 2524 9732 2576
rect 12808 2524 12860 2576
rect 8300 2320 8352 2372
rect 9956 2456 10008 2508
rect 11244 2499 11296 2508
rect 11244 2465 11253 2499
rect 11253 2465 11287 2499
rect 11287 2465 11296 2499
rect 11244 2456 11296 2465
rect 296 2252 348 2304
rect 1308 2252 1360 2304
rect 6552 2252 6604 2304
rect 10876 2388 10928 2440
rect 14464 2456 14516 2508
rect 18696 2524 18748 2576
rect 22008 2592 22060 2644
rect 22560 2635 22612 2644
rect 22560 2601 22569 2635
rect 22569 2601 22603 2635
rect 22603 2601 22612 2635
rect 22560 2592 22612 2601
rect 23756 2635 23808 2644
rect 23756 2601 23765 2635
rect 23765 2601 23799 2635
rect 23799 2601 23808 2635
rect 23756 2592 23808 2601
rect 24216 2635 24268 2644
rect 24216 2601 24225 2635
rect 24225 2601 24259 2635
rect 24259 2601 24268 2635
rect 24216 2592 24268 2601
rect 21916 2524 21968 2576
rect 18144 2388 18196 2440
rect 24492 2388 24544 2440
rect 24768 2431 24820 2440
rect 24768 2397 24777 2431
rect 24777 2397 24811 2431
rect 24811 2397 24820 2431
rect 24768 2388 24820 2397
rect 9772 2320 9824 2372
rect 11704 2320 11756 2372
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 2044 2048 2096 2100
rect 6368 2048 6420 2100
rect 11796 1640 11848 1692
rect 18880 1640 18932 1692
rect 3792 552 3844 604
rect 4528 552 4580 604
rect 7748 552 7800 604
rect 9036 552 9088 604
rect 10692 552 10744 604
rect 10784 552 10836 604
rect 11336 552 11388 604
rect 12348 552 12400 604
rect 21272 552 21324 604
rect 21548 552 21600 604
rect 4344 484 4396 536
rect 5172 484 5224 536
<< metal2 >>
rect 2778 27568 2834 27577
rect 4618 27520 4674 28000
rect 13910 27520 13966 28000
rect 23202 27520 23258 28000
rect 23478 27568 23534 27577
rect 2778 27503 2834 27512
rect 1950 26208 2006 26217
rect 1950 26143 2006 26152
rect 1582 24848 1638 24857
rect 1582 24783 1638 24792
rect 1596 22778 1624 24783
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1768 22568 1820 22574
rect 1768 22510 1820 22516
rect 1582 22128 1638 22137
rect 1582 22063 1638 22072
rect 1490 21448 1546 21457
rect 1490 21383 1546 21392
rect 1398 20768 1454 20777
rect 1398 20703 1454 20712
rect 1412 19174 1440 20703
rect 1504 20058 1532 21383
rect 1596 20602 1624 22063
rect 1780 21146 1808 22510
rect 1768 21140 1820 21146
rect 1768 21082 1820 21088
rect 1858 20768 1914 20777
rect 1858 20703 1914 20712
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1582 20088 1638 20097
rect 1492 20052 1544 20058
rect 1582 20023 1638 20032
rect 1492 19994 1544 20000
rect 1400 19168 1452 19174
rect 1400 19110 1452 19116
rect 1490 18728 1546 18737
rect 1490 18663 1546 18672
rect 1398 17368 1454 17377
rect 1504 17338 1532 18663
rect 1596 18426 1624 20023
rect 1674 19408 1730 19417
rect 1674 19343 1730 19352
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 1582 18048 1638 18057
rect 1582 17983 1638 17992
rect 1398 17303 1454 17312
rect 1492 17332 1544 17338
rect 1412 15706 1440 17303
rect 1492 17274 1544 17280
rect 1596 16794 1624 17983
rect 1688 17882 1716 19343
rect 1780 18970 1808 20198
rect 1768 18964 1820 18970
rect 1768 18906 1820 18912
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1582 16008 1638 16017
rect 1582 15943 1638 15952
rect 1400 15700 1452 15706
rect 1400 15642 1452 15648
rect 1490 14648 1546 14657
rect 1596 14618 1624 15943
rect 1872 15688 1900 20703
rect 1964 16810 1992 26143
rect 2226 24168 2282 24177
rect 2226 24103 2282 24112
rect 2042 23488 2098 23497
rect 2042 23423 2098 23432
rect 2056 20777 2084 23423
rect 2042 20768 2098 20777
rect 2042 20703 2098 20712
rect 2136 19916 2188 19922
rect 2136 19858 2188 19864
rect 2148 19174 2176 19858
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 2044 18080 2096 18086
rect 2042 18048 2044 18057
rect 2096 18048 2098 18057
rect 2042 17983 2098 17992
rect 2148 17241 2176 19110
rect 2134 17232 2190 17241
rect 2134 17167 2190 17176
rect 1964 16782 2176 16810
rect 1950 16688 2006 16697
rect 1950 16623 2006 16632
rect 1780 15660 1900 15688
rect 1674 15328 1730 15337
rect 1674 15263 1730 15272
rect 1490 14583 1546 14592
rect 1584 14612 1636 14618
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1412 14074 1440 14418
rect 1400 14068 1452 14074
rect 1400 14010 1452 14016
rect 1400 13524 1452 13530
rect 1400 13466 1452 13472
rect 1412 12782 1440 13466
rect 1504 12986 1532 14583
rect 1584 14554 1636 14560
rect 1582 13968 1638 13977
rect 1582 13903 1638 13912
rect 1492 12980 1544 12986
rect 1492 12922 1544 12928
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1400 12640 1452 12646
rect 1400 12582 1452 12588
rect 1308 9376 1360 9382
rect 1308 9318 1360 9324
rect 846 2816 902 2825
rect 846 2751 902 2760
rect 296 2304 348 2310
rect 296 2246 348 2252
rect 308 480 336 2246
rect 860 480 888 2751
rect 1320 2310 1348 9318
rect 1412 9042 1440 12582
rect 1492 12436 1544 12442
rect 1492 12378 1544 12384
rect 1504 11354 1532 12378
rect 1492 11348 1544 11354
rect 1492 11290 1544 11296
rect 1492 9988 1544 9994
rect 1492 9930 1544 9936
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1400 7744 1452 7750
rect 1400 7686 1452 7692
rect 1412 6866 1440 7686
rect 1504 7018 1532 9930
rect 1596 9654 1624 13903
rect 1688 13190 1716 15263
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1584 9648 1636 9654
rect 1584 9590 1636 9596
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1596 9178 1624 9454
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1688 8022 1716 12922
rect 1780 12442 1808 15660
rect 1860 15564 1912 15570
rect 1860 15506 1912 15512
rect 1872 14822 1900 15506
rect 1964 15162 1992 16623
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 2056 14929 2084 15846
rect 2042 14920 2098 14929
rect 2042 14855 2098 14864
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 1872 12986 1900 14758
rect 1952 14272 2004 14278
rect 1952 14214 2004 14220
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1964 12306 1992 14214
rect 2148 14006 2176 16782
rect 2240 16130 2268 24103
rect 2504 21004 2556 21010
rect 2504 20946 2556 20952
rect 2516 20262 2544 20946
rect 2504 20256 2556 20262
rect 2504 20198 2556 20204
rect 2410 19272 2466 19281
rect 2410 19207 2412 19216
rect 2464 19207 2466 19216
rect 2412 19178 2464 19184
rect 2410 18864 2466 18873
rect 2410 18799 2412 18808
rect 2464 18799 2466 18808
rect 2412 18770 2464 18776
rect 2424 18426 2452 18770
rect 2516 18737 2544 20198
rect 2502 18728 2558 18737
rect 2502 18663 2558 18672
rect 2412 18420 2464 18426
rect 2412 18362 2464 18368
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 2332 17338 2360 17682
rect 2320 17332 2372 17338
rect 2320 17274 2372 17280
rect 2332 16250 2360 17274
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2240 16102 2360 16130
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 2136 14000 2188 14006
rect 2136 13942 2188 13948
rect 2044 13864 2096 13870
rect 2042 13832 2044 13841
rect 2136 13864 2188 13870
rect 2096 13832 2098 13841
rect 2136 13806 2188 13812
rect 2042 13767 2098 13776
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2056 12782 2084 13330
rect 2044 12776 2096 12782
rect 2042 12744 2044 12753
rect 2096 12744 2098 12753
rect 2042 12679 2098 12688
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 2056 12306 2084 12582
rect 1952 12300 2004 12306
rect 1952 12242 2004 12248
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 1860 12232 1912 12238
rect 1860 12174 1912 12180
rect 1964 12186 1992 12242
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1676 8016 1728 8022
rect 1676 7958 1728 7964
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1688 7546 1716 7822
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1504 6990 1716 7018
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1412 5953 1440 6802
rect 1582 6760 1638 6769
rect 1582 6695 1584 6704
rect 1636 6695 1638 6704
rect 1584 6666 1636 6672
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1398 5944 1454 5953
rect 1596 5914 1624 6054
rect 1398 5879 1454 5888
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1596 5166 1624 5850
rect 1584 5160 1636 5166
rect 1490 5128 1546 5137
rect 1400 5092 1452 5098
rect 1584 5102 1636 5108
rect 1490 5063 1546 5072
rect 1400 5034 1452 5040
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1412 480 1440 5034
rect 1504 5030 1532 5063
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 1504 4826 1532 4966
rect 1492 4820 1544 4826
rect 1492 4762 1544 4768
rect 1688 4729 1716 6990
rect 1674 4720 1730 4729
rect 1674 4655 1730 4664
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1688 2650 1716 2926
rect 1780 2802 1808 9862
rect 1872 9450 1900 12174
rect 1964 12158 2084 12186
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1964 11762 1992 12038
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 2056 11286 2084 12158
rect 2044 11280 2096 11286
rect 2044 11222 2096 11228
rect 2042 10704 2098 10713
rect 2042 10639 2044 10648
rect 2096 10639 2098 10648
rect 2044 10610 2096 10616
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1872 7721 1900 8978
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1964 8362 1992 8774
rect 1952 8356 2004 8362
rect 1952 8298 2004 8304
rect 2148 8090 2176 13806
rect 2240 12646 2268 14010
rect 2332 13274 2360 16102
rect 2424 15910 2452 16594
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2424 15473 2452 15846
rect 2410 15464 2466 15473
rect 2410 15399 2466 15408
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2516 14618 2544 14758
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 2792 14482 2820 27503
rect 4632 27418 4660 27520
rect 4172 27390 4660 27418
rect 3054 26888 3110 26897
rect 3054 26823 3110 26832
rect 2870 25528 2926 25537
rect 2870 25463 2926 25472
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2780 14340 2832 14346
rect 2780 14282 2832 14288
rect 2688 13728 2740 13734
rect 2688 13670 2740 13676
rect 2700 13530 2728 13670
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 2792 13410 2820 14282
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2700 13382 2820 13410
rect 2332 13246 2452 13274
rect 2320 12844 2372 12850
rect 2320 12786 2372 12792
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2226 12472 2282 12481
rect 2226 12407 2282 12416
rect 2240 11898 2268 12407
rect 2332 11898 2360 12786
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 2332 11354 2360 11562
rect 2424 11354 2452 13246
rect 2516 12170 2544 13330
rect 2596 13252 2648 13258
rect 2596 13194 2648 13200
rect 2608 12850 2636 13194
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2700 12442 2728 13382
rect 2884 13326 2912 25463
rect 2962 22808 3018 22817
rect 2962 22743 3018 22752
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2870 13152 2926 13161
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2504 12164 2556 12170
rect 2504 12106 2556 12112
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2332 10470 2360 11154
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2240 8430 2268 9114
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2332 8129 2360 10406
rect 2410 10296 2466 10305
rect 2410 10231 2412 10240
rect 2464 10231 2466 10240
rect 2412 10202 2464 10208
rect 2516 8514 2544 11834
rect 2686 11656 2742 11665
rect 2686 11591 2688 11600
rect 2740 11591 2742 11600
rect 2688 11562 2740 11568
rect 2596 11552 2648 11558
rect 2594 11520 2596 11529
rect 2648 11520 2650 11529
rect 2594 11455 2650 11464
rect 2792 11098 2820 13126
rect 2870 13087 2926 13096
rect 2884 11218 2912 13087
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2700 11070 2820 11098
rect 2872 11076 2924 11082
rect 2596 9988 2648 9994
rect 2596 9930 2648 9936
rect 2608 9654 2636 9930
rect 2596 9648 2648 9654
rect 2596 9590 2648 9596
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2608 8634 2636 8910
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2424 8486 2544 8514
rect 2318 8120 2374 8129
rect 2136 8084 2188 8090
rect 2424 8106 2452 8486
rect 2502 8392 2558 8401
rect 2502 8327 2504 8336
rect 2556 8327 2558 8336
rect 2504 8298 2556 8304
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2424 8090 2544 8106
rect 2424 8084 2556 8090
rect 2424 8078 2504 8084
rect 2318 8055 2374 8064
rect 2136 8026 2188 8032
rect 2504 8026 2556 8032
rect 2228 8016 2280 8022
rect 2226 7984 2228 7993
rect 2412 8016 2464 8022
rect 2280 7984 2282 7993
rect 2412 7958 2464 7964
rect 2226 7919 2282 7928
rect 1858 7712 1914 7721
rect 1858 7647 1914 7656
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1860 5636 1912 5642
rect 1860 5578 1912 5584
rect 1872 5234 1900 5578
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1872 3398 1900 5170
rect 1964 4146 1992 7278
rect 2228 7268 2280 7274
rect 2228 7210 2280 7216
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 2042 5672 2098 5681
rect 2042 5607 2098 5616
rect 2056 4826 2084 5607
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1872 2990 1900 3334
rect 1964 3194 1992 4082
rect 2056 3738 2084 4762
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 2148 3466 2176 7142
rect 2240 6662 2268 7210
rect 2424 7002 2452 7958
rect 2516 7290 2544 8026
rect 2608 7886 2636 8230
rect 2700 8022 2728 11070
rect 2872 11018 2924 11024
rect 2884 10538 2912 11018
rect 2976 10810 3004 22743
rect 3068 16182 3096 26823
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3056 16176 3108 16182
rect 3056 16118 3108 16124
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 3068 12986 3096 14758
rect 3148 14272 3200 14278
rect 3148 14214 3200 14220
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3160 12850 3188 14214
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3344 12646 3372 16934
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3896 14550 3924 14758
rect 4172 14550 4200 27390
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 13924 22114 13952 27520
rect 17224 26852 17276 26858
rect 17224 26794 17276 26800
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 13740 22086 13952 22114
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 10874 21448 10930 21457
rect 10874 21383 10930 21392
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 9678 18864 9734 18873
rect 9678 18799 9734 18808
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 9126 18048 9182 18057
rect 9126 17983 9182 17992
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 8022 16960 8078 16969
rect 8022 16895 8078 16904
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 7654 16008 7710 16017
rect 7564 15972 7616 15978
rect 7654 15943 7710 15952
rect 7564 15914 7616 15920
rect 4894 15464 4950 15473
rect 4894 15399 4950 15408
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 4264 14958 4292 15302
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4264 14618 4292 14894
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 3884 14544 3936 14550
rect 3884 14486 3936 14492
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3436 12782 3464 14214
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3422 12608 3478 12617
rect 3422 12543 3478 12552
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3160 11830 3188 12378
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3148 11824 3200 11830
rect 3148 11766 3200 11772
rect 3160 11218 3188 11766
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2872 10532 2924 10538
rect 2872 10474 2924 10480
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2884 10198 2912 10474
rect 2872 10192 2924 10198
rect 2778 10160 2834 10169
rect 2872 10134 2924 10140
rect 2778 10095 2780 10104
rect 2832 10095 2834 10104
rect 2780 10066 2832 10072
rect 2976 10062 3004 10474
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2884 8430 2912 9046
rect 2976 8974 3004 9386
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2688 8016 2740 8022
rect 2976 7993 3004 8910
rect 3068 8537 3096 11154
rect 3054 8528 3110 8537
rect 3054 8463 3110 8472
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 2688 7958 2740 7964
rect 2962 7984 3018 7993
rect 2962 7919 3018 7928
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2964 7812 3016 7818
rect 2964 7754 3016 7760
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2516 7262 2636 7290
rect 2608 7154 2636 7262
rect 2608 7126 2728 7154
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2240 5846 2268 6598
rect 2516 6458 2544 6666
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2608 6390 2636 6938
rect 2700 6474 2728 7126
rect 2700 6458 2820 6474
rect 2700 6452 2832 6458
rect 2700 6446 2780 6452
rect 2780 6394 2832 6400
rect 2596 6384 2648 6390
rect 2596 6326 2648 6332
rect 2502 6216 2558 6225
rect 2502 6151 2558 6160
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2228 5840 2280 5846
rect 2228 5782 2280 5788
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2136 3460 2188 3466
rect 2136 3402 2188 3408
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 1860 2984 1912 2990
rect 1858 2952 1860 2961
rect 1912 2952 1914 2961
rect 1858 2887 1914 2896
rect 1780 2774 1992 2802
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 1964 2553 1992 2774
rect 1950 2544 2006 2553
rect 2240 2514 2268 5306
rect 2424 4826 2452 5850
rect 2516 5710 2544 6151
rect 2884 6066 2912 7686
rect 2700 6038 2912 6066
rect 2700 5914 2728 6038
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2516 5098 2544 5646
rect 2504 5092 2556 5098
rect 2504 5034 2556 5040
rect 2700 5030 2728 5714
rect 2976 5370 3004 7754
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 3068 5250 3096 8366
rect 3252 6322 3280 12038
rect 3344 11898 3372 12242
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3344 10130 3372 10542
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3436 9625 3464 12543
rect 3528 12442 3556 14418
rect 4172 14006 4200 14486
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4448 14074 4476 14418
rect 4528 14340 4580 14346
rect 4528 14282 4580 14288
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4160 14000 4212 14006
rect 4160 13942 4212 13948
rect 3608 13728 3660 13734
rect 3608 13670 3660 13676
rect 3620 12850 3648 13670
rect 4172 13394 4200 13942
rect 4160 13388 4212 13394
rect 4212 13348 4292 13376
rect 4160 13330 4212 13336
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3620 12714 3648 12786
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3608 11008 3660 11014
rect 3608 10950 3660 10956
rect 3620 10606 3648 10950
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3698 10568 3754 10577
rect 3896 10538 3924 13126
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4172 12170 4200 12718
rect 4264 12306 4292 13348
rect 4448 12442 4476 14010
rect 4540 13870 4568 14282
rect 4710 13968 4766 13977
rect 4710 13903 4766 13912
rect 4528 13864 4580 13870
rect 4528 13806 4580 13812
rect 4724 13161 4752 13903
rect 4802 13288 4858 13297
rect 4802 13223 4858 13232
rect 4710 13152 4766 13161
rect 4710 13087 4766 13096
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3698 10503 3754 10512
rect 3884 10532 3936 10538
rect 3422 9616 3478 9625
rect 3422 9551 3478 9560
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 2976 5222 3096 5250
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2792 4162 2820 4966
rect 2608 4134 2820 4162
rect 2412 3664 2464 3670
rect 2412 3606 2464 3612
rect 2318 2680 2374 2689
rect 2424 2650 2452 3606
rect 2318 2615 2374 2624
rect 2412 2644 2464 2650
rect 2332 2582 2360 2615
rect 2412 2586 2464 2592
rect 2320 2576 2372 2582
rect 2320 2518 2372 2524
rect 1950 2479 2006 2488
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 2044 2100 2096 2106
rect 2044 2042 2096 2048
rect 2056 480 2084 2042
rect 2608 480 2636 4134
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2778 3768 2834 3777
rect 2778 3703 2834 3712
rect 2792 2854 2820 3703
rect 2884 3534 2912 3878
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2884 2650 2912 3470
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2976 1057 3004 5222
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 3068 2961 3096 4422
rect 3252 4010 3280 4558
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 3146 3768 3202 3777
rect 3252 3738 3280 3946
rect 3146 3703 3202 3712
rect 3240 3732 3292 3738
rect 3054 2952 3110 2961
rect 3054 2887 3110 2896
rect 2962 1048 3018 1057
rect 2962 983 3018 992
rect 3160 480 3188 3703
rect 3240 3674 3292 3680
rect 3252 3194 3280 3674
rect 3344 3670 3372 8774
rect 3436 5574 3464 9318
rect 3514 8392 3570 8401
rect 3514 8327 3570 8336
rect 3528 7546 3556 8327
rect 3712 8265 3740 10503
rect 3884 10474 3936 10480
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3698 8256 3754 8265
rect 3698 8191 3754 8200
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3528 6934 3556 7482
rect 3516 6928 3568 6934
rect 3516 6870 3568 6876
rect 3528 6322 3556 6870
rect 3620 6458 3648 7890
rect 3698 6896 3754 6905
rect 3698 6831 3754 6840
rect 3712 6730 3740 6831
rect 3700 6724 3752 6730
rect 3700 6666 3752 6672
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3528 5914 3556 6258
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3804 4758 3832 6598
rect 3896 5914 3924 8774
rect 3988 6730 4016 12038
rect 4264 11626 4292 12242
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4080 11082 4108 11562
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4066 10704 4122 10713
rect 4066 10639 4122 10648
rect 4080 9654 4108 10639
rect 4356 9654 4384 11290
rect 4528 11280 4580 11286
rect 4528 11222 4580 11228
rect 4540 10305 4568 11222
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4632 10810 4660 11086
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4526 10296 4582 10305
rect 4526 10231 4582 10240
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4080 8974 4108 9114
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4080 8566 4108 8910
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 4356 8362 4384 8978
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4250 7848 4306 7857
rect 4080 7002 4108 7822
rect 4250 7783 4306 7792
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 3988 6254 4016 6666
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 4264 5914 4292 7783
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4434 7440 4490 7449
rect 4434 7375 4436 7384
rect 4488 7375 4490 7384
rect 4436 7346 4488 7352
rect 3884 5908 3936 5914
rect 4252 5908 4304 5914
rect 3936 5868 4016 5896
rect 3884 5850 3936 5856
rect 3988 4808 4016 5868
rect 4252 5850 4304 5856
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4080 5370 4108 5714
rect 4264 5370 4292 5850
rect 4540 5681 4568 7686
rect 4526 5672 4582 5681
rect 4526 5607 4582 5616
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4252 5160 4304 5166
rect 4066 5128 4122 5137
rect 4252 5102 4304 5108
rect 4066 5063 4122 5072
rect 4080 5030 4108 5063
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4160 4820 4212 4826
rect 3988 4780 4160 4808
rect 4160 4762 4212 4768
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 4264 4570 4292 5102
rect 4172 4542 4292 4570
rect 4172 4486 4200 4542
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4080 3670 4108 3878
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 4172 3602 4200 4422
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3252 2446 3280 3130
rect 3422 3088 3478 3097
rect 3422 3023 3478 3032
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3436 1601 3464 3023
rect 3896 2922 3924 3470
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4356 2990 4384 3334
rect 4632 3194 4660 8570
rect 4710 8120 4766 8129
rect 4710 8055 4766 8064
rect 4724 7313 4752 8055
rect 4710 7304 4766 7313
rect 4710 7239 4766 7248
rect 4724 6254 4752 7239
rect 4816 7206 4844 13223
rect 4908 12594 4936 15399
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5736 14550 5764 14962
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 5724 14544 5776 14550
rect 5724 14486 5776 14492
rect 5736 14362 5764 14486
rect 5552 14334 5764 14362
rect 5552 14074 5580 14334
rect 6932 14249 6960 14758
rect 6918 14240 6974 14249
rect 5622 14172 5918 14192
rect 6918 14175 6974 14184
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 7116 13870 7144 14758
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 13870 7328 14214
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 5552 13530 5580 13806
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 6644 13456 6696 13462
rect 5998 13424 6054 13433
rect 5080 13388 5132 13394
rect 6644 13398 6696 13404
rect 5998 13359 6054 13368
rect 5080 13330 5132 13336
rect 5092 12850 5120 13330
rect 6012 13161 6040 13359
rect 5998 13152 6054 13161
rect 5622 13084 5918 13104
rect 5998 13087 6054 13096
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6656 12986 6684 13398
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6734 12880 6790 12889
rect 5080 12844 5132 12850
rect 5132 12804 5212 12832
rect 6734 12815 6790 12824
rect 5080 12786 5132 12792
rect 4986 12744 5042 12753
rect 4986 12679 4988 12688
rect 5040 12679 5042 12688
rect 4988 12650 5040 12656
rect 4908 12566 5120 12594
rect 5092 11098 5120 12566
rect 5184 12238 5212 12804
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5184 12102 5212 12174
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5184 11898 5212 12038
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5552 11626 5580 12174
rect 6000 12164 6052 12170
rect 6000 12106 6052 12112
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 5552 11529 5580 11562
rect 6012 11558 6040 12106
rect 6196 11558 6224 12242
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6000 11552 6052 11558
rect 5538 11520 5594 11529
rect 6184 11552 6236 11558
rect 6000 11494 6052 11500
rect 6182 11520 6184 11529
rect 6236 11520 6238 11529
rect 5538 11455 5594 11464
rect 6182 11455 6238 11464
rect 6288 11286 6316 12038
rect 6472 11898 6500 12174
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6092 11144 6144 11150
rect 5092 11070 5212 11098
rect 6144 11092 6224 11098
rect 6092 11086 6224 11092
rect 5184 11014 5212 11070
rect 6000 11076 6052 11082
rect 6104 11070 6224 11086
rect 6000 11018 6052 11024
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5184 10470 5212 10950
rect 5172 10464 5224 10470
rect 5092 10424 5172 10452
rect 4894 7440 4950 7449
rect 4894 7375 4950 7384
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4908 6798 4936 7375
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4816 6390 4844 6734
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4620 3188 4672 3194
rect 4540 3148 4620 3176
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 3884 2916 3936 2922
rect 3884 2858 3936 2864
rect 3896 2650 3924 2858
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3422 1592 3478 1601
rect 3422 1527 3478 1536
rect 3698 1320 3754 1329
rect 3698 1255 3754 1264
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 2042 0 2098 480
rect 2594 0 2650 480
rect 3146 0 3202 480
rect 3712 377 3740 1255
rect 4540 610 4568 3148
rect 4620 3130 4672 3136
rect 4816 2666 4844 6326
rect 4908 6322 4936 6734
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4908 5846 4936 6258
rect 4896 5840 4948 5846
rect 4896 5782 4948 5788
rect 5092 3913 5120 10424
rect 5172 10406 5224 10412
rect 5356 10192 5408 10198
rect 5262 10160 5318 10169
rect 5356 10134 5408 10140
rect 5262 10095 5318 10104
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5184 9586 5212 9862
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5276 8634 5304 10095
rect 5368 9382 5396 10134
rect 5460 9518 5488 10950
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6012 10674 6040 11018
rect 6092 11008 6144 11014
rect 6090 10976 6092 10985
rect 6144 10976 6146 10985
rect 6090 10911 6146 10920
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5540 10600 5592 10606
rect 5538 10568 5540 10577
rect 5592 10568 5594 10577
rect 5538 10503 5594 10512
rect 6012 10130 6040 10610
rect 6196 10470 6224 11070
rect 6472 10810 6500 11154
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6196 10198 6224 10406
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6012 9926 6040 10066
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 6012 9382 6040 9862
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5368 8566 5396 9318
rect 5460 8838 5488 9318
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5460 8498 5488 8774
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5368 8090 5396 8366
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5170 7712 5226 7721
rect 5170 7647 5226 7656
rect 5184 7546 5212 7647
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5172 6928 5224 6934
rect 5172 6870 5224 6876
rect 5184 5778 5212 6870
rect 5460 6390 5488 8230
rect 5552 7886 5580 8502
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5552 7528 5580 7822
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5552 7500 5764 7528
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5644 7002 5672 7346
rect 5736 7342 5764 7500
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5920 7002 5948 7210
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5264 5636 5316 5642
rect 5264 5578 5316 5584
rect 5276 5098 5304 5578
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5078 3904 5134 3913
rect 5078 3839 5134 3848
rect 4816 2638 4936 2666
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4632 2009 4660 2450
rect 4618 2000 4674 2009
rect 4618 1935 4674 1944
rect 3792 604 3844 610
rect 3792 546 3844 552
rect 4528 604 4580 610
rect 4528 546 4580 552
rect 3804 480 3832 546
rect 4344 536 4396 542
rect 4344 480 4396 484
rect 4908 480 4936 2638
rect 5184 542 5212 4966
rect 5276 4690 5304 5034
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5276 3738 5304 4626
rect 5368 4622 5396 5306
rect 5448 4820 5500 4826
rect 5552 4808 5580 5850
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6012 4865 6040 8774
rect 6196 8362 6224 9046
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6104 7546 6132 7890
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6104 6458 6132 6734
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6090 6080 6146 6089
rect 6090 6015 6146 6024
rect 6104 5710 6132 6015
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6104 5030 6132 5646
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 5500 4780 5580 4808
rect 5998 4856 6054 4865
rect 5998 4791 6054 4800
rect 5448 4762 5500 4768
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5368 4214 5396 4558
rect 5448 4480 5500 4486
rect 5446 4448 5448 4457
rect 5500 4448 5502 4457
rect 5446 4383 5502 4392
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 5552 3738 5580 4626
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6012 4078 6040 4791
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6104 3777 6132 3878
rect 6090 3768 6146 3777
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5540 3732 5592 3738
rect 6090 3703 6146 3712
rect 5540 3674 5592 3680
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5354 3088 5410 3097
rect 5354 3023 5410 3032
rect 5368 2825 5396 3023
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5552 2938 5580 3334
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5630 2952 5686 2961
rect 5354 2816 5410 2825
rect 5354 2751 5410 2760
rect 5460 2650 5488 2926
rect 5552 2910 5630 2938
rect 5630 2887 5686 2896
rect 6092 2916 6144 2922
rect 5644 2854 5672 2887
rect 6092 2858 6144 2864
rect 5632 2848 5684 2854
rect 5538 2816 5594 2825
rect 5632 2790 5684 2796
rect 5538 2751 5594 2760
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5172 536 5224 542
rect 3698 368 3754 377
rect 3698 303 3754 312
rect 3790 0 3846 480
rect 4342 0 4398 480
rect 4894 0 4950 480
rect 5172 478 5224 484
rect 5552 480 5580 2751
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6104 480 6132 2858
rect 6196 2825 6224 8298
rect 6288 7274 6316 9318
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6288 6458 6316 6802
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6380 5914 6408 8774
rect 6472 6798 6500 10746
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6564 6610 6592 11562
rect 6656 11354 6684 12038
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6472 6582 6592 6610
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6288 4468 6316 5782
rect 6366 5400 6422 5409
rect 6366 5335 6422 5344
rect 6380 4826 6408 5335
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6368 4480 6420 4486
rect 6288 4440 6368 4468
rect 6368 4422 6420 4428
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6380 3942 6408 4014
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6182 2816 6238 2825
rect 6182 2751 6238 2760
rect 6380 2106 6408 3878
rect 6472 2922 6500 6582
rect 6748 5846 6776 12815
rect 7116 12374 7144 13806
rect 7300 13530 7328 13806
rect 7576 13530 7604 15914
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7300 13433 7328 13466
rect 7286 13424 7342 13433
rect 7286 13359 7342 13368
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7576 12986 7604 13330
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7104 12368 7156 12374
rect 7104 12310 7156 12316
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 7024 11354 7052 12174
rect 7116 11694 7144 12310
rect 7392 12102 7420 12718
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 7300 10606 7328 11630
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 7194 9888 7250 9897
rect 6932 8344 6960 9862
rect 7194 9823 7250 9832
rect 7208 9178 7236 9823
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7116 8498 7144 8774
rect 7208 8634 7236 8774
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 6840 8316 6960 8344
rect 6840 7002 6868 8316
rect 7300 7936 7328 8502
rect 7208 7908 7328 7936
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 7449 6960 7686
rect 6918 7440 6974 7449
rect 6918 7375 6974 7384
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6932 6662 6960 7210
rect 7116 6730 7144 7210
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 7010 6624 7066 6633
rect 7010 6559 7066 6568
rect 6736 5840 6788 5846
rect 6736 5782 6788 5788
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6826 5672 6882 5681
rect 6550 5264 6606 5273
rect 6550 5199 6606 5208
rect 6564 4758 6592 5199
rect 6642 4992 6698 5001
rect 6642 4927 6698 4936
rect 6656 4826 6684 4927
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6552 4752 6604 4758
rect 6552 4694 6604 4700
rect 6564 4282 6592 4694
rect 6656 4622 6684 4762
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6564 2922 6592 3538
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 6564 2310 6592 2858
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6368 2100 6420 2106
rect 6368 2042 6420 2048
rect 6656 480 6684 4422
rect 6748 4214 6776 5646
rect 6826 5607 6882 5616
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6840 3942 6868 5607
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6828 3936 6880 3942
rect 6734 3904 6790 3913
rect 6828 3878 6880 3884
rect 6734 3839 6790 3848
rect 6748 3534 6776 3839
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6748 2514 6776 3470
rect 6828 3188 6880 3194
rect 6932 3176 6960 5510
rect 7024 4486 7052 6559
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7116 5370 7144 5646
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 7116 5166 7144 5306
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7208 4758 7236 7908
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7196 4752 7248 4758
rect 7196 4694 7248 4700
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7208 3777 7236 3878
rect 7194 3768 7250 3777
rect 7194 3703 7250 3712
rect 6880 3148 6960 3176
rect 6828 3130 6880 3136
rect 6932 2689 6960 3148
rect 6918 2680 6974 2689
rect 6918 2615 6974 2624
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6748 2281 6776 2450
rect 6734 2272 6790 2281
rect 6734 2207 6790 2216
rect 7300 480 7328 7754
rect 7392 4049 7420 12038
rect 7484 8566 7512 12650
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7576 11354 7604 11630
rect 7668 11354 7696 15943
rect 7838 15600 7894 15609
rect 7838 15535 7894 15544
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 7760 12442 7788 13398
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7746 12336 7802 12345
rect 7746 12271 7802 12280
rect 7760 12238 7788 12271
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7562 10840 7618 10849
rect 7562 10775 7618 10784
rect 7576 10266 7604 10775
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7668 10470 7696 10542
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7576 9382 7604 10066
rect 7668 9518 7696 10406
rect 7748 9988 7800 9994
rect 7748 9930 7800 9936
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7472 8560 7524 8566
rect 7472 8502 7524 8508
rect 7576 8401 7604 9318
rect 7562 8392 7618 8401
rect 7484 8350 7562 8378
rect 7484 5817 7512 8350
rect 7562 8327 7618 8336
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7576 7750 7604 8230
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7576 6304 7604 7686
rect 7668 7342 7696 9454
rect 7760 8974 7788 9930
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7760 8090 7788 8910
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7746 7712 7802 7721
rect 7746 7647 7802 7656
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7760 7177 7788 7647
rect 7746 7168 7802 7177
rect 7746 7103 7802 7112
rect 7576 6276 7788 6304
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7470 5808 7526 5817
rect 7470 5743 7526 5752
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 7484 4214 7512 4490
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7576 4146 7604 6122
rect 7760 5778 7788 6276
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7378 4040 7434 4049
rect 7378 3975 7434 3984
rect 7656 3528 7708 3534
rect 7654 3496 7656 3505
rect 7708 3496 7710 3505
rect 7380 3460 7432 3466
rect 7654 3431 7710 3440
rect 7380 3402 7432 3408
rect 7392 3058 7420 3402
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7484 2417 7512 2926
rect 7668 2582 7696 3431
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 7470 2408 7526 2417
rect 7470 2343 7526 2352
rect 7760 610 7788 5714
rect 7748 604 7800 610
rect 7748 546 7800 552
rect 7852 480 7880 15535
rect 8036 15434 8064 16895
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 8404 15910 8432 16050
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8668 15904 8720 15910
rect 8668 15846 8720 15852
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8024 15428 8076 15434
rect 8024 15370 8076 15376
rect 8312 15162 8340 15438
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8312 15065 8340 15098
rect 8298 15056 8354 15065
rect 8298 14991 8354 15000
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8116 13796 8168 13802
rect 8116 13738 8168 13744
rect 8128 13326 8156 13738
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7944 11744 7972 12582
rect 8128 12442 8156 13262
rect 8220 12782 8248 14350
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8116 12436 8168 12442
rect 8116 12378 8168 12384
rect 8116 12164 8168 12170
rect 8116 12106 8168 12112
rect 7944 11716 8064 11744
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7944 7818 7972 11562
rect 8036 11132 8064 11716
rect 8128 11286 8156 12106
rect 8404 12102 8432 15846
rect 8680 15706 8708 15846
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 8576 14884 8628 14890
rect 8576 14826 8628 14832
rect 8588 14346 8616 14826
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 8588 13734 8616 14282
rect 8680 14278 8708 15506
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8588 13190 8616 13670
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8588 12850 8616 13126
rect 8576 12844 8628 12850
rect 8496 12804 8576 12832
rect 8496 12238 8524 12804
rect 8576 12786 8628 12792
rect 8576 12640 8628 12646
rect 8680 12617 8708 14214
rect 8850 13016 8906 13025
rect 8850 12951 8906 12960
rect 8576 12582 8628 12588
rect 8666 12608 8722 12617
rect 8588 12481 8616 12582
rect 8666 12543 8722 12552
rect 8574 12472 8630 12481
rect 8574 12407 8630 12416
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8390 11792 8446 11801
rect 8390 11727 8392 11736
rect 8444 11727 8446 11736
rect 8392 11698 8444 11704
rect 8864 11626 8892 12951
rect 9048 11898 9076 15846
rect 9140 13530 9168 17983
rect 9220 16448 9272 16454
rect 9220 16390 9272 16396
rect 9232 15910 9260 16390
rect 9692 16250 9720 18799
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 10152 16998 10180 17138
rect 10796 17134 10824 17682
rect 10784 17128 10836 17134
rect 10690 17096 10746 17105
rect 10784 17070 10836 17076
rect 10690 17031 10746 17040
rect 10704 16998 10732 17031
rect 10140 16992 10192 16998
rect 10138 16960 10140 16969
rect 10692 16992 10744 16998
rect 10192 16960 10194 16969
rect 10692 16934 10744 16940
rect 10138 16895 10194 16904
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10796 16794 10824 17070
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9784 16182 9812 16594
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 9772 16176 9824 16182
rect 9772 16118 9824 16124
rect 10138 16144 10194 16153
rect 10336 16114 10364 16390
rect 10796 16114 10824 16730
rect 10138 16079 10194 16088
rect 10324 16108 10376 16114
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9140 12986 9168 13466
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9048 11694 9076 11834
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 8852 11620 8904 11626
rect 8852 11562 8904 11568
rect 8300 11552 8352 11558
rect 9232 11529 9260 15846
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9692 15162 9720 15438
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9692 14414 9720 14826
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9968 14482 9996 14758
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9692 14074 9720 14350
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9968 13870 9996 14418
rect 10046 14104 10102 14113
rect 10046 14039 10102 14048
rect 9956 13864 10008 13870
rect 9310 13832 9366 13841
rect 9956 13806 10008 13812
rect 9310 13767 9366 13776
rect 9324 13394 9352 13767
rect 9494 13424 9550 13433
rect 9312 13388 9364 13394
rect 9494 13359 9550 13368
rect 9312 13330 9364 13336
rect 9324 12986 9352 13330
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9312 11552 9364 11558
rect 8300 11494 8352 11500
rect 9218 11520 9274 11529
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 8036 11104 8156 11132
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8036 8498 8064 8978
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 8128 8265 8156 11104
rect 8208 10600 8260 10606
rect 8312 10588 8340 11494
rect 9312 11494 9364 11500
rect 9218 11455 9274 11464
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8260 10560 8340 10588
rect 8208 10542 8260 10548
rect 8220 10062 8248 10542
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8206 9344 8262 9353
rect 8206 9279 8262 9288
rect 8220 8945 8248 9279
rect 8404 9042 8432 10066
rect 8496 9518 8524 10746
rect 8680 10266 8708 11086
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8956 10810 8984 10950
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 8758 10432 8814 10441
rect 8758 10367 8814 10376
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8680 9722 8708 10202
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8206 8936 8262 8945
rect 8206 8871 8262 8880
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8114 8256 8170 8265
rect 8114 8191 8170 8200
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 8036 7449 8064 7686
rect 8022 7440 8078 7449
rect 8022 7375 8078 7384
rect 8114 7032 8170 7041
rect 8312 7002 8340 8842
rect 8300 6996 8352 7002
rect 8114 6967 8170 6976
rect 8128 6934 8156 6967
rect 8220 6956 8300 6984
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8036 6118 8064 6190
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 8036 5098 8064 6054
rect 8128 5846 8156 6598
rect 8220 5914 8248 6956
rect 8300 6938 8352 6944
rect 8404 6361 8432 8978
rect 8588 8974 8616 9386
rect 8680 9178 8708 9658
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8588 8566 8616 8910
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8588 8430 8616 8502
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8680 8362 8708 9114
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 8680 7274 8708 7958
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8496 6458 8524 6734
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8390 6352 8446 6361
rect 8390 6287 8446 6296
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8128 5658 8156 5782
rect 8128 5630 8248 5658
rect 8404 5642 8432 6122
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8220 5522 8248 5630
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8220 5494 8340 5522
rect 8312 5302 8340 5494
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 7930 4856 7986 4865
rect 7930 4791 7932 4800
rect 7984 4791 7986 4800
rect 7932 4762 7984 4768
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 7930 4584 7986 4593
rect 7930 4519 7986 4528
rect 7944 4078 7972 4519
rect 8036 4457 8064 4694
rect 8220 4622 8248 4966
rect 8298 4720 8354 4729
rect 8298 4655 8300 4664
rect 8352 4655 8354 4664
rect 8300 4626 8352 4632
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8022 4448 8078 4457
rect 8022 4383 8078 4392
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7930 3904 7986 3913
rect 7930 3839 7986 3848
rect 7944 3194 7972 3839
rect 8036 3738 8064 4383
rect 8312 4026 8340 4626
rect 8220 3998 8340 4026
rect 8220 3942 8248 3998
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 8220 3398 8248 3878
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 7944 2854 7972 3130
rect 8220 3097 8248 3334
rect 8404 3233 8432 3878
rect 8390 3224 8446 3233
rect 8496 3194 8524 5102
rect 8588 5030 8616 5646
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8680 3777 8708 7210
rect 8772 6730 8800 10367
rect 8944 10192 8996 10198
rect 8942 10160 8944 10169
rect 8996 10160 8998 10169
rect 8942 10095 8998 10104
rect 9232 9636 9260 11455
rect 9324 11354 9352 11494
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9310 10976 9366 10985
rect 9310 10911 9366 10920
rect 9324 10266 9352 10911
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9416 9761 9444 13126
rect 9508 12238 9536 13359
rect 10060 13274 10088 14039
rect 9968 13246 10088 13274
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9588 12436 9640 12442
rect 9692 12424 9720 12582
rect 9640 12396 9720 12424
rect 9588 12378 9640 12384
rect 9784 12345 9812 13126
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9770 12336 9826 12345
rect 9876 12306 9904 12650
rect 9770 12271 9826 12280
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9496 12096 9548 12102
rect 9494 12064 9496 12073
rect 9548 12064 9550 12073
rect 9494 11999 9550 12008
rect 9586 11928 9642 11937
rect 9586 11863 9588 11872
rect 9640 11863 9642 11872
rect 9772 11892 9824 11898
rect 9588 11834 9640 11840
rect 9772 11834 9824 11840
rect 9588 11756 9640 11762
rect 9784 11744 9812 11834
rect 9640 11716 9812 11744
rect 9588 11698 9640 11704
rect 9494 11656 9550 11665
rect 9494 11591 9550 11600
rect 9508 11558 9536 11591
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9784 11286 9812 11494
rect 9772 11280 9824 11286
rect 9772 11222 9824 11228
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9508 10452 9536 11154
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9600 10588 9628 11018
rect 9680 10600 9732 10606
rect 9600 10560 9680 10588
rect 9680 10542 9732 10548
rect 9588 10464 9640 10470
rect 9508 10424 9588 10452
rect 9588 10406 9640 10412
rect 9600 10169 9628 10406
rect 9586 10160 9642 10169
rect 9586 10095 9642 10104
rect 9402 9752 9458 9761
rect 9402 9687 9458 9696
rect 9140 9608 9260 9636
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8864 6662 8892 7822
rect 8956 7206 8984 7890
rect 9140 7886 9168 9608
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9232 8090 9260 9318
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9404 8832 9456 8838
rect 9600 8809 9628 8978
rect 9404 8774 9456 8780
rect 9586 8800 9642 8809
rect 9416 8673 9444 8774
rect 9586 8735 9642 8744
rect 9402 8664 9458 8673
rect 9402 8599 9458 8608
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8864 6118 8892 6598
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8666 3768 8722 3777
rect 8666 3703 8722 3712
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8390 3159 8446 3168
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8206 3088 8262 3097
rect 8206 3023 8262 3032
rect 8496 2990 8524 3130
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 8496 2650 8524 2926
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 8312 2009 8340 2314
rect 8588 2122 8616 3470
rect 8666 2136 8722 2145
rect 8588 2094 8666 2122
rect 8666 2071 8722 2080
rect 8298 2000 8354 2009
rect 8772 1986 8800 5646
rect 8864 4486 8892 6054
rect 8956 4593 8984 7142
rect 9048 5273 9076 7686
rect 9034 5264 9090 5273
rect 9034 5199 9090 5208
rect 9036 5024 9088 5030
rect 9140 5001 9168 7686
rect 9218 7576 9274 7585
rect 9218 7511 9274 7520
rect 9232 7274 9260 7511
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9232 5681 9260 6598
rect 9218 5672 9274 5681
rect 9218 5607 9274 5616
rect 9220 5296 9272 5302
rect 9218 5264 9220 5273
rect 9272 5264 9274 5273
rect 9218 5199 9274 5208
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9036 4966 9088 4972
rect 9126 4992 9182 5001
rect 9048 4706 9076 4966
rect 9126 4927 9182 4936
rect 9232 4826 9260 5102
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9048 4678 9260 4706
rect 8942 4584 8998 4593
rect 8942 4519 8998 4528
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9140 4214 9168 4422
rect 9128 4208 9180 4214
rect 9128 4150 9180 4156
rect 9034 3632 9090 3641
rect 9034 3567 9090 3576
rect 9048 2990 9076 3567
rect 9140 3505 9168 4150
rect 9126 3496 9182 3505
rect 9126 3431 9182 3440
rect 9036 2984 9088 2990
rect 9232 2961 9260 4678
rect 9324 2990 9352 8366
rect 9402 8120 9458 8129
rect 9692 8090 9720 10542
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9784 8673 9812 10406
rect 9876 10305 9904 12242
rect 9862 10296 9918 10305
rect 9862 10231 9918 10240
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9876 9926 9904 10134
rect 9864 9920 9916 9926
rect 9862 9888 9864 9897
rect 9916 9888 9918 9897
rect 9862 9823 9918 9832
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9770 8664 9826 8673
rect 9770 8599 9826 8608
rect 9402 8055 9458 8064
rect 9588 8084 9640 8090
rect 9416 6497 9444 8055
rect 9588 8026 9640 8032
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9402 6488 9458 6497
rect 9402 6423 9458 6432
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5098 9444 5510
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9404 4072 9456 4078
rect 9508 4060 9536 7822
rect 9600 6746 9628 8026
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9692 6905 9720 7278
rect 9784 7177 9812 7346
rect 9770 7168 9826 7177
rect 9770 7103 9826 7112
rect 9876 7041 9904 8774
rect 9862 7032 9918 7041
rect 9862 6967 9918 6976
rect 9678 6896 9734 6905
rect 9678 6831 9734 6840
rect 9772 6792 9824 6798
rect 9770 6760 9772 6769
rect 9824 6760 9826 6769
rect 9600 6718 9720 6746
rect 9692 5710 9720 6718
rect 9770 6695 9826 6704
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9784 6089 9812 6326
rect 9770 6080 9826 6089
rect 9770 6015 9826 6024
rect 9876 5914 9904 6967
rect 9968 6866 9996 13246
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 10060 12102 10088 12582
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10060 11830 10088 12038
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 10060 11082 10088 11630
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 10152 10146 10180 16079
rect 10324 16050 10376 16056
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10244 14890 10272 15438
rect 10232 14884 10284 14890
rect 10232 14826 10284 14832
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14074 10732 16050
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10796 15094 10824 15914
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10888 14906 10916 21383
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13280 19718 13308 20402
rect 13740 20330 13768 22086
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 14740 20256 14792 20262
rect 14740 20198 14792 20204
rect 13268 19712 13320 19718
rect 13268 19654 13320 19660
rect 11702 19272 11758 19281
rect 11702 19207 11758 19216
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11072 17678 11100 18022
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 11072 17082 11100 17614
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 11348 17202 11376 17478
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11072 17054 11284 17082
rect 11256 16998 11284 17054
rect 11060 16992 11112 16998
rect 11058 16960 11060 16969
rect 11244 16992 11296 16998
rect 11112 16960 11114 16969
rect 11244 16934 11296 16940
rect 11058 16895 11114 16904
rect 11256 16454 11284 16934
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11256 15910 11284 16390
rect 11336 16176 11388 16182
rect 11336 16118 11388 16124
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 10966 15056 11022 15065
rect 10966 14991 11022 15000
rect 10796 14878 10916 14906
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10690 13560 10746 13569
rect 10690 13495 10746 13504
rect 10230 13424 10286 13433
rect 10704 13394 10732 13495
rect 10230 13359 10286 13368
rect 10692 13388 10744 13394
rect 10244 13326 10272 13359
rect 10692 13330 10744 13336
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10244 12850 10272 13262
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10428 11626 10456 12174
rect 10690 12064 10746 12073
rect 10690 11999 10746 12008
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10704 11286 10732 11999
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10232 11076 10284 11082
rect 10232 11018 10284 11024
rect 10244 10985 10272 11018
rect 10692 11008 10744 11014
rect 10230 10976 10286 10985
rect 10692 10950 10744 10956
rect 10230 10911 10286 10920
rect 10704 10470 10732 10950
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10690 10296 10746 10305
rect 10690 10231 10746 10240
rect 10060 10118 10180 10146
rect 10060 7834 10088 10118
rect 10140 10056 10192 10062
rect 10704 10033 10732 10231
rect 10140 9998 10192 10004
rect 10690 10024 10746 10033
rect 10152 9489 10180 9998
rect 10690 9959 10746 9968
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10138 9480 10194 9489
rect 10138 9415 10194 9424
rect 10140 9376 10192 9382
rect 10138 9344 10140 9353
rect 10612 9364 10640 9658
rect 10704 9586 10732 9862
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10192 9344 10194 9353
rect 10612 9336 10732 9364
rect 10138 9279 10194 9288
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10414 8936 10470 8945
rect 10244 8498 10272 8910
rect 10414 8871 10470 8880
rect 10428 8838 10456 8871
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10520 8634 10548 8978
rect 10704 8945 10732 9336
rect 10690 8936 10746 8945
rect 10690 8871 10746 8880
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10506 7984 10562 7993
rect 10506 7919 10508 7928
rect 10560 7919 10562 7928
rect 10508 7890 10560 7896
rect 10060 7806 10180 7834
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10060 6905 10088 7686
rect 10046 6896 10102 6905
rect 9956 6860 10008 6866
rect 10046 6831 10102 6840
rect 9956 6802 10008 6808
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9968 4690 9996 6802
rect 10046 6080 10102 6089
rect 10046 6015 10102 6024
rect 10060 5778 10088 6015
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 10060 4486 10088 5714
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 10152 4162 10180 7806
rect 10520 7410 10548 7890
rect 10704 7886 10732 8570
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10612 7342 10640 7822
rect 10704 7478 10732 7822
rect 10796 7546 10824 14878
rect 10980 14385 11008 14991
rect 11072 14618 11100 15574
rect 11256 15570 11284 15846
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11348 15366 11376 16118
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 11348 15026 11376 15302
rect 11716 15026 11744 19207
rect 13280 19174 13308 19654
rect 14096 19236 14148 19242
rect 14096 19178 14148 19184
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 12438 18728 12494 18737
rect 12438 18663 12440 18672
rect 12492 18663 12494 18672
rect 12440 18634 12492 18640
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12360 18170 12388 18566
rect 12820 18426 12848 18770
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 12360 18142 12480 18170
rect 12452 17338 12480 18142
rect 12716 18148 12768 18154
rect 12716 18090 12768 18096
rect 12728 17610 12756 18090
rect 12820 17882 12848 18362
rect 13096 18086 13124 18702
rect 13280 18222 13308 19110
rect 14004 18760 14056 18766
rect 14004 18702 14056 18708
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 14016 17882 14044 18702
rect 14108 18630 14136 19178
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14108 18086 14136 18566
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 13266 17232 13322 17241
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 12532 17196 12584 17202
rect 13266 17167 13322 17176
rect 12532 17138 12584 17144
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 10966 14376 11022 14385
rect 11072 14346 11100 14554
rect 10966 14311 11022 14320
rect 11060 14340 11112 14346
rect 10980 14226 11008 14311
rect 11060 14282 11112 14288
rect 10888 14198 11008 14226
rect 10888 12374 10916 14198
rect 11072 14074 11100 14282
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10966 13968 11022 13977
rect 10966 13903 10968 13912
rect 11020 13903 11022 13912
rect 11060 13932 11112 13938
rect 10968 13874 11020 13880
rect 11060 13874 11112 13880
rect 11072 13818 11100 13874
rect 10980 13790 11100 13818
rect 10980 13530 11008 13790
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 11152 13456 11204 13462
rect 11152 13398 11204 13404
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 10980 12617 11008 13330
rect 11164 13025 11192 13398
rect 11150 13016 11206 13025
rect 11150 12951 11152 12960
rect 11204 12951 11206 12960
rect 11152 12922 11204 12928
rect 11256 12714 11284 14758
rect 11348 14618 11376 14962
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11348 13938 11376 14554
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 11426 13696 11482 13705
rect 11426 13631 11482 13640
rect 11334 13288 11390 13297
rect 11334 13223 11390 13232
rect 11348 13190 11376 13223
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11348 12782 11376 13126
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11336 12640 11388 12646
rect 10966 12608 11022 12617
rect 11336 12582 11388 12588
rect 10966 12543 11022 12552
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 11058 12336 11114 12345
rect 10888 11558 10916 12310
rect 10968 12300 11020 12306
rect 11058 12271 11114 12280
rect 10968 12242 11020 12248
rect 10980 12073 11008 12242
rect 10966 12064 11022 12073
rect 10966 11999 11022 12008
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10980 11370 11008 11766
rect 10888 11342 11008 11370
rect 10888 11257 10916 11342
rect 11072 11286 11100 12271
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 11060 11280 11112 11286
rect 10874 11248 10930 11257
rect 11060 11222 11112 11228
rect 10874 11183 10930 11192
rect 10888 9722 10916 11183
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10888 7818 10916 9522
rect 10980 9160 11008 10542
rect 11072 10130 11100 11222
rect 11164 11200 11192 11562
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11256 11354 11284 11494
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11244 11212 11296 11218
rect 11164 11172 11244 11200
rect 11244 11154 11296 11160
rect 11256 10470 11284 11154
rect 11244 10464 11296 10470
rect 11150 10432 11206 10441
rect 11244 10406 11296 10412
rect 11150 10367 11206 10376
rect 11164 10266 11192 10367
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 11060 9172 11112 9178
rect 10980 9132 11060 9160
rect 11060 9114 11112 9120
rect 10966 8936 11022 8945
rect 10966 8871 11022 8880
rect 10980 8838 11008 8871
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10692 7472 10744 7478
rect 10692 7414 10744 7420
rect 10600 7336 10652 7342
rect 10652 7284 10732 7290
rect 10600 7278 10732 7284
rect 10612 7262 10732 7278
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10704 6458 10732 7262
rect 10888 6866 10916 7754
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 10980 7041 11008 7210
rect 10966 7032 11022 7041
rect 11072 7002 11100 8434
rect 11164 8401 11192 9590
rect 11256 8498 11284 10406
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11150 8392 11206 8401
rect 11150 8327 11206 8336
rect 11164 7342 11192 8327
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11256 8090 11284 8230
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11256 7410 11284 7686
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11256 7002 11284 7346
rect 10966 6967 11022 6976
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10692 6112 10744 6118
rect 10796 6089 10824 6190
rect 10692 6054 10744 6060
rect 10782 6080 10838 6089
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9968 4134 10180 4162
rect 9508 4032 9720 4060
rect 9404 4014 9456 4020
rect 9312 2984 9364 2990
rect 9036 2926 9088 2932
rect 9218 2952 9274 2961
rect 9312 2926 9364 2932
rect 9218 2887 9274 2896
rect 8298 1935 8354 1944
rect 8404 1958 8800 1986
rect 8404 480 8432 1958
rect 9416 1465 9444 4014
rect 9588 3392 9640 3398
rect 9692 3369 9720 4032
rect 9770 4040 9826 4049
rect 9770 3975 9826 3984
rect 9588 3334 9640 3340
rect 9678 3360 9734 3369
rect 9600 3074 9628 3334
rect 9678 3295 9734 3304
rect 9678 3088 9734 3097
rect 9600 3046 9678 3074
rect 9678 3023 9734 3032
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9402 1456 9458 1465
rect 9402 1391 9458 1400
rect 9036 604 9088 610
rect 9036 546 9088 552
rect 9048 480 9076 546
rect 9600 480 9628 2926
rect 9692 2582 9720 3023
rect 9784 2650 9812 3975
rect 9876 3482 9904 4082
rect 9968 3670 9996 4134
rect 10244 4026 10272 4218
rect 10704 4078 10732 6054
rect 10782 6015 10838 6024
rect 10888 5914 10916 6802
rect 11072 6746 11100 6938
rect 10980 6718 11100 6746
rect 10980 6390 11008 6718
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10796 5001 10824 5646
rect 10888 5370 10916 5714
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10980 5216 11008 6326
rect 11072 6118 11100 6598
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 10888 5188 11008 5216
rect 10782 4992 10838 5001
rect 10782 4927 10838 4936
rect 10796 4826 10824 4927
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10888 4690 10916 5188
rect 11072 5148 11100 6054
rect 10980 5120 11100 5148
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10152 3998 10272 4026
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10060 3738 10088 3878
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9876 3454 9996 3482
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9772 2372 9824 2378
rect 9772 2314 9824 2320
rect 9784 2281 9812 2314
rect 9770 2272 9826 2281
rect 9770 2207 9826 2216
rect 9876 1873 9904 3334
rect 9968 3126 9996 3454
rect 10046 3360 10102 3369
rect 10046 3295 10102 3304
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 9968 2514 9996 3062
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 9862 1864 9918 1873
rect 9862 1799 9918 1808
rect 10060 1170 10088 3295
rect 10152 2650 10180 3998
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10704 3738 10732 4014
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10796 3618 10824 4490
rect 10888 4214 10916 4626
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10704 3590 10824 3618
rect 10888 3602 10916 4150
rect 10876 3596 10928 3602
rect 10230 3496 10286 3505
rect 10230 3431 10286 3440
rect 10244 3194 10272 3431
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 10704 1737 10732 3590
rect 10876 3538 10928 3544
rect 10888 3194 10916 3538
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10888 3058 10916 3130
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10888 2446 10916 2994
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 10874 2000 10930 2009
rect 10980 1986 11008 5120
rect 11256 4758 11284 6938
rect 11348 5914 11376 12582
rect 11440 11762 11468 13631
rect 11808 12442 11836 17138
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12176 15910 12204 16526
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12176 15609 12204 15846
rect 12162 15600 12218 15609
rect 12162 15535 12218 15544
rect 12268 15502 12296 16934
rect 12544 16794 12572 17138
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12714 16688 12770 16697
rect 12714 16623 12770 16632
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11808 11937 11836 12378
rect 11794 11928 11850 11937
rect 11794 11863 11850 11872
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11808 10742 11836 11494
rect 11796 10736 11848 10742
rect 11702 10704 11758 10713
rect 11796 10678 11848 10684
rect 11702 10639 11704 10648
rect 11756 10639 11758 10648
rect 11704 10610 11756 10616
rect 11808 10266 11836 10678
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11624 9382 11652 9998
rect 11702 9752 11758 9761
rect 11702 9687 11758 9696
rect 11612 9376 11664 9382
rect 11426 9344 11482 9353
rect 11612 9318 11664 9324
rect 11426 9279 11482 9288
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 4282 11100 4422
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11256 4214 11284 4694
rect 11244 4208 11296 4214
rect 11244 4150 11296 4156
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 11150 3632 11206 3641
rect 11072 2650 11100 3606
rect 11150 3567 11206 3576
rect 11164 3398 11192 3567
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11348 2990 11376 5850
rect 11440 5409 11468 9279
rect 11518 8528 11574 8537
rect 11624 8498 11652 9318
rect 11518 8463 11574 8472
rect 11612 8492 11664 8498
rect 11426 5400 11482 5409
rect 11426 5335 11482 5344
rect 11532 4758 11560 8463
rect 11612 8434 11664 8440
rect 11612 8016 11664 8022
rect 11612 7958 11664 7964
rect 11624 5778 11652 7958
rect 11716 7750 11744 9687
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11704 7744 11756 7750
rect 11808 7721 11836 7822
rect 11704 7686 11756 7692
rect 11794 7712 11850 7721
rect 11716 7206 11744 7686
rect 11794 7647 11850 7656
rect 11808 7546 11836 7647
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11520 4752 11572 4758
rect 11426 4720 11482 4729
rect 11520 4694 11572 4700
rect 11426 4655 11482 4664
rect 11440 4457 11468 4655
rect 11426 4448 11482 4457
rect 11426 4383 11482 4392
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11440 3913 11468 4014
rect 11426 3904 11482 3913
rect 11426 3839 11482 3848
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11426 2952 11482 2961
rect 11426 2887 11482 2896
rect 11440 2854 11468 2887
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11242 2544 11298 2553
rect 11242 2479 11244 2488
rect 11296 2479 11298 2488
rect 11244 2450 11296 2456
rect 10930 1958 11008 1986
rect 10874 1935 10930 1944
rect 10690 1728 10746 1737
rect 10690 1663 10746 1672
rect 11426 1592 11482 1601
rect 11532 1578 11560 2790
rect 11716 2496 11744 5510
rect 11794 3224 11850 3233
rect 11794 3159 11796 3168
rect 11848 3159 11850 3168
rect 11796 3130 11848 3136
rect 11716 2468 11836 2496
rect 11702 2408 11758 2417
rect 11702 2343 11704 2352
rect 11756 2343 11758 2352
rect 11704 2314 11756 2320
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 1601 11652 2246
rect 11808 1698 11836 2468
rect 11796 1692 11848 1698
rect 11796 1634 11848 1640
rect 11482 1550 11560 1578
rect 11610 1592 11666 1601
rect 11426 1527 11482 1536
rect 11610 1527 11666 1536
rect 10690 1184 10746 1193
rect 10060 1142 10180 1170
rect 10152 480 10180 1142
rect 10690 1119 10746 1128
rect 10704 610 10732 1119
rect 10692 604 10744 610
rect 10692 546 10744 552
rect 10784 604 10836 610
rect 10784 546 10836 552
rect 11336 604 11388 610
rect 11336 546 11388 552
rect 10796 480 10824 546
rect 11348 480 11376 546
rect 11900 480 11928 15438
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12346 14920 12402 14929
rect 12346 14855 12348 14864
rect 12400 14855 12402 14864
rect 12348 14826 12400 14832
rect 12636 14822 12664 14962
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11992 13870 12020 14214
rect 12268 14074 12296 14418
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 12268 13530 12296 14010
rect 12452 13977 12480 14758
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12636 14006 12664 14350
rect 12624 14000 12676 14006
rect 12438 13968 12494 13977
rect 12624 13942 12676 13948
rect 12438 13903 12494 13912
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12268 12986 12296 13466
rect 12544 13326 12572 13874
rect 12636 13394 12664 13942
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12532 13320 12584 13326
rect 12452 13268 12532 13274
rect 12452 13262 12584 13268
rect 12452 13246 12572 13262
rect 12346 13152 12402 13161
rect 12346 13087 12402 13096
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 12176 12209 12204 12310
rect 12162 12200 12218 12209
rect 12162 12135 12218 12144
rect 11978 11656 12034 11665
rect 11978 11591 12034 11600
rect 11992 5778 12020 11591
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12084 10849 12112 11494
rect 12070 10840 12126 10849
rect 12126 10798 12204 10826
rect 12070 10775 12126 10784
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 12084 5114 12112 10610
rect 12176 9897 12204 10798
rect 12162 9888 12218 9897
rect 12162 9823 12218 9832
rect 12164 9648 12216 9654
rect 12162 9616 12164 9625
rect 12216 9616 12218 9625
rect 12162 9551 12218 9560
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12176 7546 12204 8026
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 12162 6624 12218 6633
rect 12162 6559 12218 6568
rect 11992 5086 12112 5114
rect 11992 3670 12020 5086
rect 12176 4078 12204 6559
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 12176 3890 12204 4014
rect 12268 3992 12296 12922
rect 12360 11393 12388 13087
rect 12452 12442 12480 13246
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12346 11384 12402 11393
rect 12346 11319 12402 11328
rect 12360 10130 12480 10146
rect 12348 10124 12480 10130
rect 12400 10118 12480 10124
rect 12348 10066 12400 10072
rect 12452 9654 12480 10118
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12452 9518 12480 9549
rect 12440 9512 12492 9518
rect 12438 9480 12440 9489
rect 12492 9480 12494 9489
rect 12438 9415 12494 9424
rect 12452 9178 12480 9415
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12452 8430 12480 8910
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12544 8242 12572 12582
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12636 11121 12664 11630
rect 12622 11112 12678 11121
rect 12622 11047 12678 11056
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12636 9926 12664 10542
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12622 9616 12678 9625
rect 12622 9551 12678 9560
rect 12636 8537 12664 9551
rect 12622 8528 12678 8537
rect 12622 8463 12678 8472
rect 12728 8378 12756 16623
rect 13280 16590 13308 17167
rect 13372 17134 13400 17478
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13372 16794 13400 17070
rect 13556 16998 13584 17614
rect 13636 17604 13688 17610
rect 13636 17546 13688 17552
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13360 16788 13412 16794
rect 13360 16730 13412 16736
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 12808 15088 12860 15094
rect 12808 15030 12860 15036
rect 12820 13870 12848 15030
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 13004 14414 13032 14962
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 13096 14260 13124 16390
rect 13280 15910 13308 16526
rect 13556 15978 13584 16934
rect 13648 16590 13676 17546
rect 13912 17060 13964 17066
rect 13912 17002 13964 17008
rect 13636 16584 13688 16590
rect 13924 16538 13952 17002
rect 14016 16794 14044 17818
rect 14108 17678 14136 18022
rect 14752 17882 14780 20198
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14922 19272 14978 19281
rect 14922 19207 14978 19216
rect 14936 19174 14964 19207
rect 14924 19168 14976 19174
rect 14924 19110 14976 19116
rect 14936 18834 14964 19110
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14740 17876 14792 17882
rect 14740 17818 14792 17824
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 14108 16726 14136 17614
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14096 16720 14148 16726
rect 14096 16662 14148 16668
rect 13636 16526 13688 16532
rect 13648 16250 13676 16526
rect 13740 16522 13952 16538
rect 13728 16516 13952 16522
rect 13780 16510 13952 16516
rect 13728 16458 13780 16464
rect 13636 16244 13688 16250
rect 13636 16186 13688 16192
rect 13924 16114 13952 16510
rect 14096 16516 14148 16522
rect 14096 16458 14148 16464
rect 14004 16176 14056 16182
rect 14004 16118 14056 16124
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13450 15872 13506 15881
rect 12898 14240 12954 14249
rect 12898 14175 12954 14184
rect 13004 14232 13124 14260
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12820 13530 12848 13806
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12820 12782 12848 13126
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12360 8214 12572 8242
rect 12636 8350 12756 8378
rect 12360 8022 12388 8214
rect 12348 8016 12400 8022
rect 12348 7958 12400 7964
rect 12438 7848 12494 7857
rect 12438 7783 12494 7792
rect 12452 6100 12480 7783
rect 12636 7528 12664 8350
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12728 7818 12756 8230
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12728 7546 12756 7754
rect 12544 7500 12664 7528
rect 12716 7540 12768 7546
rect 12544 6254 12572 7500
rect 12716 7482 12768 7488
rect 12622 7440 12678 7449
rect 12622 7375 12678 7384
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12452 6072 12572 6100
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12452 5166 12480 5850
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12268 3964 12388 3992
rect 12176 3862 12296 3890
rect 12162 3768 12218 3777
rect 12162 3703 12164 3712
rect 12216 3703 12218 3712
rect 12164 3674 12216 3680
rect 12268 3670 12296 3862
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 12256 3664 12308 3670
rect 12256 3606 12308 3612
rect 11992 2825 12020 3606
rect 11978 2816 12034 2825
rect 11978 2751 12034 2760
rect 12360 610 12388 3964
rect 12452 3942 12480 4966
rect 12544 4826 12572 6072
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12440 3120 12492 3126
rect 12438 3088 12440 3097
rect 12492 3088 12494 3097
rect 12438 3023 12494 3032
rect 12348 604 12400 610
rect 12348 546 12400 552
rect 12544 480 12572 4422
rect 12636 3738 12664 7375
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12728 5710 12756 6326
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12728 5234 12756 5646
rect 12820 5370 12848 12718
rect 12912 10282 12940 14175
rect 13004 12374 13032 14232
rect 13082 12608 13138 12617
rect 13082 12543 13138 12552
rect 12992 12368 13044 12374
rect 12992 12310 13044 12316
rect 13004 11354 13032 12310
rect 13096 12209 13124 12543
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13082 12200 13138 12209
rect 13082 12135 13138 12144
rect 13188 11937 13216 12242
rect 13174 11928 13230 11937
rect 13174 11863 13176 11872
rect 13228 11863 13230 11872
rect 13176 11834 13228 11840
rect 13174 11792 13230 11801
rect 13174 11727 13230 11736
rect 13082 11656 13138 11665
rect 13082 11591 13138 11600
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13096 11286 13124 11591
rect 13188 11354 13216 11727
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 13096 10606 13124 11222
rect 13280 10962 13308 15846
rect 13372 15502 13400 15846
rect 13450 15807 13506 15816
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13464 15042 13492 15807
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13634 15464 13690 15473
rect 13556 15162 13584 15438
rect 13832 15450 13860 15642
rect 14016 15570 14044 16118
rect 14108 15706 14136 16458
rect 14384 16114 14412 17138
rect 14752 17066 14780 17818
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14752 16794 14780 17002
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14752 16674 14780 16730
rect 14752 16646 14872 16674
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14752 16250 14780 16526
rect 14740 16244 14792 16250
rect 14740 16186 14792 16192
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 14384 15706 14412 16050
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 13634 15399 13636 15408
rect 13688 15399 13690 15408
rect 13740 15422 13860 15450
rect 13636 15370 13688 15376
rect 13544 15156 13596 15162
rect 13544 15098 13596 15104
rect 13464 15014 13584 15042
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13372 13870 13400 14350
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13372 12458 13400 12718
rect 13363 12430 13400 12458
rect 13363 12356 13391 12430
rect 13363 12328 13400 12356
rect 13188 10934 13308 10962
rect 13188 10713 13216 10934
rect 13266 10840 13322 10849
rect 13266 10775 13322 10784
rect 13174 10704 13230 10713
rect 13174 10639 13230 10648
rect 13084 10600 13136 10606
rect 13084 10542 13136 10548
rect 12912 10254 13216 10282
rect 12898 10160 12954 10169
rect 12898 10095 12900 10104
rect 12952 10095 12954 10104
rect 13084 10124 13136 10130
rect 12900 10066 12952 10072
rect 13084 10066 13136 10072
rect 12898 10024 12954 10033
rect 12898 9959 12954 9968
rect 12912 9654 12940 9959
rect 12992 9920 13044 9926
rect 13096 9897 13124 10066
rect 12992 9862 13044 9868
rect 13082 9888 13138 9897
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 13004 9586 13032 9862
rect 13082 9823 13138 9832
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12900 9512 12952 9518
rect 12898 9480 12900 9489
rect 12952 9480 12954 9489
rect 12898 9415 12954 9424
rect 13004 9042 13032 9522
rect 13082 9072 13138 9081
rect 12992 9036 13044 9042
rect 13082 9007 13138 9016
rect 12992 8978 13044 8984
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12912 8090 12940 8298
rect 13004 8090 13032 8978
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12912 7546 12940 8026
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12912 5574 12940 7278
rect 13096 6610 13124 9007
rect 13188 7154 13216 10254
rect 13280 10062 13308 10775
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13280 9722 13308 9998
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13268 9580 13320 9586
rect 13372 9568 13400 12328
rect 13450 12200 13506 12209
rect 13450 12135 13452 12144
rect 13504 12135 13506 12144
rect 13452 12106 13504 12112
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13320 9540 13400 9568
rect 13268 9522 13320 9528
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 13280 7449 13308 9386
rect 13266 7440 13322 7449
rect 13266 7375 13322 7384
rect 13464 7342 13492 11494
rect 13556 8090 13584 15014
rect 13740 14618 13768 15422
rect 14016 14618 14044 15506
rect 14384 15162 14412 15642
rect 14554 15600 14610 15609
rect 14554 15535 14610 15544
rect 14372 15156 14424 15162
rect 14372 15098 14424 15104
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14108 14550 14136 14826
rect 14096 14544 14148 14550
rect 14096 14486 14148 14492
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 14200 13530 14228 14418
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14384 14113 14412 14214
rect 14370 14104 14426 14113
rect 14370 14039 14426 14048
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14002 13424 14058 13433
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13912 13388 13964 13394
rect 14292 13410 14320 13670
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14002 13359 14058 13368
rect 14200 13382 14320 13410
rect 13912 13330 13964 13336
rect 13648 11694 13676 13330
rect 13924 12986 13952 13330
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13726 12472 13782 12481
rect 13726 12407 13782 12416
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13740 11286 13768 12407
rect 13924 12374 13952 12922
rect 14016 12782 14044 13359
rect 14200 13326 14228 13382
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14200 12442 14228 13262
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 13912 12368 13964 12374
rect 13912 12310 13964 12316
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13924 11694 13952 12174
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13728 11280 13780 11286
rect 13634 11248 13690 11257
rect 13728 11222 13780 11228
rect 13818 11248 13874 11257
rect 13634 11183 13636 11192
rect 13688 11183 13690 11192
rect 13636 11154 13688 11160
rect 13648 10810 13676 11154
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13740 10538 13768 11222
rect 13818 11183 13874 11192
rect 13832 10985 13860 11183
rect 13924 11150 13952 11630
rect 14004 11620 14056 11626
rect 14004 11562 14056 11568
rect 14016 11150 14044 11562
rect 14292 11506 14320 13194
rect 14108 11478 14320 11506
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 13818 10976 13874 10985
rect 13818 10911 13874 10920
rect 13924 10810 13952 11086
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13648 8537 13676 10406
rect 14108 10010 14136 11478
rect 14278 11384 14334 11393
rect 14278 11319 14334 11328
rect 13740 9982 14136 10010
rect 13634 8528 13690 8537
rect 13634 8463 13690 8472
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13544 7200 13596 7206
rect 13188 7126 13308 7154
rect 13544 7142 13596 7148
rect 13174 7032 13230 7041
rect 13174 6967 13176 6976
rect 13228 6967 13230 6976
rect 13176 6938 13228 6944
rect 13174 6896 13230 6905
rect 13174 6831 13230 6840
rect 13188 6662 13216 6831
rect 13004 6582 13124 6610
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 13004 5250 13032 6582
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12820 5222 13032 5250
rect 12820 4978 12848 5222
rect 12728 4950 12848 4978
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 12728 4078 12756 4950
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12636 2922 12664 3674
rect 12728 3641 12756 4014
rect 12714 3632 12770 3641
rect 12714 3567 12770 3576
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 12820 2582 12848 4762
rect 13004 3641 13032 4966
rect 12990 3632 13046 3641
rect 12990 3567 13046 3576
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 12912 2990 12940 3130
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 13096 480 13124 6394
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 13188 5302 13216 5782
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 13188 4486 13216 5238
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13188 4214 13216 4422
rect 13176 4208 13228 4214
rect 13176 4150 13228 4156
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13188 3602 13216 4014
rect 13280 3992 13308 7126
rect 13556 7041 13584 7142
rect 13542 7032 13598 7041
rect 13542 6967 13598 6976
rect 13648 6934 13676 7346
rect 13636 6928 13688 6934
rect 13636 6870 13688 6876
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13372 6497 13400 6734
rect 13358 6488 13414 6497
rect 13358 6423 13360 6432
rect 13412 6423 13414 6432
rect 13360 6394 13412 6400
rect 13634 6352 13690 6361
rect 13634 6287 13690 6296
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13556 5681 13584 6054
rect 13542 5672 13598 5681
rect 13542 5607 13598 5616
rect 13358 5536 13414 5545
rect 13358 5471 13414 5480
rect 13372 4146 13400 5471
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13280 3964 13400 3992
rect 13266 3904 13322 3913
rect 13266 3839 13322 3848
rect 13280 3738 13308 3839
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13372 3602 13400 3964
rect 13556 3913 13584 4422
rect 13542 3904 13598 3913
rect 13542 3839 13598 3848
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13372 3126 13400 3538
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 13648 480 13676 6287
rect 13740 5914 13768 9982
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 13818 8800 13874 8809
rect 13818 8735 13874 8744
rect 13832 7177 13860 8735
rect 13818 7168 13874 7177
rect 13818 7103 13874 7112
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13740 4049 13768 5510
rect 13832 5098 13860 6598
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13924 4758 13952 9862
rect 14016 5234 14044 9862
rect 14292 9654 14320 11319
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14292 9450 14320 9590
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 14384 9353 14412 13466
rect 14464 13388 14516 13394
rect 14464 13330 14516 13336
rect 14476 12442 14504 13330
rect 14568 13258 14596 15535
rect 14844 14618 14872 16646
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15396 16046 15424 16934
rect 15474 16416 15530 16425
rect 15474 16351 15530 16360
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15396 15706 15424 15982
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15396 15502 15424 15642
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 15212 14414 15240 14758
rect 15304 14618 15332 15302
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15396 14414 15424 15438
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15200 13864 15252 13870
rect 15488 13852 15516 16351
rect 15568 15972 15620 15978
rect 15568 15914 15620 15920
rect 15580 13954 15608 15914
rect 15672 14550 15700 17614
rect 17040 16788 17092 16794
rect 17040 16730 17092 16736
rect 17052 16697 17080 16730
rect 17038 16688 17094 16697
rect 17038 16623 17094 16632
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15856 15502 15884 16526
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16776 16250 16804 16390
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 17144 15910 17172 16594
rect 17236 16454 17264 26794
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 23216 19281 23244 27520
rect 23478 27503 23534 27512
rect 23492 26858 23520 27503
rect 23570 26888 23626 26897
rect 23480 26852 23532 26858
rect 23570 26823 23626 26832
rect 23480 26794 23532 26800
rect 23478 20088 23534 20097
rect 23478 20023 23534 20032
rect 23202 19272 23258 19281
rect 23202 19207 23258 19216
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 23492 17218 23520 20023
rect 23400 17190 23520 17218
rect 18050 16960 18106 16969
rect 18050 16895 18106 16904
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 16580 15904 16632 15910
rect 17132 15904 17184 15910
rect 16580 15846 16632 15852
rect 17130 15872 17132 15881
rect 17184 15872 17186 15881
rect 16028 15632 16080 15638
rect 16028 15574 16080 15580
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 16040 15337 16068 15574
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16026 15328 16082 15337
rect 16026 15263 16082 15272
rect 16040 15162 16068 15263
rect 16408 15201 16436 15506
rect 16592 15434 16620 15846
rect 17130 15807 17186 15816
rect 17592 15564 17644 15570
rect 17592 15506 17644 15512
rect 17316 15496 17368 15502
rect 17314 15464 17316 15473
rect 17368 15464 17370 15473
rect 16580 15428 16632 15434
rect 17314 15399 17370 15408
rect 16580 15370 16632 15376
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16394 15192 16450 15201
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 16120 15156 16172 15162
rect 16394 15127 16396 15136
rect 16120 15098 16172 15104
rect 16448 15127 16450 15136
rect 16396 15098 16448 15104
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15660 14544 15712 14550
rect 15660 14486 15712 14492
rect 15672 14074 15700 14486
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15764 14074 15792 14350
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15580 13926 15792 13954
rect 15488 13824 15700 13852
rect 15200 13806 15252 13812
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14660 12986 14688 13738
rect 15212 13546 15240 13806
rect 15120 13530 15240 13546
rect 15108 13524 15240 13530
rect 15160 13518 15240 13524
rect 15108 13466 15160 13472
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 15580 12850 15608 13126
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15672 12730 15700 13824
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 15580 12702 15700 12730
rect 15304 12442 15332 12650
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15382 12336 15438 12345
rect 15382 12271 15438 12280
rect 15396 12073 15424 12271
rect 15382 12064 15438 12073
rect 14956 11996 15252 12016
rect 15382 11999 15438 12008
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15108 11824 15160 11830
rect 15108 11766 15160 11772
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14660 11354 14688 11698
rect 15120 11354 15148 11766
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10606 15332 11086
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 14556 10532 14608 10538
rect 14556 10474 14608 10480
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14476 10266 14504 10406
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14476 9518 14504 10202
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14464 9376 14516 9382
rect 14370 9344 14426 9353
rect 14464 9318 14516 9324
rect 14370 9279 14426 9288
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14108 8430 14136 8774
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14200 7857 14228 8570
rect 14278 8256 14334 8265
rect 14278 8191 14334 8200
rect 14186 7848 14242 7857
rect 14186 7783 14242 7792
rect 14096 6724 14148 6730
rect 14096 6666 14148 6672
rect 14108 6186 14136 6666
rect 14096 6180 14148 6186
rect 14096 6122 14148 6128
rect 14108 5914 14136 6122
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 14016 4826 14044 5170
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 13912 4752 13964 4758
rect 13912 4694 13964 4700
rect 13924 4282 13952 4694
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 14016 4282 14044 4626
rect 14108 4622 14136 5850
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 13726 4040 13782 4049
rect 13726 3975 13782 3984
rect 14108 3738 14136 4558
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 13728 3528 13780 3534
rect 13820 3528 13872 3534
rect 13728 3470 13780 3476
rect 13818 3496 13820 3505
rect 13872 3496 13874 3505
rect 13740 3369 13768 3470
rect 13818 3431 13874 3440
rect 13726 3360 13782 3369
rect 13726 3295 13782 3304
rect 13740 2854 13768 3295
rect 13832 3194 13860 3431
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 14002 2816 14058 2825
rect 14200 2802 14228 5714
rect 14292 5250 14320 8191
rect 14476 8090 14504 9318
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14370 7848 14426 7857
rect 14370 7783 14426 7792
rect 14384 7585 14412 7783
rect 14370 7576 14426 7585
rect 14370 7511 14426 7520
rect 14372 7268 14424 7274
rect 14372 7210 14424 7216
rect 14384 6458 14412 7210
rect 14476 7002 14504 8026
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14568 6882 14596 10474
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 14832 9988 14884 9994
rect 14832 9930 14884 9936
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14646 8528 14702 8537
rect 14646 8463 14702 8472
rect 14476 6854 14596 6882
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14384 5370 14412 6394
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14292 5222 14412 5250
rect 14002 2751 14058 2760
rect 14108 2774 14228 2802
rect 14016 2650 14044 2751
rect 14108 2666 14136 2774
rect 14004 2644 14056 2650
rect 14108 2638 14320 2666
rect 14004 2586 14056 2592
rect 14292 480 14320 2638
rect 14384 2145 14412 5222
rect 14476 3754 14504 6854
rect 14554 6080 14610 6089
rect 14554 6015 14610 6024
rect 14568 4146 14596 6015
rect 14660 4826 14688 8463
rect 14752 8430 14780 8978
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14738 8120 14794 8129
rect 14844 8090 14872 9930
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 15028 9178 15056 9522
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 15304 8922 15332 10134
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15396 9178 15424 9998
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15120 8906 15332 8922
rect 15108 8900 15332 8906
rect 15160 8894 15332 8900
rect 15108 8842 15160 8848
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 14738 8055 14794 8064
rect 14832 8084 14884 8090
rect 14752 5914 14780 8055
rect 14832 8026 14884 8032
rect 15028 8022 15056 8366
rect 15120 8090 15148 8366
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15016 8016 15068 8022
rect 15016 7958 15068 7964
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15304 7478 15332 8894
rect 15396 8362 15424 9114
rect 15384 8356 15436 8362
rect 15384 8298 15436 8304
rect 15292 7472 15344 7478
rect 15292 7414 15344 7420
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 15382 5808 15438 5817
rect 15382 5743 15438 5752
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 14752 4146 14780 4422
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15304 4185 15332 4422
rect 15290 4176 15346 4185
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14740 4140 14792 4146
rect 15290 4111 15346 4120
rect 14740 4082 14792 4088
rect 14476 3726 14688 3754
rect 14752 3738 14780 4082
rect 15290 4040 15346 4049
rect 15016 4004 15068 4010
rect 15290 3975 15346 3984
rect 15016 3946 15068 3952
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 14476 2514 14504 2790
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 14370 2136 14426 2145
rect 14370 2071 14426 2080
rect 14568 1329 14596 3334
rect 14660 1442 14688 3726
rect 14740 3732 14792 3738
rect 14792 3692 14872 3720
rect 14740 3674 14792 3680
rect 14844 2922 14872 3692
rect 15028 3466 15056 3946
rect 15304 3602 15332 3975
rect 15396 3738 15424 5743
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15488 3618 15516 12582
rect 15580 12102 15608 12702
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15580 11694 15608 12038
rect 15672 11898 15700 12582
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15580 11529 15608 11630
rect 15566 11520 15622 11529
rect 15566 11455 15622 11464
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 15580 10266 15608 10542
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15568 8424 15620 8430
rect 15568 8366 15620 8372
rect 15580 7954 15608 8366
rect 15672 8294 15700 9046
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15580 7002 15608 7754
rect 15672 7750 15700 8230
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15672 7546 15700 7686
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15660 4548 15712 4554
rect 15660 4490 15712 4496
rect 15568 4004 15620 4010
rect 15568 3946 15620 3952
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15396 3590 15516 3618
rect 15016 3460 15068 3466
rect 15016 3402 15068 3408
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 15016 2916 15068 2922
rect 15016 2858 15068 2864
rect 15028 2689 15056 2858
rect 15396 2802 15424 3590
rect 15580 2825 15608 3946
rect 15672 3942 15700 4490
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15672 3777 15700 3878
rect 15658 3768 15714 3777
rect 15658 3703 15714 3712
rect 15764 2836 15792 13926
rect 15856 13530 15884 14554
rect 16040 13841 16068 15098
rect 16026 13832 16082 13841
rect 15936 13796 15988 13802
rect 16026 13767 16082 13776
rect 15936 13738 15988 13744
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 15948 13410 15976 13738
rect 15856 13382 15976 13410
rect 15856 12442 15884 13382
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15934 13016 15990 13025
rect 16040 12986 16068 13262
rect 15934 12951 15936 12960
rect 15988 12951 15990 12960
rect 16028 12980 16080 12986
rect 15936 12922 15988 12928
rect 16028 12922 16080 12928
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15948 12345 15976 12786
rect 15934 12336 15990 12345
rect 15934 12271 15990 12280
rect 15948 11830 15976 12271
rect 16040 12238 16068 12922
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 15936 11824 15988 11830
rect 15936 11766 15988 11772
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15948 10305 15976 11494
rect 15934 10296 15990 10305
rect 15934 10231 15990 10240
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 15948 9518 15976 10066
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15844 9376 15896 9382
rect 15842 9344 15844 9353
rect 15896 9344 15898 9353
rect 15842 9279 15898 9288
rect 15948 7993 15976 9454
rect 16132 9450 16160 15098
rect 16500 14958 16528 15302
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 15934 7984 15990 7993
rect 15844 7948 15896 7954
rect 15934 7919 15990 7928
rect 15844 7890 15896 7896
rect 15856 7857 15884 7890
rect 15842 7848 15898 7857
rect 15842 7783 15898 7792
rect 15856 7546 15884 7783
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15856 6254 15884 6734
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 15856 5778 15884 6190
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 15844 5092 15896 5098
rect 15844 5034 15896 5040
rect 15856 3534 15884 5034
rect 15948 4049 15976 5510
rect 16040 4826 16068 9318
rect 16316 8673 16344 14894
rect 16592 14890 16620 15370
rect 17328 15162 17356 15399
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 16580 14884 16632 14890
rect 16580 14826 16632 14832
rect 17604 14822 17632 15506
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 16580 14544 16632 14550
rect 16580 14486 16632 14492
rect 16592 14278 16620 14486
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16408 13938 16436 14214
rect 16488 14000 16540 14006
rect 16488 13942 16540 13948
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16500 12866 16528 13942
rect 16592 13394 16620 14214
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16684 13530 16712 13874
rect 16776 13802 16804 14214
rect 16868 13977 16896 14758
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 16854 13968 16910 13977
rect 16854 13903 16910 13912
rect 17236 13870 17264 14418
rect 17328 14074 17356 14554
rect 17604 14346 17632 14758
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 16764 13796 16816 13802
rect 16764 13738 16816 13744
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16592 12986 16620 13330
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16500 12838 16620 12866
rect 16592 12782 16620 12838
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16592 11558 16620 12174
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 16394 10704 16450 10713
rect 16394 10639 16450 10648
rect 16408 10010 16436 10639
rect 16488 10600 16540 10606
rect 16592 10588 16620 11222
rect 16540 10560 16620 10588
rect 16488 10542 16540 10548
rect 16684 10146 16712 12650
rect 16854 12064 16910 12073
rect 16854 11999 16910 12008
rect 16868 10810 16896 11999
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 16592 10118 16712 10146
rect 16408 9982 16528 10010
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16408 9382 16436 9862
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16302 8664 16358 8673
rect 16302 8599 16358 8608
rect 16304 8560 16356 8566
rect 16304 8502 16356 8508
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16132 4865 16160 7142
rect 16118 4856 16174 4865
rect 16028 4820 16080 4826
rect 16118 4791 16174 4800
rect 16224 4808 16252 7482
rect 16316 6866 16344 8502
rect 16408 8265 16436 9318
rect 16394 8256 16450 8265
rect 16394 8191 16450 8200
rect 16394 7168 16450 7177
rect 16394 7103 16450 7112
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16316 5914 16344 6802
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16224 4780 16344 4808
rect 16028 4762 16080 4768
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 16224 4282 16252 4626
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 15934 4040 15990 4049
rect 15934 3975 15990 3984
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15948 3738 15976 3878
rect 16224 3738 16252 4218
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 16212 3596 16264 3602
rect 16212 3538 16264 3544
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15856 3194 15884 3470
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 16224 3126 16252 3538
rect 16316 3369 16344 4780
rect 16408 4010 16436 7103
rect 16500 6633 16528 9982
rect 16486 6624 16542 6633
rect 16486 6559 16542 6568
rect 16500 6322 16528 6559
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16500 5914 16528 6258
rect 16592 6225 16620 10118
rect 16672 10056 16724 10062
rect 16670 10024 16672 10033
rect 16724 10024 16726 10033
rect 16670 9959 16726 9968
rect 17144 9654 17172 12786
rect 17328 12306 17356 13466
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17328 11898 17356 12242
rect 17224 11892 17276 11898
rect 17224 11834 17276 11840
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17236 11354 17264 11834
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17512 11150 17540 11494
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17406 10568 17462 10577
rect 17406 10503 17462 10512
rect 17314 10296 17370 10305
rect 17314 10231 17370 10240
rect 17132 9648 17184 9654
rect 17132 9590 17184 9596
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16684 8634 16712 9522
rect 16946 8664 17002 8673
rect 16672 8628 16724 8634
rect 16946 8599 17002 8608
rect 16672 8570 16724 8576
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16776 7886 16804 8298
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16776 7002 16804 7822
rect 16960 7750 16988 8599
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16868 7410 16896 7686
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16960 7290 16988 7686
rect 17328 7478 17356 10231
rect 17420 8090 17448 10503
rect 17512 10470 17540 11086
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17512 9654 17540 10406
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17500 9648 17552 9654
rect 17500 9590 17552 9596
rect 17604 9178 17632 9862
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17512 8634 17540 8842
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17420 7546 17448 8026
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17316 7472 17368 7478
rect 17316 7414 17368 7420
rect 16868 7262 16988 7290
rect 16868 7206 16896 7262
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 16868 6361 16896 7142
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17420 6458 17448 6598
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 16854 6352 16910 6361
rect 16854 6287 16910 6296
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16578 6216 16634 6225
rect 16578 6151 16634 6160
rect 16854 6216 16910 6225
rect 16854 6151 16910 6160
rect 16868 6118 16896 6151
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16488 5024 16540 5030
rect 16486 4992 16488 5001
rect 16540 4992 16542 5001
rect 16486 4927 16542 4936
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16500 4060 16528 4762
rect 16592 4758 16620 6054
rect 17052 5846 17080 6258
rect 17040 5840 17092 5846
rect 17040 5782 17092 5788
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16868 5370 16896 5714
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 17052 4826 17080 5782
rect 17500 5092 17552 5098
rect 17500 5034 17552 5040
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 16580 4752 16632 4758
rect 16580 4694 16632 4700
rect 17408 4752 17460 4758
rect 17408 4694 17460 4700
rect 16580 4072 16632 4078
rect 16500 4032 16580 4060
rect 16580 4014 16632 4020
rect 17130 4040 17186 4049
rect 16396 4004 16448 4010
rect 17130 3975 17186 3984
rect 17314 4040 17370 4049
rect 17314 3975 17370 3984
rect 16396 3946 16448 3952
rect 16408 3602 16436 3946
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 16302 3360 16358 3369
rect 16302 3295 16358 3304
rect 16212 3120 16264 3126
rect 16212 3062 16264 3068
rect 15365 2774 15424 2802
rect 15566 2816 15622 2825
rect 14738 2680 14794 2689
rect 14738 2615 14794 2624
rect 15014 2680 15070 2689
rect 15365 2666 15393 2774
rect 15566 2751 15622 2760
rect 15755 2808 15792 2836
rect 15755 2666 15783 2808
rect 16854 2680 16910 2689
rect 15365 2638 15424 2666
rect 15755 2638 16068 2666
rect 15014 2615 15070 2624
rect 14752 2009 14780 2615
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14738 2000 14794 2009
rect 14738 1935 14794 1944
rect 14660 1414 14872 1442
rect 14554 1320 14610 1329
rect 14554 1255 14610 1264
rect 14844 480 14872 1414
rect 15396 480 15424 2638
rect 16040 480 16068 2638
rect 16854 2615 16856 2624
rect 16908 2615 16910 2624
rect 16856 2586 16908 2592
rect 16578 1592 16634 1601
rect 16578 1527 16634 1536
rect 16592 480 16620 1527
rect 17144 480 17172 3975
rect 17224 3732 17276 3738
rect 17328 3720 17356 3975
rect 17420 3738 17448 4694
rect 17512 4622 17540 5034
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 17512 4282 17540 4558
rect 17696 4554 17724 15982
rect 17774 15056 17830 15065
rect 17774 14991 17830 15000
rect 17788 14618 17816 14991
rect 17960 14884 18012 14890
rect 17880 14844 17960 14872
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17788 12986 17816 14418
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17774 11248 17830 11257
rect 17774 11183 17830 11192
rect 17788 10130 17816 11183
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17788 9654 17816 10066
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17788 8430 17816 9454
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17788 8022 17816 8366
rect 17880 8090 17908 14844
rect 17960 14826 18012 14832
rect 18064 14074 18092 16895
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 20074 16552 20130 16561
rect 20074 16487 20130 16496
rect 18236 16176 18288 16182
rect 18234 16144 18236 16153
rect 18288 16144 18290 16153
rect 18234 16079 18290 16088
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19444 15609 19472 15642
rect 19430 15600 19486 15609
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 19340 15564 19392 15570
rect 19430 15535 19486 15544
rect 19340 15506 19392 15512
rect 18236 15360 18288 15366
rect 18236 15302 18288 15308
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 17960 12912 18012 12918
rect 17960 12854 18012 12860
rect 17972 12442 18000 12854
rect 18144 12708 18196 12714
rect 18144 12650 18196 12656
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17972 11762 18000 12038
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 18064 11665 18092 12582
rect 18050 11656 18106 11665
rect 18050 11591 18106 11600
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17972 10538 18000 10950
rect 17960 10532 18012 10538
rect 17960 10474 18012 10480
rect 17972 10266 18000 10474
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18064 10198 18092 11494
rect 18156 11354 18184 12650
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18052 10192 18104 10198
rect 18052 10134 18104 10140
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17972 8838 18000 9386
rect 18052 9036 18104 9042
rect 18052 8978 18104 8984
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17972 8634 18000 8774
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17972 7954 18000 8570
rect 18064 8566 18092 8978
rect 18052 8560 18104 8566
rect 18052 8502 18104 8508
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 18064 7546 18092 8026
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 18156 7342 18184 9998
rect 18248 9194 18276 15302
rect 18432 14890 18460 15506
rect 19352 14958 19380 15506
rect 20088 15473 20116 16487
rect 23400 16266 23428 17190
rect 23478 17096 23534 17105
rect 23478 17031 23534 17040
rect 23308 16238 23428 16266
rect 22284 15496 22336 15502
rect 20074 15464 20130 15473
rect 22284 15438 22336 15444
rect 20074 15399 20130 15408
rect 18880 14952 18932 14958
rect 19340 14952 19392 14958
rect 18880 14894 18932 14900
rect 19168 14900 19340 14906
rect 19168 14894 19392 14900
rect 18420 14884 18472 14890
rect 18420 14826 18472 14832
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18616 14521 18644 14554
rect 18602 14512 18658 14521
rect 18602 14447 18658 14456
rect 18602 14376 18658 14385
rect 18602 14311 18658 14320
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18432 13734 18460 14214
rect 18616 13938 18644 14311
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18602 13832 18658 13841
rect 18602 13767 18658 13776
rect 18420 13728 18472 13734
rect 18418 13696 18420 13705
rect 18472 13696 18474 13705
rect 18418 13631 18474 13640
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18340 12646 18368 13126
rect 18524 12889 18552 13126
rect 18510 12880 18566 12889
rect 18510 12815 18566 12824
rect 18616 12730 18644 13767
rect 18524 12702 18644 12730
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18248 9166 18368 9194
rect 18236 9036 18288 9042
rect 18236 8978 18288 8984
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18156 7002 18184 7278
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18052 6928 18104 6934
rect 18052 6870 18104 6876
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17788 5370 17816 6122
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 17684 4548 17736 4554
rect 17684 4490 17736 4496
rect 17500 4276 17552 4282
rect 17500 4218 17552 4224
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17276 3692 17356 3720
rect 17408 3732 17460 3738
rect 17224 3674 17276 3680
rect 17408 3674 17460 3680
rect 17500 3664 17552 3670
rect 17500 3606 17552 3612
rect 17512 3194 17540 3606
rect 17500 3188 17552 3194
rect 17500 3130 17552 3136
rect 17696 2553 17724 4082
rect 17788 3194 17816 5306
rect 18064 3738 18092 6870
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18156 5166 18184 5510
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18248 4146 18276 8978
rect 18340 6254 18368 9166
rect 18524 7818 18552 12702
rect 18602 12608 18658 12617
rect 18602 12543 18658 12552
rect 18616 8838 18644 12543
rect 18708 10554 18736 14758
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18800 13025 18828 13330
rect 18786 13016 18842 13025
rect 18786 12951 18842 12960
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18800 11354 18828 11494
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18800 10674 18828 11290
rect 18892 10810 18920 14894
rect 19168 14878 19380 14894
rect 18972 13320 19024 13326
rect 18970 13288 18972 13297
rect 19064 13320 19116 13326
rect 19024 13288 19026 13297
rect 19064 13262 19116 13268
rect 18970 13223 19026 13232
rect 18984 12594 19012 13223
rect 19076 12714 19104 13262
rect 19064 12708 19116 12714
rect 19064 12650 19116 12656
rect 18984 12566 19104 12594
rect 19076 12442 19104 12566
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 18970 12336 19026 12345
rect 18970 12271 19026 12280
rect 18984 12102 19012 12271
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18972 11824 19024 11830
rect 18972 11766 19024 11772
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18708 10526 18828 10554
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18708 9178 18736 10406
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18694 7440 18750 7449
rect 18694 7375 18750 7384
rect 18708 6798 18736 7375
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18340 5778 18368 6190
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18340 4146 18368 4422
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 18236 3936 18288 3942
rect 18234 3904 18236 3913
rect 18288 3904 18290 3913
rect 18234 3839 18290 3848
rect 18248 3738 18276 3839
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18142 3496 18198 3505
rect 18142 3431 18144 3440
rect 18196 3431 18198 3440
rect 18144 3402 18196 3408
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 17774 2952 17830 2961
rect 18064 2922 18092 2994
rect 18156 2990 18184 3402
rect 18432 3097 18460 6054
rect 18524 4826 18552 6598
rect 18708 6390 18736 6734
rect 18696 6384 18748 6390
rect 18696 6326 18748 6332
rect 18800 5250 18828 10526
rect 18984 7721 19012 11766
rect 19064 11212 19116 11218
rect 19064 11154 19116 11160
rect 19076 10470 19104 11154
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 19076 8090 19104 8774
rect 19064 8084 19116 8090
rect 19064 8026 19116 8032
rect 18970 7712 19026 7721
rect 18970 7647 19026 7656
rect 18970 7440 19026 7449
rect 18970 7375 19026 7384
rect 18984 7274 19012 7375
rect 18972 7268 19024 7274
rect 18972 7210 19024 7216
rect 18970 7032 19026 7041
rect 18970 6967 19026 6976
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 18892 6769 18920 6802
rect 18878 6760 18934 6769
rect 18878 6695 18934 6704
rect 18892 5914 18920 6695
rect 18984 5914 19012 6967
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 19076 6458 19104 6734
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18972 5908 19024 5914
rect 18972 5850 19024 5856
rect 18616 5222 18828 5250
rect 19064 5296 19116 5302
rect 19064 5238 19116 5244
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 18616 3670 18644 5222
rect 18786 5128 18842 5137
rect 18786 5063 18842 5072
rect 18800 4321 18828 5063
rect 19076 4758 19104 5238
rect 19168 4826 19196 14878
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19248 14272 19300 14278
rect 19300 14232 19380 14260
rect 19248 14214 19300 14220
rect 19248 13864 19300 13870
rect 19352 13852 19380 14232
rect 19444 14074 19472 14418
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19300 13824 19380 13852
rect 19248 13806 19300 13812
rect 19352 12986 19380 13824
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19430 13560 19486 13569
rect 19622 13552 19918 13572
rect 19430 13495 19486 13504
rect 19444 13462 19472 13495
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19800 13456 19852 13462
rect 19800 13398 19852 13404
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19260 11830 19288 12582
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19248 11824 19300 11830
rect 19352 11801 19380 12242
rect 19248 11766 19300 11772
rect 19338 11792 19394 11801
rect 19338 11727 19394 11736
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 19338 11656 19394 11665
rect 19260 11558 19288 11630
rect 19338 11591 19394 11600
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19260 11286 19288 11494
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19352 10554 19380 11591
rect 19260 10526 19380 10554
rect 19444 10554 19472 13262
rect 19616 13184 19668 13190
rect 19614 13152 19616 13161
rect 19812 13161 19840 13398
rect 19668 13152 19670 13161
rect 19614 13087 19670 13096
rect 19798 13152 19854 13161
rect 19798 13087 19854 13096
rect 19628 12782 19656 13087
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19524 12232 19576 12238
rect 19522 12200 19524 12209
rect 19616 12232 19668 12238
rect 19576 12200 19578 12209
rect 19616 12174 19668 12180
rect 19522 12135 19578 12144
rect 19628 12102 19656 12174
rect 19616 12096 19668 12102
rect 19616 12038 19668 12044
rect 19996 11642 20024 14214
rect 20088 13326 20116 15399
rect 20444 15088 20496 15094
rect 20444 15030 20496 15036
rect 20352 14952 20404 14958
rect 20352 14894 20404 14900
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 20180 13870 20208 14418
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 20088 12850 20116 13126
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 20088 12073 20116 12786
rect 20074 12064 20130 12073
rect 20074 11999 20130 12008
rect 20180 11801 20208 13806
rect 20166 11792 20222 11801
rect 20166 11727 20222 11736
rect 19996 11614 20208 11642
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 19444 10526 19564 10554
rect 19260 10010 19288 10526
rect 19432 10464 19484 10470
rect 19338 10432 19394 10441
rect 19432 10406 19484 10412
rect 19338 10367 19394 10376
rect 19352 10130 19380 10367
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19260 9982 19380 10010
rect 19444 9994 19472 10406
rect 19246 8528 19302 8537
rect 19246 8463 19302 8472
rect 19260 8362 19288 8463
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19260 8090 19288 8298
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19260 7410 19288 8026
rect 19352 7426 19380 9982
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 19444 9722 19472 9930
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19444 8401 19472 8774
rect 19430 8392 19486 8401
rect 19430 8327 19486 8336
rect 19248 7404 19300 7410
rect 19352 7398 19472 7426
rect 19248 7346 19300 7352
rect 19444 6934 19472 7398
rect 19432 6928 19484 6934
rect 19432 6870 19484 6876
rect 19536 5914 19564 10526
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19892 10124 19944 10130
rect 19892 10066 19944 10072
rect 19904 9722 19932 10066
rect 19982 10024 20038 10033
rect 19982 9959 19984 9968
rect 20036 9959 20038 9968
rect 19984 9930 20036 9936
rect 19892 9716 19944 9722
rect 19892 9658 19944 9664
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19812 7546 19840 7822
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19996 7478 20024 7890
rect 19984 7472 20036 7478
rect 19984 7414 20036 7420
rect 19890 7304 19946 7313
rect 19890 7239 19892 7248
rect 19944 7239 19946 7248
rect 19892 7210 19944 7216
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19996 7002 20024 7414
rect 19984 6996 20036 7002
rect 19984 6938 20036 6944
rect 19616 6656 19668 6662
rect 19616 6598 19668 6604
rect 19628 6186 19656 6598
rect 19616 6180 19668 6186
rect 19616 6122 19668 6128
rect 19984 6180 20036 6186
rect 19984 6122 20036 6128
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19430 5672 19486 5681
rect 19430 5607 19486 5616
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19352 4826 19380 5510
rect 19156 4820 19208 4826
rect 19156 4762 19208 4768
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19064 4752 19116 4758
rect 19444 4706 19472 5607
rect 19536 5370 19564 5850
rect 19892 5704 19944 5710
rect 19996 5692 20024 6122
rect 19944 5664 20024 5692
rect 19892 5646 19944 5652
rect 19524 5364 19576 5370
rect 19524 5306 19576 5312
rect 19904 5234 19932 5646
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19064 4694 19116 4700
rect 19352 4678 19472 4706
rect 19524 4684 19576 4690
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18786 4312 18842 4321
rect 18786 4247 18842 4256
rect 18892 4146 18920 4422
rect 18696 4140 18748 4146
rect 18880 4140 18932 4146
rect 18748 4100 18828 4128
rect 18696 4082 18748 4088
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18418 3088 18474 3097
rect 18418 3023 18474 3032
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 17774 2887 17830 2896
rect 18052 2916 18104 2922
rect 17682 2544 17738 2553
rect 17682 2479 17738 2488
rect 17314 2000 17370 2009
rect 17314 1935 17370 1944
rect 17328 1465 17356 1935
rect 17314 1456 17370 1465
rect 17314 1391 17370 1400
rect 17788 480 17816 2887
rect 18052 2858 18104 2864
rect 18064 2650 18092 2858
rect 18524 2650 18552 3470
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18156 2446 18184 2586
rect 18708 2582 18736 3674
rect 18696 2576 18748 2582
rect 18696 2518 18748 2524
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18326 1728 18382 1737
rect 18326 1663 18382 1672
rect 18340 480 18368 1663
rect 5538 0 5594 480
rect 6090 0 6146 480
rect 6642 0 6698 480
rect 7286 0 7342 480
rect 7838 0 7894 480
rect 8390 0 8446 480
rect 9034 0 9090 480
rect 9586 0 9642 480
rect 10138 0 10194 480
rect 10782 0 10838 480
rect 11334 0 11390 480
rect 11886 0 11942 480
rect 12530 0 12586 480
rect 13082 0 13138 480
rect 13634 0 13690 480
rect 14278 0 14334 480
rect 14830 0 14886 480
rect 15382 0 15438 480
rect 16026 0 16082 480
rect 16578 0 16634 480
rect 17130 0 17186 480
rect 17774 0 17830 480
rect 18326 0 18382 480
rect 18800 377 18828 4100
rect 18880 4082 18932 4088
rect 18892 3738 18920 4082
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 19352 3074 19380 4678
rect 19524 4626 19576 4632
rect 19536 3738 19564 4626
rect 19708 4616 19760 4622
rect 19708 4558 19760 4564
rect 19720 4282 19748 4558
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19444 3194 19472 3674
rect 20088 3602 20116 10950
rect 20180 5137 20208 11614
rect 20272 9178 20300 14214
rect 20364 13841 20392 14894
rect 20350 13832 20406 13841
rect 20350 13767 20406 13776
rect 20350 13696 20406 13705
rect 20350 13631 20406 13640
rect 20364 13258 20392 13631
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 20352 12708 20404 12714
rect 20352 12650 20404 12656
rect 20364 12345 20392 12650
rect 20350 12336 20406 12345
rect 20350 12271 20406 12280
rect 20364 11257 20392 12271
rect 20350 11248 20406 11257
rect 20350 11183 20406 11192
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20364 9994 20392 10406
rect 20456 10266 20484 15030
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20352 9988 20404 9994
rect 20352 9930 20404 9936
rect 20364 9722 20392 9930
rect 20352 9716 20404 9722
rect 20352 9658 20404 9664
rect 20456 9518 20484 10202
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20272 7342 20300 9114
rect 20364 8634 20392 9114
rect 20548 9042 20576 14758
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20640 13734 20668 14418
rect 20810 14104 20866 14113
rect 20810 14039 20866 14048
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 20640 10810 20668 13670
rect 20718 13288 20774 13297
rect 20718 13223 20774 13232
rect 20732 12986 20760 13223
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20732 10606 20760 11018
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 20732 10266 20760 10542
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 20628 9104 20680 9110
rect 20628 9046 20680 9052
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20444 8832 20496 8838
rect 20444 8774 20496 8780
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 20364 7886 20392 8230
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 20166 5128 20222 5137
rect 20166 5063 20222 5072
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 20272 4593 20300 4966
rect 20258 4584 20314 4593
rect 20258 4519 20314 4528
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 19352 3046 19472 3074
rect 19444 2666 19472 3046
rect 19904 2961 19932 3334
rect 19890 2952 19946 2961
rect 19890 2887 19946 2896
rect 20364 2825 20392 7142
rect 20456 5370 20484 8774
rect 20548 8022 20576 8978
rect 20640 8945 20668 9046
rect 20626 8936 20682 8945
rect 20626 8871 20682 8880
rect 20640 8634 20668 8871
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20628 8424 20680 8430
rect 20626 8392 20628 8401
rect 20680 8392 20682 8401
rect 20626 8327 20682 8336
rect 20628 8084 20680 8090
rect 20732 8072 20760 8774
rect 20680 8044 20760 8072
rect 20628 8026 20680 8032
rect 20536 8016 20588 8022
rect 20536 7958 20588 7964
rect 20640 7002 20668 8026
rect 20718 7712 20774 7721
rect 20718 7647 20774 7656
rect 20732 7206 20760 7647
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20640 6118 20668 6802
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20640 5574 20668 6054
rect 20628 5568 20680 5574
rect 20628 5510 20680 5516
rect 20444 5364 20496 5370
rect 20444 5306 20496 5312
rect 20442 5264 20498 5273
rect 20442 5199 20498 5208
rect 20456 5098 20484 5199
rect 20444 5092 20496 5098
rect 20444 5034 20496 5040
rect 20456 4826 20484 5034
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 20548 4758 20576 4966
rect 20536 4752 20588 4758
rect 20536 4694 20588 4700
rect 20640 4622 20668 5510
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 20732 4321 20760 7142
rect 20824 4826 20852 14039
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 20902 13016 20958 13025
rect 20902 12951 20904 12960
rect 20956 12951 20958 12960
rect 20904 12922 20956 12928
rect 21100 12186 21128 13262
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 20916 12158 21128 12186
rect 20916 9058 20944 12158
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 21008 11762 21036 12038
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 21008 11558 21036 11698
rect 21088 11620 21140 11626
rect 21088 11562 21140 11568
rect 20996 11552 21048 11558
rect 21100 11529 21128 11562
rect 20996 11494 21048 11500
rect 21086 11520 21142 11529
rect 21008 11218 21036 11494
rect 21086 11455 21142 11464
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 21008 9994 21036 11154
rect 21100 10674 21128 11290
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20996 9988 21048 9994
rect 20996 9930 21048 9936
rect 21192 9178 21220 12582
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21284 10266 21312 12174
rect 21456 11824 21508 11830
rect 21456 11766 21508 11772
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21376 10674 21404 11630
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21364 10260 21416 10266
rect 21364 10202 21416 10208
rect 21284 9722 21312 10202
rect 21272 9716 21324 9722
rect 21272 9658 21324 9664
rect 21376 9586 21404 10202
rect 21364 9580 21416 9586
rect 21364 9522 21416 9528
rect 21362 9208 21418 9217
rect 21180 9172 21232 9178
rect 21362 9143 21364 9152
rect 21180 9114 21232 9120
rect 21416 9143 21418 9152
rect 21364 9114 21416 9120
rect 20916 9030 21036 9058
rect 20904 8968 20956 8974
rect 20904 8910 20956 8916
rect 20916 8362 20944 8910
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 20902 8256 20958 8265
rect 20902 8191 20958 8200
rect 20916 7886 20944 8191
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 20916 6798 20944 7822
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 21008 4842 21036 9030
rect 21272 8900 21324 8906
rect 21272 8842 21324 8848
rect 21284 8022 21312 8842
rect 21364 8832 21416 8838
rect 21364 8774 21416 8780
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 21178 7712 21234 7721
rect 21178 7647 21234 7656
rect 21192 7274 21220 7647
rect 21284 7410 21312 7958
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 21284 7002 21312 7346
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21376 5817 21404 8774
rect 21362 5808 21418 5817
rect 21362 5743 21418 5752
rect 21468 5658 21496 11766
rect 21560 7313 21588 14758
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 21640 13864 21692 13870
rect 21640 13806 21692 13812
rect 21652 11830 21680 13806
rect 21822 13152 21878 13161
rect 21822 13087 21878 13096
rect 21730 13016 21786 13025
rect 21730 12951 21786 12960
rect 21640 11824 21692 11830
rect 21640 11766 21692 11772
rect 21744 11642 21772 12951
rect 21836 12442 21864 13087
rect 21824 12436 21876 12442
rect 21824 12378 21876 12384
rect 21836 11801 21864 12378
rect 22100 12368 22152 12374
rect 22100 12310 22152 12316
rect 22112 11898 22140 12310
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 21822 11792 21878 11801
rect 21822 11727 21878 11736
rect 21652 11614 21772 11642
rect 21546 7304 21602 7313
rect 21546 7239 21602 7248
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21560 6662 21588 7142
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21560 5914 21588 6598
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 20812 4820 20864 4826
rect 20812 4762 20864 4768
rect 20916 4814 21036 4842
rect 21284 5630 21496 5658
rect 20718 4312 20774 4321
rect 20718 4247 20774 4256
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20548 3942 20576 4014
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20548 3369 20576 3878
rect 20732 3738 20760 3878
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20916 3670 20944 4814
rect 20996 4752 21048 4758
rect 20996 4694 21048 4700
rect 20904 3664 20956 3670
rect 20626 3632 20682 3641
rect 20904 3606 20956 3612
rect 20626 3567 20682 3576
rect 20534 3360 20590 3369
rect 20534 3295 20590 3304
rect 20350 2816 20406 2825
rect 19622 2748 19918 2768
rect 20350 2751 20406 2760
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19444 2638 19564 2666
rect 18880 1692 18932 1698
rect 18880 1634 18932 1640
rect 18892 480 18920 1634
rect 19536 480 19564 2638
rect 20074 1864 20130 1873
rect 20074 1799 20130 1808
rect 20088 480 20116 1799
rect 20640 480 20668 3567
rect 20718 3224 20774 3233
rect 20916 3194 20944 3606
rect 21008 3602 21036 4694
rect 21180 3936 21232 3942
rect 21178 3904 21180 3913
rect 21232 3904 21234 3913
rect 21178 3839 21234 3848
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 21284 3466 21312 5630
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21468 3777 21496 5510
rect 21548 5364 21600 5370
rect 21548 5306 21600 5312
rect 21454 3768 21510 3777
rect 21364 3732 21416 3738
rect 21454 3703 21510 3712
rect 21364 3674 21416 3680
rect 21376 3641 21404 3674
rect 21362 3632 21418 3641
rect 21362 3567 21418 3576
rect 21456 3528 21508 3534
rect 21454 3496 21456 3505
rect 21508 3496 21510 3505
rect 21272 3460 21324 3466
rect 21454 3431 21510 3440
rect 21272 3402 21324 3408
rect 21468 3194 21496 3431
rect 20718 3159 20774 3168
rect 20904 3188 20956 3194
rect 20732 2922 20760 3159
rect 20904 3130 20956 3136
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 20732 2650 20760 2858
rect 20904 2848 20956 2854
rect 20904 2790 20956 2796
rect 20916 2650 20944 2790
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 21560 610 21588 5306
rect 21652 4826 21680 11614
rect 21732 11552 21784 11558
rect 21836 11540 21864 11727
rect 21916 11552 21968 11558
rect 21836 11512 21916 11540
rect 21732 11494 21784 11500
rect 21916 11494 21968 11500
rect 21744 11354 21772 11494
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 22112 11286 22140 11834
rect 22100 11280 22152 11286
rect 21730 11248 21786 11257
rect 22100 11222 22152 11228
rect 21730 11183 21786 11192
rect 21744 8838 21772 11183
rect 21914 11112 21970 11121
rect 21914 11047 21970 11056
rect 21928 10266 21956 11047
rect 22100 11008 22152 11014
rect 22100 10950 22152 10956
rect 22112 10266 22140 10950
rect 21916 10260 21968 10266
rect 21916 10202 21968 10208
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 22008 9716 22060 9722
rect 22008 9658 22060 9664
rect 21824 9648 21876 9654
rect 21824 9590 21876 9596
rect 21732 8832 21784 8838
rect 21732 8774 21784 8780
rect 21732 8560 21784 8566
rect 21730 8528 21732 8537
rect 21784 8528 21786 8537
rect 21730 8463 21786 8472
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 21744 6118 21772 6190
rect 21732 6112 21784 6118
rect 21732 6054 21784 6060
rect 21744 5166 21772 6054
rect 21732 5160 21784 5166
rect 21732 5102 21784 5108
rect 21640 4820 21692 4826
rect 21640 4762 21692 4768
rect 21652 4282 21680 4762
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 21836 3369 21864 9590
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 21928 9081 21956 9454
rect 21914 9072 21970 9081
rect 21914 9007 21970 9016
rect 22020 7324 22048 9658
rect 22112 9654 22140 10202
rect 22100 9648 22152 9654
rect 22100 9590 22152 9596
rect 22020 7296 22140 7324
rect 22006 7168 22062 7177
rect 22006 7103 22062 7112
rect 22020 6633 22048 7103
rect 22006 6624 22062 6633
rect 22006 6559 22062 6568
rect 21916 6112 21968 6118
rect 21916 6054 21968 6060
rect 21928 4758 21956 6054
rect 22112 5914 22140 7296
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 22008 5636 22060 5642
rect 22008 5578 22060 5584
rect 22020 5030 22048 5578
rect 22008 5024 22060 5030
rect 22008 4966 22060 4972
rect 21916 4752 21968 4758
rect 21916 4694 21968 4700
rect 22020 4690 22048 4966
rect 22008 4684 22060 4690
rect 22008 4626 22060 4632
rect 21916 4140 21968 4146
rect 21916 4082 21968 4088
rect 21928 3738 21956 4082
rect 22020 4026 22048 4626
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22112 4026 22140 4082
rect 22020 3998 22140 4026
rect 21916 3732 21968 3738
rect 21916 3674 21968 3680
rect 21822 3360 21878 3369
rect 21822 3295 21878 3304
rect 21928 3126 21956 3674
rect 21916 3120 21968 3126
rect 21822 3088 21878 3097
rect 21916 3062 21968 3068
rect 21822 3023 21878 3032
rect 21272 604 21324 610
rect 21272 546 21324 552
rect 21548 604 21600 610
rect 21548 546 21600 552
rect 21284 480 21312 546
rect 21836 480 21864 3023
rect 21928 2582 21956 3062
rect 22020 2650 22048 3998
rect 22204 3738 22232 14010
rect 22296 13025 22324 15438
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22374 13832 22430 13841
rect 22374 13767 22430 13776
rect 22282 13016 22338 13025
rect 22282 12951 22338 12960
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 22296 11694 22324 12242
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22296 11354 22324 11630
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22284 11212 22336 11218
rect 22284 11154 22336 11160
rect 22296 10538 22324 11154
rect 22284 10532 22336 10538
rect 22284 10474 22336 10480
rect 22296 10062 22324 10474
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 22284 8288 22336 8294
rect 22284 8230 22336 8236
rect 22296 8090 22324 8230
rect 22284 8084 22336 8090
rect 22284 8026 22336 8032
rect 22388 6610 22416 13767
rect 22480 11082 22508 15302
rect 22834 14920 22890 14929
rect 22834 14855 22890 14864
rect 22744 14816 22796 14822
rect 22744 14758 22796 14764
rect 22560 14476 22612 14482
rect 22560 14418 22612 14424
rect 22572 14113 22600 14418
rect 22558 14104 22614 14113
rect 22558 14039 22560 14048
rect 22612 14039 22614 14048
rect 22560 14010 22612 14016
rect 22572 13979 22600 14010
rect 22652 13728 22704 13734
rect 22652 13670 22704 13676
rect 22558 12880 22614 12889
rect 22558 12815 22614 12824
rect 22572 12782 22600 12815
rect 22560 12776 22612 12782
rect 22560 12718 22612 12724
rect 22468 11076 22520 11082
rect 22468 11018 22520 11024
rect 22468 10600 22520 10606
rect 22468 10542 22520 10548
rect 22480 9625 22508 10542
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22572 10130 22600 10406
rect 22560 10124 22612 10130
rect 22560 10066 22612 10072
rect 22664 9722 22692 13670
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22466 9616 22522 9625
rect 22466 9551 22522 9560
rect 22560 8288 22612 8294
rect 22560 8230 22612 8236
rect 22572 7546 22600 8230
rect 22756 8090 22784 14758
rect 22848 11286 22876 14855
rect 23204 14816 23256 14822
rect 23204 14758 23256 14764
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 22836 11280 22888 11286
rect 22836 11222 22888 11228
rect 22836 10056 22888 10062
rect 22836 9998 22888 10004
rect 22848 9722 22876 9998
rect 22836 9716 22888 9722
rect 22836 9658 22888 9664
rect 22848 9042 22876 9658
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 22744 8084 22796 8090
rect 22744 8026 22796 8032
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 22572 7002 22600 7482
rect 22756 7342 22784 8026
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 22560 6996 22612 7002
rect 22560 6938 22612 6944
rect 22744 6656 22796 6662
rect 22388 6582 22508 6610
rect 22744 6598 22796 6604
rect 22376 5772 22428 5778
rect 22376 5714 22428 5720
rect 22388 4826 22416 5714
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 22284 4616 22336 4622
rect 22284 4558 22336 4564
rect 22296 4010 22324 4558
rect 22480 4078 22508 6582
rect 22756 6322 22784 6598
rect 22744 6316 22796 6322
rect 22744 6258 22796 6264
rect 22756 5574 22784 6258
rect 22744 5568 22796 5574
rect 22744 5510 22796 5516
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22664 4185 22692 4966
rect 22756 4690 22784 5510
rect 22940 5370 22968 14214
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 23032 8401 23060 13806
rect 23112 13320 23164 13326
rect 23112 13262 23164 13268
rect 23124 10606 23152 13262
rect 23112 10600 23164 10606
rect 23112 10542 23164 10548
rect 23124 10266 23152 10542
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 23124 9586 23152 10066
rect 23216 9636 23244 14758
rect 23308 10810 23336 16238
rect 23492 14770 23520 17031
rect 23584 14890 23612 26823
rect 24030 26208 24086 26217
rect 24030 26143 24086 26152
rect 23848 22092 23900 22098
rect 23848 22034 23900 22040
rect 23860 21486 23888 22034
rect 23848 21480 23900 21486
rect 23846 21448 23848 21457
rect 23940 21480 23992 21486
rect 23900 21448 23902 21457
rect 23940 21422 23992 21428
rect 23846 21383 23902 21392
rect 23664 17128 23716 17134
rect 23664 17070 23716 17076
rect 23572 14884 23624 14890
rect 23572 14826 23624 14832
rect 23400 14742 23520 14770
rect 23400 14498 23428 14742
rect 23400 14470 23520 14498
rect 23492 13394 23520 14470
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 23584 13870 23612 14418
rect 23572 13864 23624 13870
rect 23572 13806 23624 13812
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23492 12986 23520 13330
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23478 12744 23534 12753
rect 23478 12679 23534 12688
rect 23492 11257 23520 12679
rect 23478 11248 23534 11257
rect 23478 11183 23534 11192
rect 23296 10804 23348 10810
rect 23296 10746 23348 10752
rect 23480 9648 23532 9654
rect 23216 9608 23480 9636
rect 23480 9590 23532 9596
rect 23112 9580 23164 9586
rect 23112 9522 23164 9528
rect 23124 9178 23152 9522
rect 23112 9172 23164 9178
rect 23112 9114 23164 9120
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23018 8392 23074 8401
rect 23018 8327 23074 8336
rect 23112 7336 23164 7342
rect 23112 7278 23164 7284
rect 23124 6458 23152 7278
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 22928 5364 22980 5370
rect 22928 5306 22980 5312
rect 22940 5166 22968 5306
rect 22928 5160 22980 5166
rect 22928 5102 22980 5108
rect 22744 4684 22796 4690
rect 22744 4626 22796 4632
rect 22756 4282 22784 4626
rect 22744 4276 22796 4282
rect 22744 4218 22796 4224
rect 22650 4176 22706 4185
rect 22650 4111 22706 4120
rect 22468 4072 22520 4078
rect 22468 4014 22520 4020
rect 22284 4004 22336 4010
rect 22284 3946 22336 3952
rect 22480 3738 22508 4014
rect 23216 3942 23244 8910
rect 23480 8356 23532 8362
rect 23480 8298 23532 8304
rect 23492 7449 23520 8298
rect 23478 7440 23534 7449
rect 23478 7375 23534 7384
rect 23478 7304 23534 7313
rect 23478 7239 23480 7248
rect 23532 7239 23534 7248
rect 23480 7210 23532 7216
rect 23296 7200 23348 7206
rect 23296 7142 23348 7148
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 22468 3732 22520 3738
rect 22468 3674 22520 3680
rect 22664 3505 22692 3878
rect 22650 3496 22706 3505
rect 22650 3431 22706 3440
rect 22652 3392 22704 3398
rect 22374 3360 22430 3369
rect 22652 3334 22704 3340
rect 22374 3295 22430 3304
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 21916 2576 21968 2582
rect 21916 2518 21968 2524
rect 22388 480 22416 3295
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 22572 2650 22600 3130
rect 22664 2825 22692 3334
rect 23308 3108 23336 7142
rect 23388 6248 23440 6254
rect 23440 6208 23520 6236
rect 23388 6190 23440 6196
rect 23492 5137 23520 6208
rect 23478 5128 23534 5137
rect 23478 5063 23534 5072
rect 23584 4264 23612 13806
rect 23676 13705 23704 17070
rect 23848 16652 23900 16658
rect 23848 16594 23900 16600
rect 23860 16046 23888 16594
rect 23952 16561 23980 21422
rect 23938 16552 23994 16561
rect 23938 16487 23994 16496
rect 23848 16040 23900 16046
rect 23846 16008 23848 16017
rect 23900 16008 23902 16017
rect 23846 15943 23902 15952
rect 23848 15904 23900 15910
rect 23848 15846 23900 15852
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 23768 13841 23796 14214
rect 23754 13832 23810 13841
rect 23754 13767 23810 13776
rect 23662 13696 23718 13705
rect 23662 13631 23718 13640
rect 23860 13326 23888 15846
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 23952 14822 23980 15506
rect 23940 14816 23992 14822
rect 23940 14758 23992 14764
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 23846 13152 23902 13161
rect 23846 13087 23902 13096
rect 23860 11354 23888 13087
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23952 11234 23980 14758
rect 24044 12442 24072 26143
rect 25226 25528 25282 25537
rect 25226 25463 25282 25472
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24766 24848 24822 24857
rect 24766 24783 24822 24792
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24780 23322 24808 24783
rect 24768 23316 24820 23322
rect 24768 23258 24820 23264
rect 24766 23216 24822 23225
rect 24676 23180 24728 23186
rect 24766 23151 24822 23160
rect 24676 23122 24728 23128
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24688 22658 24716 23122
rect 24596 22630 24716 22658
rect 24596 22438 24624 22630
rect 24674 22536 24730 22545
rect 24674 22471 24730 22480
rect 24584 22432 24636 22438
rect 24584 22374 24636 22380
rect 24596 22234 24624 22374
rect 24584 22228 24636 22234
rect 24584 22170 24636 22176
rect 24124 22092 24176 22098
rect 24124 22034 24176 22040
rect 24136 21350 24164 22034
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24688 21690 24716 22471
rect 24780 21962 24808 23151
rect 24768 21956 24820 21962
rect 24768 21898 24820 21904
rect 24676 21684 24728 21690
rect 24676 21626 24728 21632
rect 24674 21448 24730 21457
rect 24674 21383 24730 21392
rect 24124 21344 24176 21350
rect 24124 21286 24176 21292
rect 24136 19961 24164 21286
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24122 19952 24178 19961
rect 24122 19887 24178 19896
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24214 18728 24270 18737
rect 24214 18663 24270 18672
rect 24228 17338 24256 18663
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 18193 24716 21383
rect 24766 19408 24822 19417
rect 24766 19343 24822 19352
rect 24674 18184 24730 18193
rect 24674 18119 24730 18128
rect 24780 17882 24808 19343
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 24766 17776 24822 17785
rect 24676 17740 24728 17746
rect 24766 17711 24822 17720
rect 24676 17682 24728 17688
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24216 17332 24268 17338
rect 24216 17274 24268 17280
rect 24688 17218 24716 17682
rect 24412 17190 24716 17218
rect 24412 16998 24440 17190
rect 24674 17096 24730 17105
rect 24674 17031 24730 17040
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24412 16794 24440 16934
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 24214 16688 24270 16697
rect 24124 16652 24176 16658
rect 24214 16623 24270 16632
rect 24124 16594 24176 16600
rect 24136 16425 24164 16594
rect 24122 16416 24178 16425
rect 24122 16351 24178 16360
rect 24136 16250 24164 16351
rect 24124 16244 24176 16250
rect 24124 16186 24176 16192
rect 24122 15192 24178 15201
rect 24122 15127 24178 15136
rect 24136 14958 24164 15127
rect 24124 14952 24176 14958
rect 24124 14894 24176 14900
rect 24124 14816 24176 14822
rect 24124 14758 24176 14764
rect 24136 13433 24164 14758
rect 24228 14618 24256 16623
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24688 15706 24716 17031
rect 24780 16794 24808 17711
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24766 16008 24822 16017
rect 24766 15943 24822 15952
rect 24676 15700 24728 15706
rect 24676 15642 24728 15648
rect 24674 15328 24730 15337
rect 24289 15260 24585 15280
rect 24674 15263 24730 15272
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 14634 24716 15263
rect 24780 15162 24808 15943
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24872 14822 24900 15506
rect 24952 14884 25004 14890
rect 24952 14826 25004 14832
rect 24860 14816 24912 14822
rect 24860 14758 24912 14764
rect 24216 14612 24268 14618
rect 24688 14606 24808 14634
rect 24216 14554 24268 14560
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24582 13968 24638 13977
rect 24582 13903 24638 13912
rect 24596 13870 24624 13903
rect 24584 13864 24636 13870
rect 24584 13806 24636 13812
rect 24688 13734 24716 14418
rect 24780 14090 24808 14606
rect 24780 14062 24900 14090
rect 24768 14000 24820 14006
rect 24766 13968 24768 13977
rect 24820 13968 24822 13977
rect 24766 13903 24822 13912
rect 24872 13852 24900 14062
rect 24780 13824 24900 13852
rect 24400 13728 24452 13734
rect 24400 13670 24452 13676
rect 24676 13728 24728 13734
rect 24676 13670 24728 13676
rect 24412 13530 24440 13670
rect 24780 13530 24808 13824
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24768 13524 24820 13530
rect 24768 13466 24820 13472
rect 24122 13424 24178 13433
rect 24122 13359 24178 13368
rect 24216 13388 24268 13394
rect 24216 13330 24268 13336
rect 24228 12918 24256 13330
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24216 12912 24268 12918
rect 24216 12854 24268 12860
rect 24124 12776 24176 12782
rect 24124 12718 24176 12724
rect 24032 12436 24084 12442
rect 24032 12378 24084 12384
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 24044 11626 24072 12038
rect 24032 11620 24084 11626
rect 24032 11562 24084 11568
rect 23860 11206 23980 11234
rect 23756 10532 23808 10538
rect 23756 10474 23808 10480
rect 23664 10464 23716 10470
rect 23664 10406 23716 10412
rect 23676 10198 23704 10406
rect 23664 10192 23716 10198
rect 23664 10134 23716 10140
rect 23676 9518 23704 10134
rect 23664 9512 23716 9518
rect 23768 9489 23796 10474
rect 23664 9454 23716 9460
rect 23754 9480 23810 9489
rect 23754 9415 23810 9424
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 23662 8392 23718 8401
rect 23662 8327 23718 8336
rect 23676 7546 23704 8327
rect 23768 8090 23796 8978
rect 23860 8378 23888 11206
rect 24044 11150 24072 11562
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 24136 10538 24164 12718
rect 24676 12300 24728 12306
rect 24676 12242 24728 12248
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11812 24716 12242
rect 24596 11784 24716 11812
rect 24596 11150 24624 11784
rect 24676 11280 24728 11286
rect 24676 11222 24728 11228
rect 24584 11144 24636 11150
rect 24582 11112 24584 11121
rect 24636 11112 24638 11121
rect 24582 11047 24638 11056
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10810 24716 11222
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24674 10704 24730 10713
rect 24308 10668 24360 10674
rect 24674 10639 24730 10648
rect 24308 10610 24360 10616
rect 24124 10532 24176 10538
rect 24124 10474 24176 10480
rect 24320 10130 24348 10610
rect 24308 10124 24360 10130
rect 24308 10066 24360 10072
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24122 9208 24178 9217
rect 24122 9143 24178 9152
rect 24030 8528 24086 8537
rect 24030 8463 24086 8472
rect 23860 8350 23980 8378
rect 23848 8288 23900 8294
rect 23848 8230 23900 8236
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 23768 7546 23796 8026
rect 23664 7540 23716 7546
rect 23664 7482 23716 7488
rect 23756 7540 23808 7546
rect 23756 7482 23808 7488
rect 23662 6896 23718 6905
rect 23768 6866 23796 7482
rect 23860 7410 23888 8230
rect 23848 7404 23900 7410
rect 23848 7346 23900 7352
rect 23860 7002 23888 7346
rect 23848 6996 23900 7002
rect 23848 6938 23900 6944
rect 23662 6831 23718 6840
rect 23756 6860 23808 6866
rect 23676 5817 23704 6831
rect 23756 6802 23808 6808
rect 23768 6458 23796 6802
rect 23756 6452 23808 6458
rect 23756 6394 23808 6400
rect 23768 5846 23796 6394
rect 23756 5840 23808 5846
rect 23662 5808 23718 5817
rect 23756 5782 23808 5788
rect 23662 5743 23718 5752
rect 23952 5642 23980 8350
rect 23940 5636 23992 5642
rect 23940 5578 23992 5584
rect 24044 5409 24072 8463
rect 24136 7721 24164 9143
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24492 8492 24544 8498
rect 24492 8434 24544 8440
rect 24504 8022 24532 8434
rect 24688 8430 24716 10639
rect 24780 10010 24808 13262
rect 24964 12986 24992 14826
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 24950 12608 25006 12617
rect 24950 12543 25006 12552
rect 24860 11552 24912 11558
rect 24860 11494 24912 11500
rect 24872 10674 24900 11494
rect 24964 11286 24992 12543
rect 25042 12336 25098 12345
rect 25042 12271 25098 12280
rect 24952 11280 25004 11286
rect 24952 11222 25004 11228
rect 25056 11218 25084 12271
rect 25240 11354 25268 25463
rect 25502 24168 25558 24177
rect 25502 24103 25558 24112
rect 25410 22128 25466 22137
rect 25410 22063 25466 22072
rect 25318 18184 25374 18193
rect 25318 18119 25374 18128
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 25044 11212 25096 11218
rect 25044 11154 25096 11160
rect 25056 10810 25084 11154
rect 25044 10804 25096 10810
rect 25044 10746 25096 10752
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 25228 10600 25280 10606
rect 25228 10542 25280 10548
rect 25240 10169 25268 10542
rect 25226 10160 25282 10169
rect 25226 10095 25282 10104
rect 25226 10024 25282 10033
rect 24780 9982 24992 10010
rect 24768 9920 24820 9926
rect 24768 9862 24820 9868
rect 24780 9518 24808 9862
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 24780 9364 24808 9454
rect 24860 9376 24912 9382
rect 24780 9336 24860 9364
rect 24780 9110 24808 9336
rect 24860 9318 24912 9324
rect 24768 9104 24820 9110
rect 24768 9046 24820 9052
rect 24872 8634 24900 9318
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24676 8424 24728 8430
rect 24676 8366 24728 8372
rect 24492 8016 24544 8022
rect 24492 7958 24544 7964
rect 24766 7848 24822 7857
rect 24766 7783 24822 7792
rect 24676 7744 24728 7750
rect 24122 7712 24178 7721
rect 24676 7686 24728 7692
rect 24122 7647 24178 7656
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24688 7410 24716 7686
rect 24676 7404 24728 7410
rect 24676 7346 24728 7352
rect 24688 6934 24716 7346
rect 24676 6928 24728 6934
rect 24676 6870 24728 6876
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24400 6248 24452 6254
rect 24214 6216 24270 6225
rect 24400 6190 24452 6196
rect 24214 6151 24270 6160
rect 24030 5400 24086 5409
rect 24030 5335 24086 5344
rect 24228 5302 24256 6151
rect 24412 5914 24440 6190
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 24676 5908 24728 5914
rect 24676 5850 24728 5856
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24216 5296 24268 5302
rect 24216 5238 24268 5244
rect 24228 5098 24256 5238
rect 24688 5234 24716 5850
rect 24780 5794 24808 7783
rect 24964 5914 24992 9982
rect 25226 9959 25282 9968
rect 25240 9518 25268 9959
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 25148 8634 25176 8774
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25148 7546 25176 8570
rect 25332 7546 25360 18119
rect 25424 9654 25452 22063
rect 25516 10810 25544 24103
rect 25594 20768 25650 20777
rect 25594 20703 25650 20712
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25412 9648 25464 9654
rect 25412 9590 25464 9596
rect 25608 8634 25636 20703
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 25412 8424 25464 8430
rect 25412 8366 25464 8372
rect 25424 7993 25452 8366
rect 25410 7984 25466 7993
rect 25410 7919 25466 7928
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 25226 7440 25282 7449
rect 25226 7375 25282 7384
rect 25240 7342 25268 7375
rect 25228 7336 25280 7342
rect 25228 7278 25280 7284
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25148 6254 25176 6598
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 25136 6112 25188 6118
rect 25136 6054 25188 6060
rect 24952 5908 25004 5914
rect 24952 5850 25004 5856
rect 24780 5766 24900 5794
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 24780 5370 24808 5646
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24676 5228 24728 5234
rect 24676 5170 24728 5176
rect 24872 5166 24900 5766
rect 24964 5370 24992 5850
rect 25148 5710 25176 6054
rect 25136 5704 25188 5710
rect 25136 5646 25188 5652
rect 24952 5364 25004 5370
rect 24952 5306 25004 5312
rect 24860 5160 24912 5166
rect 24780 5120 24860 5148
rect 24216 5092 24268 5098
rect 24216 5034 24268 5040
rect 24780 4826 24808 5120
rect 24860 5102 24912 5108
rect 24950 4992 25006 5001
rect 24950 4927 25006 4936
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 24964 4690 24992 4927
rect 25148 4758 25176 5646
rect 25136 4752 25188 4758
rect 25136 4694 25188 4700
rect 24952 4684 25004 4690
rect 24952 4626 25004 4632
rect 23848 4480 23900 4486
rect 23848 4422 23900 4428
rect 23754 4312 23810 4321
rect 23584 4236 23704 4264
rect 23754 4247 23810 4256
rect 23572 4140 23624 4146
rect 23572 4082 23624 4088
rect 23584 3602 23612 4082
rect 23676 4078 23704 4236
rect 23664 4072 23716 4078
rect 23664 4014 23716 4020
rect 23662 3904 23718 3913
rect 23662 3839 23718 3848
rect 23572 3596 23624 3602
rect 23572 3538 23624 3544
rect 23584 3194 23612 3538
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 23308 3080 23520 3108
rect 23492 3074 23520 3080
rect 23492 3046 23612 3074
rect 23480 2848 23532 2854
rect 22650 2816 22706 2825
rect 23480 2790 23532 2796
rect 22650 2751 22706 2760
rect 23018 2680 23074 2689
rect 22560 2644 22612 2650
rect 23018 2615 23074 2624
rect 22560 2586 22612 2592
rect 23032 480 23060 2615
rect 23492 2145 23520 2790
rect 23478 2136 23534 2145
rect 23478 2071 23534 2080
rect 23584 480 23612 3046
rect 23676 1057 23704 3839
rect 23768 2650 23796 4247
rect 23860 4010 23888 4422
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24964 4282 24992 4626
rect 27068 4480 27120 4486
rect 27068 4422 27120 4428
rect 24952 4276 25004 4282
rect 24952 4218 25004 4224
rect 25318 4176 25374 4185
rect 25136 4140 25188 4146
rect 25318 4111 25374 4120
rect 25136 4082 25188 4088
rect 24032 4072 24084 4078
rect 24032 4014 24084 4020
rect 23848 4004 23900 4010
rect 23848 3946 23900 3952
rect 23860 3670 23888 3946
rect 24044 3942 24072 4014
rect 24216 4004 24268 4010
rect 24216 3946 24268 3952
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 24122 3904 24178 3913
rect 24122 3839 24178 3848
rect 23938 3768 23994 3777
rect 23938 3703 23994 3712
rect 23848 3664 23900 3670
rect 23848 3606 23900 3612
rect 23860 3126 23888 3606
rect 23848 3120 23900 3126
rect 23848 3062 23900 3068
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 23952 2281 23980 3703
rect 24030 3224 24086 3233
rect 24030 3159 24032 3168
rect 24084 3159 24086 3168
rect 24032 3130 24084 3136
rect 24030 3088 24086 3097
rect 24030 3023 24086 3032
rect 24044 2854 24072 3023
rect 24032 2848 24084 2854
rect 24032 2790 24084 2796
rect 23938 2272 23994 2281
rect 23938 2207 23994 2216
rect 23662 1048 23718 1057
rect 23662 983 23718 992
rect 24136 480 24164 3839
rect 24228 2650 24256 3946
rect 25148 3942 25176 4082
rect 25136 3936 25188 3942
rect 25136 3878 25188 3884
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24780 2990 24808 3334
rect 25148 3194 25176 3878
rect 25136 3188 25188 3194
rect 25136 3130 25188 3136
rect 24768 2984 24820 2990
rect 24582 2952 24638 2961
rect 24768 2926 24820 2932
rect 24582 2887 24638 2896
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 24492 2440 24544 2446
rect 24490 2408 24492 2417
rect 24544 2408 24546 2417
rect 24596 2394 24624 2887
rect 24780 2446 24808 2926
rect 24768 2440 24820 2446
rect 24596 2366 24716 2394
rect 24768 2382 24820 2388
rect 24490 2343 24546 2352
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24688 1442 24716 2366
rect 24688 1414 24808 1442
rect 24780 480 24808 1414
rect 25332 480 25360 4111
rect 26054 3632 26110 3641
rect 26054 3567 26110 3576
rect 25870 3496 25926 3505
rect 25870 3431 25926 3440
rect 25884 480 25912 3431
rect 26068 3194 26096 3567
rect 26056 3188 26108 3194
rect 26056 3130 26108 3136
rect 26514 2816 26570 2825
rect 26514 2751 26570 2760
rect 26528 480 26556 2751
rect 27080 480 27108 4422
rect 27618 4040 27674 4049
rect 27618 3975 27674 3984
rect 27632 480 27660 3975
rect 18786 368 18842 377
rect 18786 303 18842 312
rect 18878 0 18934 480
rect 19522 0 19578 480
rect 20074 0 20130 480
rect 20626 0 20682 480
rect 21270 0 21326 480
rect 21822 0 21878 480
rect 22374 0 22430 480
rect 23018 0 23074 480
rect 23570 0 23626 480
rect 24122 0 24178 480
rect 24766 0 24822 480
rect 25318 0 25374 480
rect 25870 0 25926 480
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 2778 27512 2834 27568
rect 1950 26152 2006 26208
rect 1582 24792 1638 24848
rect 1582 22072 1638 22128
rect 1490 21392 1546 21448
rect 1398 20712 1454 20768
rect 1858 20712 1914 20768
rect 1582 20032 1638 20088
rect 1490 18672 1546 18728
rect 1398 17312 1454 17368
rect 1674 19352 1730 19408
rect 1582 17992 1638 18048
rect 1582 15952 1638 16008
rect 1490 14592 1546 14648
rect 2226 24112 2282 24168
rect 2042 23432 2098 23488
rect 2042 20712 2098 20768
rect 2042 18028 2044 18048
rect 2044 18028 2096 18048
rect 2096 18028 2098 18048
rect 2042 17992 2098 18028
rect 2134 17176 2190 17232
rect 1950 16632 2006 16688
rect 1674 15272 1730 15328
rect 1582 13912 1638 13968
rect 846 2760 902 2816
rect 2042 14864 2098 14920
rect 2410 19236 2466 19272
rect 2410 19216 2412 19236
rect 2412 19216 2464 19236
rect 2464 19216 2466 19236
rect 2410 18828 2466 18864
rect 2410 18808 2412 18828
rect 2412 18808 2464 18828
rect 2464 18808 2466 18828
rect 2502 18672 2558 18728
rect 2042 13812 2044 13832
rect 2044 13812 2096 13832
rect 2096 13812 2098 13832
rect 2042 13776 2098 13812
rect 2042 12724 2044 12744
rect 2044 12724 2096 12744
rect 2096 12724 2098 12744
rect 2042 12688 2098 12724
rect 1582 6724 1638 6760
rect 1582 6704 1584 6724
rect 1584 6704 1636 6724
rect 1636 6704 1638 6724
rect 1398 5888 1454 5944
rect 1490 5072 1546 5128
rect 1674 4664 1730 4720
rect 2042 10668 2098 10704
rect 2042 10648 2044 10668
rect 2044 10648 2096 10668
rect 2096 10648 2098 10668
rect 2410 15408 2466 15464
rect 3054 26832 3110 26888
rect 2870 25472 2926 25528
rect 2226 12416 2282 12472
rect 2962 22752 3018 22808
rect 2410 10260 2466 10296
rect 2410 10240 2412 10260
rect 2412 10240 2464 10260
rect 2464 10240 2466 10260
rect 2686 11620 2742 11656
rect 2686 11600 2688 11620
rect 2688 11600 2740 11620
rect 2740 11600 2742 11620
rect 2594 11500 2596 11520
rect 2596 11500 2648 11520
rect 2648 11500 2650 11520
rect 2594 11464 2650 11500
rect 2870 13096 2926 13152
rect 2318 8064 2374 8120
rect 2502 8356 2558 8392
rect 2502 8336 2504 8356
rect 2504 8336 2556 8356
rect 2556 8336 2558 8356
rect 2226 7964 2228 7984
rect 2228 7964 2280 7984
rect 2280 7964 2282 7984
rect 2226 7928 2282 7964
rect 1858 7656 1914 7712
rect 2042 5616 2098 5672
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 10874 21392 10930 21448
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 9678 18808 9734 18864
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 9126 17992 9182 18048
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 8022 16904 8078 16960
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 7654 15952 7710 16008
rect 4894 15408 4950 15464
rect 3422 12552 3478 12608
rect 2778 10124 2834 10160
rect 2778 10104 2780 10124
rect 2780 10104 2832 10124
rect 2832 10104 2834 10124
rect 3054 8472 3110 8528
rect 2962 7928 3018 7984
rect 2502 6160 2558 6216
rect 1858 2932 1860 2952
rect 1860 2932 1912 2952
rect 1912 2932 1914 2952
rect 1858 2896 1914 2932
rect 1950 2488 2006 2544
rect 3698 10512 3754 10568
rect 4710 13912 4766 13968
rect 4802 13232 4858 13288
rect 4710 13096 4766 13152
rect 3422 9560 3478 9616
rect 2318 2624 2374 2680
rect 2778 3712 2834 3768
rect 3146 3712 3202 3768
rect 3054 2896 3110 2952
rect 2962 992 3018 1048
rect 3514 8336 3570 8392
rect 3698 8200 3754 8256
rect 3698 6840 3754 6896
rect 4066 10648 4122 10704
rect 4526 10240 4582 10296
rect 4250 7792 4306 7848
rect 4434 7404 4490 7440
rect 4434 7384 4436 7404
rect 4436 7384 4488 7404
rect 4488 7384 4490 7404
rect 4526 5616 4582 5672
rect 4066 5072 4122 5128
rect 3422 3032 3478 3088
rect 4710 8064 4766 8120
rect 4710 7248 4766 7304
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 6918 14184 6974 14240
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5998 13368 6054 13424
rect 5998 13096 6054 13152
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 6734 12824 6790 12880
rect 4986 12708 5042 12744
rect 4986 12688 4988 12708
rect 4988 12688 5040 12708
rect 5040 12688 5042 12708
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5538 11464 5594 11520
rect 6182 11500 6184 11520
rect 6184 11500 6236 11520
rect 6236 11500 6238 11520
rect 6182 11464 6238 11500
rect 4894 7384 4950 7440
rect 3422 1536 3478 1592
rect 3698 1264 3754 1320
rect 5262 10104 5318 10160
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 6090 10956 6092 10976
rect 6092 10956 6144 10976
rect 6144 10956 6146 10976
rect 6090 10920 6146 10956
rect 5538 10548 5540 10568
rect 5540 10548 5592 10568
rect 5592 10548 5594 10568
rect 5538 10512 5594 10548
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5170 7656 5226 7712
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5078 3848 5134 3904
rect 4618 1944 4674 2000
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 6090 6024 6146 6080
rect 5998 4800 6054 4856
rect 5446 4428 5448 4448
rect 5448 4428 5500 4448
rect 5500 4428 5502 4448
rect 5446 4392 5502 4428
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 6090 3712 6146 3768
rect 5354 3032 5410 3088
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5354 2760 5410 2816
rect 5630 2896 5686 2952
rect 5538 2760 5594 2816
rect 3698 312 3754 368
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6366 5344 6422 5400
rect 6182 2760 6238 2816
rect 7286 13368 7342 13424
rect 7194 9832 7250 9888
rect 6918 7384 6974 7440
rect 7010 6568 7066 6624
rect 6550 5208 6606 5264
rect 6642 4936 6698 4992
rect 6826 5616 6882 5672
rect 6734 3848 6790 3904
rect 7194 3712 7250 3768
rect 6918 2624 6974 2680
rect 6734 2216 6790 2272
rect 7838 15544 7894 15600
rect 7746 12280 7802 12336
rect 7562 10784 7618 10840
rect 7562 8336 7618 8392
rect 7746 7656 7802 7712
rect 7746 7112 7802 7168
rect 7470 5752 7526 5808
rect 7378 3984 7434 4040
rect 7654 3476 7656 3496
rect 7656 3476 7708 3496
rect 7708 3476 7710 3496
rect 7654 3440 7710 3476
rect 7470 2352 7526 2408
rect 8298 15000 8354 15056
rect 8850 12960 8906 13016
rect 8666 12552 8722 12608
rect 8574 12416 8630 12472
rect 8390 11756 8446 11792
rect 8390 11736 8392 11756
rect 8392 11736 8444 11756
rect 8444 11736 8446 11756
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10690 17040 10746 17096
rect 10138 16940 10140 16960
rect 10140 16940 10192 16960
rect 10192 16940 10194 16960
rect 10138 16904 10194 16940
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10138 16088 10194 16144
rect 10046 14048 10102 14104
rect 9310 13776 9366 13832
rect 9494 13368 9550 13424
rect 9218 11464 9274 11520
rect 8206 9288 8262 9344
rect 8758 10376 8814 10432
rect 8206 8880 8262 8936
rect 8114 8200 8170 8256
rect 8022 7384 8078 7440
rect 8114 6976 8170 7032
rect 8390 6296 8446 6352
rect 7930 4820 7986 4856
rect 7930 4800 7932 4820
rect 7932 4800 7984 4820
rect 7984 4800 7986 4820
rect 7930 4528 7986 4584
rect 8298 4684 8354 4720
rect 8298 4664 8300 4684
rect 8300 4664 8352 4684
rect 8352 4664 8354 4684
rect 8022 4392 8078 4448
rect 7930 3848 7986 3904
rect 8390 3168 8446 3224
rect 8942 10140 8944 10160
rect 8944 10140 8996 10160
rect 8996 10140 8998 10160
rect 8942 10104 8998 10140
rect 9310 10920 9366 10976
rect 9770 12280 9826 12336
rect 9494 12044 9496 12064
rect 9496 12044 9548 12064
rect 9548 12044 9550 12064
rect 9494 12008 9550 12044
rect 9586 11892 9642 11928
rect 9586 11872 9588 11892
rect 9588 11872 9640 11892
rect 9640 11872 9642 11892
rect 9494 11600 9550 11656
rect 9586 10104 9642 10160
rect 9402 9696 9458 9752
rect 9586 8744 9642 8800
rect 9402 8608 9458 8664
rect 8666 3712 8722 3768
rect 8206 3032 8262 3088
rect 8666 2080 8722 2136
rect 8298 1944 8354 2000
rect 9034 5208 9090 5264
rect 9218 7520 9274 7576
rect 9218 5616 9274 5672
rect 9218 5244 9220 5264
rect 9220 5244 9272 5264
rect 9272 5244 9274 5264
rect 9218 5208 9274 5244
rect 9126 4936 9182 4992
rect 8942 4528 8998 4584
rect 9034 3576 9090 3632
rect 9126 3440 9182 3496
rect 9402 8064 9458 8120
rect 9862 10240 9918 10296
rect 9862 9868 9864 9888
rect 9864 9868 9916 9888
rect 9916 9868 9918 9888
rect 9862 9832 9918 9868
rect 9770 8608 9826 8664
rect 9402 6432 9458 6488
rect 9770 7112 9826 7168
rect 9862 6976 9918 7032
rect 9678 6840 9734 6896
rect 9770 6740 9772 6760
rect 9772 6740 9824 6760
rect 9824 6740 9826 6760
rect 9770 6704 9826 6740
rect 9770 6024 9826 6080
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 11702 19216 11758 19272
rect 11058 16940 11060 16960
rect 11060 16940 11112 16960
rect 11112 16940 11114 16960
rect 11058 16904 11114 16940
rect 10966 15000 11022 15056
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10690 13504 10746 13560
rect 10230 13368 10286 13424
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10690 12008 10746 12064
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10230 10920 10286 10976
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10690 10240 10746 10296
rect 10690 9968 10746 10024
rect 10138 9424 10194 9480
rect 10138 9324 10140 9344
rect 10140 9324 10192 9344
rect 10192 9324 10194 9344
rect 10138 9288 10194 9324
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10414 8880 10470 8936
rect 10690 8880 10746 8936
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10506 7948 10562 7984
rect 10506 7928 10508 7948
rect 10508 7928 10560 7948
rect 10560 7928 10562 7948
rect 10046 6840 10102 6896
rect 10046 6024 10102 6080
rect 12438 18692 12494 18728
rect 12438 18672 12440 18692
rect 12440 18672 12492 18692
rect 12492 18672 12494 18692
rect 13266 17176 13322 17232
rect 10966 14320 11022 14376
rect 10966 13932 11022 13968
rect 10966 13912 10968 13932
rect 10968 13912 11020 13932
rect 11020 13912 11022 13932
rect 11150 12980 11206 13016
rect 11150 12960 11152 12980
rect 11152 12960 11204 12980
rect 11204 12960 11206 12980
rect 11426 13640 11482 13696
rect 11334 13232 11390 13288
rect 10966 12552 11022 12608
rect 11058 12280 11114 12336
rect 10966 12008 11022 12064
rect 10874 11192 10930 11248
rect 11150 10376 11206 10432
rect 10966 8880 11022 8936
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10966 6976 11022 7032
rect 11150 8336 11206 8392
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 9218 2896 9274 2952
rect 9770 3984 9826 4040
rect 9678 3304 9734 3360
rect 9678 3032 9734 3088
rect 9402 1400 9458 1456
rect 10782 6024 10838 6080
rect 10782 4936 10838 4992
rect 9770 2216 9826 2272
rect 10046 3304 10102 3360
rect 9862 1808 9918 1864
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10230 3440 10286 3496
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10874 1944 10930 2000
rect 12162 15544 12218 15600
rect 12714 16632 12770 16688
rect 11794 11872 11850 11928
rect 11702 10668 11758 10704
rect 11702 10648 11704 10668
rect 11704 10648 11756 10668
rect 11756 10648 11758 10668
rect 11702 9696 11758 9752
rect 11426 9288 11482 9344
rect 11150 3576 11206 3632
rect 11518 8472 11574 8528
rect 11426 5344 11482 5400
rect 11794 7656 11850 7712
rect 11426 4664 11482 4720
rect 11426 4392 11482 4448
rect 11426 3848 11482 3904
rect 11426 2896 11482 2952
rect 11242 2508 11298 2544
rect 11242 2488 11244 2508
rect 11244 2488 11296 2508
rect 11296 2488 11298 2508
rect 10690 1672 10746 1728
rect 11426 1536 11482 1592
rect 11794 3188 11850 3224
rect 11794 3168 11796 3188
rect 11796 3168 11848 3188
rect 11848 3168 11850 3188
rect 11702 2372 11758 2408
rect 11702 2352 11704 2372
rect 11704 2352 11756 2372
rect 11756 2352 11758 2372
rect 11610 1536 11666 1592
rect 10690 1128 10746 1184
rect 12346 14884 12402 14920
rect 12346 14864 12348 14884
rect 12348 14864 12400 14884
rect 12400 14864 12402 14884
rect 12438 13912 12494 13968
rect 12346 13096 12402 13152
rect 12162 12144 12218 12200
rect 11978 11600 12034 11656
rect 12070 10784 12126 10840
rect 12162 9832 12218 9888
rect 12162 9596 12164 9616
rect 12164 9596 12216 9616
rect 12216 9596 12218 9616
rect 12162 9560 12218 9596
rect 12162 6568 12218 6624
rect 12346 11328 12402 11384
rect 12438 9460 12440 9480
rect 12440 9460 12492 9480
rect 12492 9460 12494 9480
rect 12438 9424 12494 9460
rect 12622 11056 12678 11112
rect 12622 9560 12678 9616
rect 12622 8472 12678 8528
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14922 19216 14978 19272
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 12898 14184 12954 14240
rect 12438 7792 12494 7848
rect 12622 7384 12678 7440
rect 12162 3732 12218 3768
rect 12162 3712 12164 3732
rect 12164 3712 12216 3732
rect 12216 3712 12218 3732
rect 11978 2760 12034 2816
rect 12438 3068 12440 3088
rect 12440 3068 12492 3088
rect 12492 3068 12494 3088
rect 12438 3032 12494 3068
rect 13082 12552 13138 12608
rect 13082 12144 13138 12200
rect 13174 11892 13230 11928
rect 13174 11872 13176 11892
rect 13176 11872 13228 11892
rect 13228 11872 13230 11892
rect 13174 11736 13230 11792
rect 13082 11600 13138 11656
rect 13450 15816 13506 15872
rect 13634 15428 13690 15464
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 13634 15408 13636 15428
rect 13636 15408 13688 15428
rect 13688 15408 13690 15428
rect 13266 10784 13322 10840
rect 13174 10648 13230 10704
rect 12898 10124 12954 10160
rect 12898 10104 12900 10124
rect 12900 10104 12952 10124
rect 12952 10104 12954 10124
rect 12898 9968 12954 10024
rect 13082 9832 13138 9888
rect 12898 9460 12900 9480
rect 12900 9460 12952 9480
rect 12952 9460 12954 9480
rect 12898 9424 12954 9460
rect 13082 9016 13138 9072
rect 13450 12164 13506 12200
rect 13450 12144 13452 12164
rect 13452 12144 13504 12164
rect 13504 12144 13506 12164
rect 13266 7384 13322 7440
rect 14554 15544 14610 15600
rect 14370 14048 14426 14104
rect 14002 13368 14058 13424
rect 13726 12416 13782 12472
rect 13634 11212 13690 11248
rect 13634 11192 13636 11212
rect 13636 11192 13688 11212
rect 13688 11192 13690 11212
rect 13818 11192 13874 11248
rect 13818 10920 13874 10976
rect 14278 11328 14334 11384
rect 13634 8472 13690 8528
rect 13174 6996 13230 7032
rect 13174 6976 13176 6996
rect 13176 6976 13228 6996
rect 13228 6976 13230 6996
rect 13174 6840 13230 6896
rect 12714 3576 12770 3632
rect 12990 3576 13046 3632
rect 13542 6976 13598 7032
rect 13358 6452 13414 6488
rect 13358 6432 13360 6452
rect 13360 6432 13412 6452
rect 13412 6432 13414 6452
rect 13634 6296 13690 6352
rect 13542 5616 13598 5672
rect 13358 5480 13414 5536
rect 13266 3848 13322 3904
rect 13542 3848 13598 3904
rect 13818 8744 13874 8800
rect 13818 7112 13874 7168
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15474 16360 15530 16416
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 17038 16632 17094 16688
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 23478 27512 23534 27568
rect 23570 26832 23626 26888
rect 23478 20032 23534 20088
rect 23202 19216 23258 19272
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 18050 16904 18106 16960
rect 17130 15852 17132 15872
rect 17132 15852 17184 15872
rect 17184 15852 17186 15872
rect 16026 15272 16082 15328
rect 17130 15816 17186 15852
rect 17314 15444 17316 15464
rect 17316 15444 17368 15464
rect 17368 15444 17370 15464
rect 17314 15408 17370 15444
rect 16394 15156 16450 15192
rect 16394 15136 16396 15156
rect 16396 15136 16448 15156
rect 16448 15136 16450 15156
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15382 12280 15438 12336
rect 15382 12008 15438 12064
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14370 9288 14426 9344
rect 14278 8200 14334 8256
rect 14186 7792 14242 7848
rect 13726 3984 13782 4040
rect 13818 3476 13820 3496
rect 13820 3476 13872 3496
rect 13872 3476 13874 3496
rect 13818 3440 13874 3476
rect 13726 3304 13782 3360
rect 14002 2760 14058 2816
rect 14370 7792 14426 7848
rect 14370 7520 14426 7576
rect 14646 8472 14702 8528
rect 14554 6024 14610 6080
rect 14738 8064 14794 8120
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15382 5752 15438 5808
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15290 4120 15346 4176
rect 15290 3984 15346 4040
rect 14370 2080 14426 2136
rect 15566 11464 15622 11520
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15658 3712 15714 3768
rect 16026 13776 16082 13832
rect 15934 12980 15990 13016
rect 15934 12960 15936 12980
rect 15936 12960 15988 12980
rect 15988 12960 15990 12980
rect 15934 12280 15990 12336
rect 15934 10240 15990 10296
rect 15842 9324 15844 9344
rect 15844 9324 15896 9344
rect 15896 9324 15898 9344
rect 15842 9288 15898 9324
rect 15934 7928 15990 7984
rect 15842 7792 15898 7848
rect 16854 13912 16910 13968
rect 16394 10648 16450 10704
rect 16854 12008 16910 12064
rect 16302 8608 16358 8664
rect 16118 4800 16174 4856
rect 16394 8200 16450 8256
rect 16394 7112 16450 7168
rect 15934 3984 15990 4040
rect 16486 6568 16542 6624
rect 16670 10004 16672 10024
rect 16672 10004 16724 10024
rect 16724 10004 16726 10024
rect 16670 9968 16726 10004
rect 17406 10512 17462 10568
rect 17314 10240 17370 10296
rect 16946 8608 17002 8664
rect 16854 6296 16910 6352
rect 16578 6160 16634 6216
rect 16854 6160 16910 6216
rect 16486 4972 16488 4992
rect 16488 4972 16540 4992
rect 16540 4972 16542 4992
rect 16486 4936 16542 4972
rect 17130 3984 17186 4040
rect 17314 3984 17370 4040
rect 16302 3304 16358 3360
rect 14738 2624 14794 2680
rect 15014 2624 15070 2680
rect 15566 2760 15622 2816
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 14738 1944 14794 2000
rect 14554 1264 14610 1320
rect 16854 2644 16910 2680
rect 16854 2624 16856 2644
rect 16856 2624 16908 2644
rect 16908 2624 16910 2644
rect 16578 1536 16634 1592
rect 17774 15000 17830 15056
rect 17774 11192 17830 11248
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 20074 16496 20130 16552
rect 18234 16124 18236 16144
rect 18236 16124 18288 16144
rect 18288 16124 18290 16144
rect 18234 16088 18290 16124
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19430 15544 19486 15600
rect 18050 11600 18106 11656
rect 23478 17040 23534 17096
rect 20074 15408 20130 15464
rect 18602 14456 18658 14512
rect 18602 14320 18658 14376
rect 18602 13776 18658 13832
rect 18418 13676 18420 13696
rect 18420 13676 18472 13696
rect 18472 13676 18474 13696
rect 18418 13640 18474 13676
rect 18510 12824 18566 12880
rect 18602 12552 18658 12608
rect 18786 12960 18842 13016
rect 18970 13268 18972 13288
rect 18972 13268 19024 13288
rect 19024 13268 19026 13288
rect 18970 13232 19026 13268
rect 18970 12280 19026 12336
rect 18694 7384 18750 7440
rect 18234 3884 18236 3904
rect 18236 3884 18288 3904
rect 18288 3884 18290 3904
rect 18234 3848 18290 3884
rect 18142 3460 18198 3496
rect 18142 3440 18144 3460
rect 18144 3440 18196 3460
rect 18196 3440 18198 3460
rect 17774 2896 17830 2952
rect 18970 7656 19026 7712
rect 18970 7384 19026 7440
rect 18970 6976 19026 7032
rect 18878 6704 18934 6760
rect 18786 5072 18842 5128
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19430 13504 19486 13560
rect 19338 11736 19394 11792
rect 19338 11600 19394 11656
rect 19614 13132 19616 13152
rect 19616 13132 19668 13152
rect 19668 13132 19670 13152
rect 19614 13096 19670 13132
rect 19798 13096 19854 13152
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19522 12180 19524 12200
rect 19524 12180 19576 12200
rect 19576 12180 19578 12200
rect 19522 12144 19578 12180
rect 20074 12008 20130 12064
rect 20166 11736 20222 11792
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19338 10376 19394 10432
rect 19246 8472 19302 8528
rect 19430 8336 19486 8392
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19982 9988 20038 10024
rect 19982 9968 19984 9988
rect 19984 9968 20036 9988
rect 20036 9968 20038 9988
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19890 7268 19946 7304
rect 19890 7248 19892 7268
rect 19892 7248 19944 7268
rect 19944 7248 19946 7268
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19430 5616 19486 5672
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 18786 4256 18842 4312
rect 18418 3032 18474 3088
rect 17682 2488 17738 2544
rect 17314 1944 17370 2000
rect 17314 1400 17370 1456
rect 18326 1672 18382 1728
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20350 13776 20406 13832
rect 20350 13640 20406 13696
rect 20350 12280 20406 12336
rect 20350 11192 20406 11248
rect 20810 14048 20866 14104
rect 20718 13232 20774 13288
rect 20166 5072 20222 5128
rect 20258 4528 20314 4584
rect 19890 2896 19946 2952
rect 20626 8880 20682 8936
rect 20626 8372 20628 8392
rect 20628 8372 20680 8392
rect 20680 8372 20682 8392
rect 20626 8336 20682 8372
rect 20718 7656 20774 7712
rect 20442 5208 20498 5264
rect 20902 12980 20958 13016
rect 20902 12960 20904 12980
rect 20904 12960 20956 12980
rect 20956 12960 20958 12980
rect 21086 11464 21142 11520
rect 21362 9172 21418 9208
rect 21362 9152 21364 9172
rect 21364 9152 21416 9172
rect 21416 9152 21418 9172
rect 20902 8200 20958 8256
rect 21178 7656 21234 7712
rect 21362 5752 21418 5808
rect 21822 13096 21878 13152
rect 21730 12960 21786 13016
rect 21822 11736 21878 11792
rect 21546 7248 21602 7304
rect 20718 4256 20774 4312
rect 20626 3576 20682 3632
rect 20534 3304 20590 3360
rect 20350 2760 20406 2816
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20074 1808 20130 1864
rect 20718 3168 20774 3224
rect 21178 3884 21180 3904
rect 21180 3884 21232 3904
rect 21232 3884 21234 3904
rect 21178 3848 21234 3884
rect 21454 3712 21510 3768
rect 21362 3576 21418 3632
rect 21454 3476 21456 3496
rect 21456 3476 21508 3496
rect 21508 3476 21510 3496
rect 21454 3440 21510 3476
rect 21730 11192 21786 11248
rect 21914 11056 21970 11112
rect 21730 8508 21732 8528
rect 21732 8508 21784 8528
rect 21784 8508 21786 8528
rect 21730 8472 21786 8508
rect 21914 9016 21970 9072
rect 22006 7112 22062 7168
rect 22006 6568 22062 6624
rect 21822 3304 21878 3360
rect 21822 3032 21878 3088
rect 22374 13776 22430 13832
rect 22282 12960 22338 13016
rect 22834 14864 22890 14920
rect 22558 14068 22614 14104
rect 22558 14048 22560 14068
rect 22560 14048 22612 14068
rect 22612 14048 22614 14068
rect 22558 12824 22614 12880
rect 22466 9560 22522 9616
rect 24030 26152 24086 26208
rect 23846 21428 23848 21448
rect 23848 21428 23900 21448
rect 23900 21428 23902 21448
rect 23846 21392 23902 21428
rect 23478 12688 23534 12744
rect 23478 11192 23534 11248
rect 23018 8336 23074 8392
rect 22650 4120 22706 4176
rect 23478 7384 23534 7440
rect 23478 7268 23534 7304
rect 23478 7248 23480 7268
rect 23480 7248 23532 7268
rect 23532 7248 23534 7268
rect 22650 3440 22706 3496
rect 22374 3304 22430 3360
rect 23478 5072 23534 5128
rect 23938 16496 23994 16552
rect 23846 15988 23848 16008
rect 23848 15988 23900 16008
rect 23900 15988 23902 16008
rect 23846 15952 23902 15988
rect 23754 13776 23810 13832
rect 23662 13640 23718 13696
rect 23846 13096 23902 13152
rect 25226 25472 25282 25528
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24766 24792 24822 24848
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24766 23160 24822 23216
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24674 22480 24730 22536
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24674 21392 24730 21448
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24122 19896 24178 19952
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24214 18672 24270 18728
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24766 19352 24822 19408
rect 24674 18128 24730 18184
rect 24766 17720 24822 17776
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24674 17040 24730 17096
rect 24214 16632 24270 16688
rect 24122 16360 24178 16416
rect 24122 15136 24178 15192
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24766 15952 24822 16008
rect 24674 15272 24730 15328
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24582 13912 24638 13968
rect 24766 13948 24768 13968
rect 24768 13948 24820 13968
rect 24820 13948 24822 13968
rect 24766 13912 24822 13948
rect 24122 13368 24178 13424
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 23754 9424 23810 9480
rect 23662 8336 23718 8392
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24582 11092 24584 11112
rect 24584 11092 24636 11112
rect 24636 11092 24638 11112
rect 24582 11056 24638 11092
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24674 10648 24730 10704
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24122 9152 24178 9208
rect 24030 8472 24086 8528
rect 23662 6840 23718 6896
rect 23662 5752 23718 5808
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24950 12552 25006 12608
rect 25042 12280 25098 12336
rect 25502 24112 25558 24168
rect 25410 22072 25466 22128
rect 25318 18128 25374 18184
rect 25226 10104 25282 10160
rect 24766 7792 24822 7848
rect 24122 7656 24178 7712
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24214 6160 24270 6216
rect 24030 5344 24086 5400
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 25226 9968 25282 10024
rect 25594 20712 25650 20768
rect 25410 7928 25466 7984
rect 25226 7384 25282 7440
rect 24950 4936 25006 4992
rect 23754 4256 23810 4312
rect 23662 3848 23718 3904
rect 22650 2760 22706 2816
rect 23018 2624 23074 2680
rect 23478 2080 23534 2136
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 25318 4120 25374 4176
rect 24122 3848 24178 3904
rect 23938 3712 23994 3768
rect 24030 3188 24086 3224
rect 24030 3168 24032 3188
rect 24032 3168 24084 3188
rect 24084 3168 24086 3188
rect 24030 3032 24086 3088
rect 23938 2216 23994 2272
rect 23662 992 23718 1048
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24582 2896 24638 2952
rect 24490 2388 24492 2408
rect 24492 2388 24544 2408
rect 24544 2388 24546 2408
rect 24490 2352 24546 2388
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 26054 3576 26110 3632
rect 25870 3440 25926 3496
rect 26514 2760 26570 2816
rect 27618 3984 27674 4040
rect 18786 312 18842 368
<< metal3 >>
rect 0 27570 480 27600
rect 2773 27570 2839 27573
rect 0 27568 2839 27570
rect 0 27512 2778 27568
rect 2834 27512 2839 27568
rect 0 27510 2839 27512
rect 0 27480 480 27510
rect 2773 27507 2839 27510
rect 23473 27570 23539 27573
rect 27520 27570 28000 27600
rect 23473 27568 28000 27570
rect 23473 27512 23478 27568
rect 23534 27512 28000 27568
rect 23473 27510 28000 27512
rect 23473 27507 23539 27510
rect 27520 27480 28000 27510
rect 0 26890 480 26920
rect 3049 26890 3115 26893
rect 0 26888 3115 26890
rect 0 26832 3054 26888
rect 3110 26832 3115 26888
rect 0 26830 3115 26832
rect 0 26800 480 26830
rect 3049 26827 3115 26830
rect 23565 26890 23631 26893
rect 27520 26890 28000 26920
rect 23565 26888 28000 26890
rect 23565 26832 23570 26888
rect 23626 26832 28000 26888
rect 23565 26830 28000 26832
rect 23565 26827 23631 26830
rect 27520 26800 28000 26830
rect 0 26210 480 26240
rect 1945 26210 2011 26213
rect 0 26208 2011 26210
rect 0 26152 1950 26208
rect 2006 26152 2011 26208
rect 0 26150 2011 26152
rect 0 26120 480 26150
rect 1945 26147 2011 26150
rect 24025 26210 24091 26213
rect 27520 26210 28000 26240
rect 24025 26208 28000 26210
rect 24025 26152 24030 26208
rect 24086 26152 28000 26208
rect 24025 26150 28000 26152
rect 24025 26147 24091 26150
rect 27520 26120 28000 26150
rect 10277 25600 10597 25601
rect 0 25530 480 25560
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 2865 25530 2931 25533
rect 0 25528 2931 25530
rect 0 25472 2870 25528
rect 2926 25472 2931 25528
rect 0 25470 2931 25472
rect 0 25440 480 25470
rect 2865 25467 2931 25470
rect 25221 25530 25287 25533
rect 27520 25530 28000 25560
rect 25221 25528 28000 25530
rect 25221 25472 25226 25528
rect 25282 25472 28000 25528
rect 25221 25470 28000 25472
rect 25221 25467 25287 25470
rect 27520 25440 28000 25470
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24850 480 24880
rect 1577 24850 1643 24853
rect 0 24848 1643 24850
rect 0 24792 1582 24848
rect 1638 24792 1643 24848
rect 0 24790 1643 24792
rect 0 24760 480 24790
rect 1577 24787 1643 24790
rect 24761 24850 24827 24853
rect 27520 24850 28000 24880
rect 24761 24848 28000 24850
rect 24761 24792 24766 24848
rect 24822 24792 28000 24848
rect 24761 24790 28000 24792
rect 24761 24787 24827 24790
rect 27520 24760 28000 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 0 24170 480 24200
rect 2221 24170 2287 24173
rect 0 24168 2287 24170
rect 0 24112 2226 24168
rect 2282 24112 2287 24168
rect 0 24110 2287 24112
rect 0 24080 480 24110
rect 2221 24107 2287 24110
rect 25497 24170 25563 24173
rect 27520 24170 28000 24200
rect 25497 24168 28000 24170
rect 25497 24112 25502 24168
rect 25558 24112 28000 24168
rect 25497 24110 28000 24112
rect 25497 24107 25563 24110
rect 27520 24080 28000 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 0 23490 480 23520
rect 2037 23490 2103 23493
rect 27520 23490 28000 23520
rect 0 23488 2103 23490
rect 0 23432 2042 23488
rect 2098 23432 2103 23488
rect 0 23430 2103 23432
rect 0 23400 480 23430
rect 2037 23427 2103 23430
rect 24902 23430 28000 23490
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 24761 23218 24827 23221
rect 24902 23218 24962 23430
rect 27520 23400 28000 23430
rect 24761 23216 24962 23218
rect 24761 23160 24766 23216
rect 24822 23160 24962 23216
rect 24761 23158 24962 23160
rect 24761 23155 24827 23158
rect 5610 22880 5930 22881
rect 0 22810 480 22840
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 2957 22810 3023 22813
rect 27520 22810 28000 22840
rect 0 22808 3023 22810
rect 0 22752 2962 22808
rect 3018 22752 3023 22808
rect 0 22750 3023 22752
rect 0 22720 480 22750
rect 2957 22747 3023 22750
rect 24718 22750 28000 22810
rect 24718 22541 24778 22750
rect 27520 22720 28000 22750
rect 24669 22536 24778 22541
rect 24669 22480 24674 22536
rect 24730 22480 24778 22536
rect 24669 22478 24778 22480
rect 24669 22475 24735 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 0 22130 480 22160
rect 1577 22130 1643 22133
rect 0 22128 1643 22130
rect 0 22072 1582 22128
rect 1638 22072 1643 22128
rect 0 22070 1643 22072
rect 0 22040 480 22070
rect 1577 22067 1643 22070
rect 25405 22130 25471 22133
rect 27520 22130 28000 22160
rect 25405 22128 28000 22130
rect 25405 22072 25410 22128
rect 25466 22072 28000 22128
rect 25405 22070 28000 22072
rect 25405 22067 25471 22070
rect 27520 22040 28000 22070
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 0 21450 480 21480
rect 1485 21450 1551 21453
rect 0 21448 1551 21450
rect 0 21392 1490 21448
rect 1546 21392 1551 21448
rect 0 21390 1551 21392
rect 0 21360 480 21390
rect 1485 21387 1551 21390
rect 10869 21450 10935 21453
rect 23841 21450 23907 21453
rect 10869 21448 23907 21450
rect 10869 21392 10874 21448
rect 10930 21392 23846 21448
rect 23902 21392 23907 21448
rect 10869 21390 23907 21392
rect 10869 21387 10935 21390
rect 23841 21387 23907 21390
rect 24669 21450 24735 21453
rect 27520 21450 28000 21480
rect 24669 21448 28000 21450
rect 24669 21392 24674 21448
rect 24730 21392 28000 21448
rect 24669 21390 28000 21392
rect 24669 21387 24735 21390
rect 27520 21360 28000 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 0 20770 480 20800
rect 1393 20770 1459 20773
rect 0 20768 1459 20770
rect 0 20712 1398 20768
rect 1454 20712 1459 20768
rect 0 20710 1459 20712
rect 0 20680 480 20710
rect 1393 20707 1459 20710
rect 1853 20770 1919 20773
rect 2037 20770 2103 20773
rect 1853 20768 2103 20770
rect 1853 20712 1858 20768
rect 1914 20712 2042 20768
rect 2098 20712 2103 20768
rect 1853 20710 2103 20712
rect 1853 20707 1919 20710
rect 2037 20707 2103 20710
rect 25589 20770 25655 20773
rect 27520 20770 28000 20800
rect 25589 20768 28000 20770
rect 25589 20712 25594 20768
rect 25650 20712 28000 20768
rect 25589 20710 28000 20712
rect 25589 20707 25655 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 27520 20680 28000 20710
rect 24277 20639 24597 20640
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 1577 20090 1643 20093
rect 0 20088 1643 20090
rect 0 20032 1582 20088
rect 1638 20032 1643 20088
rect 0 20030 1643 20032
rect 0 20000 480 20030
rect 1577 20027 1643 20030
rect 23473 20090 23539 20093
rect 27520 20090 28000 20120
rect 23473 20088 28000 20090
rect 23473 20032 23478 20088
rect 23534 20032 28000 20088
rect 23473 20030 28000 20032
rect 23473 20027 23539 20030
rect 27520 20000 28000 20030
rect 21398 19892 21404 19956
rect 21468 19954 21474 19956
rect 24117 19954 24183 19957
rect 21468 19952 24183 19954
rect 21468 19896 24122 19952
rect 24178 19896 24183 19952
rect 21468 19894 24183 19896
rect 21468 19892 21474 19894
rect 24117 19891 24183 19894
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 0 19410 480 19440
rect 1669 19410 1735 19413
rect 0 19408 1735 19410
rect 0 19352 1674 19408
rect 1730 19352 1735 19408
rect 0 19350 1735 19352
rect 0 19320 480 19350
rect 1669 19347 1735 19350
rect 24761 19410 24827 19413
rect 27520 19410 28000 19440
rect 24761 19408 28000 19410
rect 24761 19352 24766 19408
rect 24822 19352 28000 19408
rect 24761 19350 28000 19352
rect 24761 19347 24827 19350
rect 27520 19320 28000 19350
rect 2405 19274 2471 19277
rect 11697 19274 11763 19277
rect 2405 19272 11763 19274
rect 2405 19216 2410 19272
rect 2466 19216 11702 19272
rect 11758 19216 11763 19272
rect 2405 19214 11763 19216
rect 2405 19211 2471 19214
rect 11697 19211 11763 19214
rect 14917 19274 14983 19277
rect 23197 19274 23263 19277
rect 14917 19272 23263 19274
rect 14917 19216 14922 19272
rect 14978 19216 23202 19272
rect 23258 19216 23263 19272
rect 14917 19214 23263 19216
rect 14917 19211 14983 19214
rect 23197 19211 23263 19214
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 2405 18866 2471 18869
rect 9673 18866 9739 18869
rect 2405 18864 9739 18866
rect 2405 18808 2410 18864
rect 2466 18808 9678 18864
rect 9734 18808 9739 18864
rect 2405 18806 9739 18808
rect 2405 18803 2471 18806
rect 9673 18803 9739 18806
rect 0 18730 480 18760
rect 1485 18730 1551 18733
rect 0 18728 1551 18730
rect 0 18672 1490 18728
rect 1546 18672 1551 18728
rect 0 18670 1551 18672
rect 0 18640 480 18670
rect 1485 18667 1551 18670
rect 2497 18730 2563 18733
rect 12433 18730 12499 18733
rect 2497 18728 12499 18730
rect 2497 18672 2502 18728
rect 2558 18672 12438 18728
rect 12494 18672 12499 18728
rect 2497 18670 12499 18672
rect 2497 18667 2563 18670
rect 12433 18667 12499 18670
rect 24209 18730 24275 18733
rect 27520 18730 28000 18760
rect 24209 18728 28000 18730
rect 24209 18672 24214 18728
rect 24270 18672 28000 18728
rect 24209 18670 28000 18672
rect 24209 18667 24275 18670
rect 27520 18640 28000 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 24669 18186 24735 18189
rect 25313 18186 25379 18189
rect 24669 18184 25379 18186
rect 24669 18128 24674 18184
rect 24730 18128 25318 18184
rect 25374 18128 25379 18184
rect 24669 18126 25379 18128
rect 24669 18123 24735 18126
rect 25313 18123 25379 18126
rect 0 18050 480 18080
rect 1577 18050 1643 18053
rect 0 18048 1643 18050
rect 0 17992 1582 18048
rect 1638 17992 1643 18048
rect 0 17990 1643 17992
rect 0 17960 480 17990
rect 1577 17987 1643 17990
rect 2037 18050 2103 18053
rect 9121 18050 9187 18053
rect 27520 18050 28000 18080
rect 2037 18048 9187 18050
rect 2037 17992 2042 18048
rect 2098 17992 9126 18048
rect 9182 17992 9187 18048
rect 2037 17990 9187 17992
rect 2037 17987 2103 17990
rect 9121 17987 9187 17990
rect 24902 17990 28000 18050
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 24761 17778 24827 17781
rect 24902 17778 24962 17990
rect 27520 17960 28000 17990
rect 24761 17776 24962 17778
rect 24761 17720 24766 17776
rect 24822 17720 24962 17776
rect 24761 17718 24962 17720
rect 24761 17715 24827 17718
rect 5610 17440 5930 17441
rect 0 17370 480 17400
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 1393 17370 1459 17373
rect 27520 17370 28000 17400
rect 0 17368 1459 17370
rect 0 17312 1398 17368
rect 1454 17312 1459 17368
rect 0 17310 1459 17312
rect 0 17280 480 17310
rect 1393 17307 1459 17310
rect 24672 17310 28000 17370
rect 2129 17234 2195 17237
rect 13261 17234 13327 17237
rect 2129 17232 13327 17234
rect 2129 17176 2134 17232
rect 2190 17176 13266 17232
rect 13322 17176 13327 17232
rect 2129 17174 13327 17176
rect 2129 17171 2195 17174
rect 13261 17171 13327 17174
rect 24672 17101 24732 17310
rect 27520 17280 28000 17310
rect 10685 17098 10751 17101
rect 23473 17098 23539 17101
rect 10685 17096 23539 17098
rect 10685 17040 10690 17096
rect 10746 17040 23478 17096
rect 23534 17040 23539 17096
rect 10685 17038 23539 17040
rect 10685 17035 10751 17038
rect 23473 17035 23539 17038
rect 24669 17096 24735 17101
rect 24669 17040 24674 17096
rect 24730 17040 24735 17096
rect 24669 17035 24735 17040
rect 8017 16962 8083 16965
rect 10133 16962 10199 16965
rect 8017 16960 10199 16962
rect 8017 16904 8022 16960
rect 8078 16904 10138 16960
rect 10194 16904 10199 16960
rect 8017 16902 10199 16904
rect 8017 16899 8083 16902
rect 10133 16899 10199 16902
rect 11053 16962 11119 16965
rect 18045 16962 18111 16965
rect 11053 16960 18111 16962
rect 11053 16904 11058 16960
rect 11114 16904 18050 16960
rect 18106 16904 18111 16960
rect 11053 16902 18111 16904
rect 11053 16899 11119 16902
rect 18045 16899 18111 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 0 16690 480 16720
rect 1945 16690 2011 16693
rect 0 16688 2011 16690
rect 0 16632 1950 16688
rect 2006 16632 2011 16688
rect 0 16630 2011 16632
rect 0 16600 480 16630
rect 1945 16627 2011 16630
rect 12709 16690 12775 16693
rect 17033 16690 17099 16693
rect 12709 16688 17099 16690
rect 12709 16632 12714 16688
rect 12770 16632 17038 16688
rect 17094 16632 17099 16688
rect 12709 16630 17099 16632
rect 12709 16627 12775 16630
rect 17033 16627 17099 16630
rect 24209 16690 24275 16693
rect 27520 16690 28000 16720
rect 24209 16688 28000 16690
rect 24209 16632 24214 16688
rect 24270 16632 28000 16688
rect 24209 16630 28000 16632
rect 24209 16627 24275 16630
rect 27520 16600 28000 16630
rect 20069 16554 20135 16557
rect 23933 16554 23999 16557
rect 20069 16552 23999 16554
rect 20069 16496 20074 16552
rect 20130 16496 23938 16552
rect 23994 16496 23999 16552
rect 20069 16494 23999 16496
rect 20069 16491 20135 16494
rect 23933 16491 23999 16494
rect 15469 16418 15535 16421
rect 24117 16418 24183 16421
rect 15469 16416 24183 16418
rect 15469 16360 15474 16416
rect 15530 16360 24122 16416
rect 24178 16360 24183 16416
rect 15469 16358 24183 16360
rect 15469 16355 15535 16358
rect 24117 16355 24183 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 10133 16146 10199 16149
rect 18229 16146 18295 16149
rect 10133 16144 18295 16146
rect 10133 16088 10138 16144
rect 10194 16088 18234 16144
rect 18290 16088 18295 16144
rect 10133 16086 18295 16088
rect 10133 16083 10199 16086
rect 18229 16083 18295 16086
rect 0 16010 480 16040
rect 1577 16010 1643 16013
rect 0 16008 1643 16010
rect 0 15952 1582 16008
rect 1638 15952 1643 16008
rect 0 15950 1643 15952
rect 0 15920 480 15950
rect 1577 15947 1643 15950
rect 7649 16010 7715 16013
rect 23841 16010 23907 16013
rect 7649 16008 23907 16010
rect 7649 15952 7654 16008
rect 7710 15952 23846 16008
rect 23902 15952 23907 16008
rect 7649 15950 23907 15952
rect 7649 15947 7715 15950
rect 23841 15947 23907 15950
rect 24761 16010 24827 16013
rect 27520 16010 28000 16040
rect 24761 16008 28000 16010
rect 24761 15952 24766 16008
rect 24822 15952 28000 16008
rect 24761 15950 28000 15952
rect 24761 15947 24827 15950
rect 27520 15920 28000 15950
rect 13445 15874 13511 15877
rect 17125 15874 17191 15877
rect 13445 15872 17191 15874
rect 13445 15816 13450 15872
rect 13506 15816 17130 15872
rect 17186 15816 17191 15872
rect 13445 15814 17191 15816
rect 13445 15811 13511 15814
rect 17125 15811 17191 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 7833 15602 7899 15605
rect 12157 15602 12223 15605
rect 7833 15600 12223 15602
rect 7833 15544 7838 15600
rect 7894 15544 12162 15600
rect 12218 15544 12223 15600
rect 7833 15542 12223 15544
rect 7833 15539 7899 15542
rect 12157 15539 12223 15542
rect 14549 15602 14615 15605
rect 19425 15602 19491 15605
rect 14549 15600 19491 15602
rect 14549 15544 14554 15600
rect 14610 15544 19430 15600
rect 19486 15544 19491 15600
rect 14549 15542 19491 15544
rect 14549 15539 14615 15542
rect 19425 15539 19491 15542
rect 2405 15466 2471 15469
rect 4889 15466 4955 15469
rect 2405 15464 4955 15466
rect 2405 15408 2410 15464
rect 2466 15408 4894 15464
rect 4950 15408 4955 15464
rect 2405 15406 4955 15408
rect 2405 15403 2471 15406
rect 4889 15403 4955 15406
rect 13629 15466 13695 15469
rect 17309 15466 17375 15469
rect 20069 15466 20135 15469
rect 13629 15464 17375 15466
rect 13629 15408 13634 15464
rect 13690 15408 17314 15464
rect 17370 15408 17375 15464
rect 13629 15406 17375 15408
rect 13629 15403 13695 15406
rect 17309 15403 17375 15406
rect 17542 15464 20135 15466
rect 17542 15408 20074 15464
rect 20130 15408 20135 15464
rect 17542 15406 20135 15408
rect 0 15330 480 15360
rect 1669 15330 1735 15333
rect 0 15328 1735 15330
rect 0 15272 1674 15328
rect 1730 15272 1735 15328
rect 0 15270 1735 15272
rect 0 15240 480 15270
rect 1669 15267 1735 15270
rect 16021 15330 16087 15333
rect 17542 15330 17602 15406
rect 20069 15403 20135 15406
rect 16021 15328 17602 15330
rect 16021 15272 16026 15328
rect 16082 15272 17602 15328
rect 16021 15270 17602 15272
rect 24669 15330 24735 15333
rect 27520 15330 28000 15360
rect 24669 15328 28000 15330
rect 24669 15272 24674 15328
rect 24730 15272 28000 15328
rect 24669 15270 28000 15272
rect 16021 15267 16087 15270
rect 24669 15267 24735 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 27520 15240 28000 15270
rect 24277 15199 24597 15200
rect 16389 15194 16455 15197
rect 24117 15194 24183 15197
rect 16389 15192 24183 15194
rect 16389 15136 16394 15192
rect 16450 15136 24122 15192
rect 24178 15136 24183 15192
rect 16389 15134 24183 15136
rect 16389 15131 16455 15134
rect 24117 15131 24183 15134
rect 8293 15058 8359 15061
rect 10961 15058 11027 15061
rect 8293 15056 11027 15058
rect 8293 15000 8298 15056
rect 8354 15000 10966 15056
rect 11022 15000 11027 15056
rect 8293 14998 11027 15000
rect 8293 14995 8359 14998
rect 10961 14995 11027 14998
rect 17769 15058 17835 15061
rect 21398 15058 21404 15060
rect 17769 15056 21404 15058
rect 17769 15000 17774 15056
rect 17830 15000 21404 15056
rect 17769 14998 21404 15000
rect 17769 14995 17835 14998
rect 21398 14996 21404 14998
rect 21468 14996 21474 15060
rect 2037 14922 2103 14925
rect 12341 14922 12407 14925
rect 22829 14922 22895 14925
rect 2037 14920 22895 14922
rect 2037 14864 2042 14920
rect 2098 14864 12346 14920
rect 12402 14864 22834 14920
rect 22890 14864 22895 14920
rect 2037 14862 22895 14864
rect 2037 14859 2103 14862
rect 12341 14859 12407 14862
rect 22829 14859 22895 14862
rect 10277 14720 10597 14721
rect 0 14650 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 1485 14650 1551 14653
rect 27520 14650 28000 14680
rect 0 14648 1551 14650
rect 0 14592 1490 14648
rect 1546 14592 1551 14648
rect 0 14590 1551 14592
rect 0 14560 480 14590
rect 1485 14587 1551 14590
rect 27478 14560 28000 14650
rect 18597 14514 18663 14517
rect 27478 14514 27538 14560
rect 18597 14512 27538 14514
rect 18597 14456 18602 14512
rect 18658 14456 27538 14512
rect 18597 14454 27538 14456
rect 18597 14451 18663 14454
rect 10961 14378 11027 14381
rect 18597 14378 18663 14381
rect 10961 14376 18663 14378
rect 10961 14320 10966 14376
rect 11022 14320 18602 14376
rect 18658 14320 18663 14376
rect 10961 14318 18663 14320
rect 10961 14315 11027 14318
rect 18597 14315 18663 14318
rect 6913 14242 6979 14245
rect 12893 14242 12959 14245
rect 6913 14240 12959 14242
rect 6913 14184 6918 14240
rect 6974 14184 12898 14240
rect 12954 14184 12959 14240
rect 6913 14182 12959 14184
rect 6913 14179 6979 14182
rect 12893 14179 12959 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 10041 14106 10107 14109
rect 14365 14106 14431 14109
rect 10041 14104 14431 14106
rect 10041 14048 10046 14104
rect 10102 14048 14370 14104
rect 14426 14048 14431 14104
rect 10041 14046 14431 14048
rect 10041 14043 10107 14046
rect 14365 14043 14431 14046
rect 20805 14106 20871 14109
rect 22553 14106 22619 14109
rect 20805 14104 22619 14106
rect 20805 14048 20810 14104
rect 20866 14048 22558 14104
rect 22614 14048 22619 14104
rect 20805 14046 22619 14048
rect 20805 14043 20871 14046
rect 22553 14043 22619 14046
rect 0 13970 480 14000
rect 1577 13970 1643 13973
rect 0 13968 1643 13970
rect 0 13912 1582 13968
rect 1638 13912 1643 13968
rect 0 13910 1643 13912
rect 0 13880 480 13910
rect 1577 13907 1643 13910
rect 4705 13970 4771 13973
rect 10961 13970 11027 13973
rect 12433 13970 12499 13973
rect 4705 13968 9506 13970
rect 4705 13912 4710 13968
rect 4766 13912 9506 13968
rect 4705 13910 9506 13912
rect 4705 13907 4771 13910
rect 2037 13834 2103 13837
rect 9305 13834 9371 13837
rect 2037 13832 9371 13834
rect 2037 13776 2042 13832
rect 2098 13776 9310 13832
rect 9366 13776 9371 13832
rect 2037 13774 9371 13776
rect 9446 13834 9506 13910
rect 10961 13968 12499 13970
rect 10961 13912 10966 13968
rect 11022 13912 12438 13968
rect 12494 13912 12499 13968
rect 10961 13910 12499 13912
rect 10961 13907 11027 13910
rect 12433 13907 12499 13910
rect 16849 13970 16915 13973
rect 24577 13970 24643 13973
rect 16849 13968 24643 13970
rect 16849 13912 16854 13968
rect 16910 13912 24582 13968
rect 24638 13912 24643 13968
rect 16849 13910 24643 13912
rect 16849 13907 16915 13910
rect 24577 13907 24643 13910
rect 24761 13970 24827 13973
rect 27520 13970 28000 14000
rect 24761 13968 28000 13970
rect 24761 13912 24766 13968
rect 24822 13912 28000 13968
rect 24761 13910 28000 13912
rect 24761 13907 24827 13910
rect 27520 13880 28000 13910
rect 16021 13834 16087 13837
rect 9446 13832 16087 13834
rect 9446 13776 16026 13832
rect 16082 13776 16087 13832
rect 9446 13774 16087 13776
rect 2037 13771 2103 13774
rect 9305 13771 9371 13774
rect 16021 13771 16087 13774
rect 18597 13834 18663 13837
rect 20345 13834 20411 13837
rect 18597 13832 20411 13834
rect 18597 13776 18602 13832
rect 18658 13776 20350 13832
rect 20406 13776 20411 13832
rect 18597 13774 20411 13776
rect 18597 13771 18663 13774
rect 20345 13771 20411 13774
rect 22369 13834 22435 13837
rect 23749 13834 23815 13837
rect 22369 13832 23815 13834
rect 22369 13776 22374 13832
rect 22430 13776 23754 13832
rect 23810 13776 23815 13832
rect 22369 13774 23815 13776
rect 22369 13771 22435 13774
rect 23749 13771 23815 13774
rect 11421 13698 11487 13701
rect 18413 13698 18479 13701
rect 11421 13696 18479 13698
rect 11421 13640 11426 13696
rect 11482 13640 18418 13696
rect 18474 13640 18479 13696
rect 11421 13638 18479 13640
rect 11421 13635 11487 13638
rect 18413 13635 18479 13638
rect 20345 13698 20411 13701
rect 23657 13698 23723 13701
rect 20345 13696 23723 13698
rect 20345 13640 20350 13696
rect 20406 13640 23662 13696
rect 23718 13640 23723 13696
rect 20345 13638 23723 13640
rect 20345 13635 20411 13638
rect 23657 13635 23723 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 10685 13562 10751 13565
rect 19425 13562 19491 13565
rect 10685 13560 19491 13562
rect 10685 13504 10690 13560
rect 10746 13504 19430 13560
rect 19486 13504 19491 13560
rect 10685 13502 19491 13504
rect 10685 13499 10751 13502
rect 19425 13499 19491 13502
rect 5993 13426 6059 13429
rect 2684 13424 6059 13426
rect 2684 13368 5998 13424
rect 6054 13368 6059 13424
rect 2684 13366 6059 13368
rect 0 13290 480 13320
rect 2684 13290 2744 13366
rect 5993 13363 6059 13366
rect 7281 13426 7347 13429
rect 9489 13426 9555 13429
rect 10225 13426 10291 13429
rect 7281 13424 10291 13426
rect 7281 13368 7286 13424
rect 7342 13368 9494 13424
rect 9550 13368 10230 13424
rect 10286 13368 10291 13424
rect 7281 13366 10291 13368
rect 7281 13363 7347 13366
rect 9489 13363 9555 13366
rect 10225 13363 10291 13366
rect 13997 13426 14063 13429
rect 24117 13426 24183 13429
rect 13997 13424 24183 13426
rect 13997 13368 14002 13424
rect 14058 13368 24122 13424
rect 24178 13368 24183 13424
rect 13997 13366 24183 13368
rect 13997 13363 14063 13366
rect 24117 13363 24183 13366
rect 0 13230 2744 13290
rect 4797 13290 4863 13293
rect 11329 13290 11395 13293
rect 4797 13288 11395 13290
rect 4797 13232 4802 13288
rect 4858 13232 11334 13288
rect 11390 13232 11395 13288
rect 4797 13230 11395 13232
rect 0 13200 480 13230
rect 4797 13227 4863 13230
rect 11329 13227 11395 13230
rect 18965 13290 19031 13293
rect 20713 13290 20779 13293
rect 27520 13290 28000 13320
rect 18965 13288 20779 13290
rect 18965 13232 18970 13288
rect 19026 13232 20718 13288
rect 20774 13232 20779 13288
rect 18965 13230 20779 13232
rect 18965 13227 19031 13230
rect 20713 13227 20779 13230
rect 23982 13230 28000 13290
rect 2865 13154 2931 13157
rect 4705 13154 4771 13157
rect 2865 13152 4771 13154
rect 2865 13096 2870 13152
rect 2926 13096 4710 13152
rect 4766 13096 4771 13152
rect 2865 13094 4771 13096
rect 2865 13091 2931 13094
rect 4705 13091 4771 13094
rect 5993 13154 6059 13157
rect 12341 13154 12407 13157
rect 19609 13154 19675 13157
rect 5993 13152 12407 13154
rect 5993 13096 5998 13152
rect 6054 13096 12346 13152
rect 12402 13096 12407 13152
rect 5993 13094 12407 13096
rect 5993 13091 6059 13094
rect 12341 13091 12407 13094
rect 15702 13152 19675 13154
rect 15702 13096 19614 13152
rect 19670 13096 19675 13152
rect 15702 13094 19675 13096
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 8845 13018 8911 13021
rect 11145 13018 11211 13021
rect 8845 13016 11211 13018
rect 8845 12960 8850 13016
rect 8906 12960 11150 13016
rect 11206 12960 11211 13016
rect 8845 12958 11211 12960
rect 8845 12955 8911 12958
rect 11145 12955 11211 12958
rect 6729 12882 6795 12885
rect 15702 12882 15762 13094
rect 19609 13091 19675 13094
rect 19793 13154 19859 13157
rect 21817 13154 21883 13157
rect 19793 13152 21883 13154
rect 19793 13096 19798 13152
rect 19854 13096 21822 13152
rect 21878 13096 21883 13152
rect 19793 13094 21883 13096
rect 19793 13091 19859 13094
rect 21817 13091 21883 13094
rect 23841 13154 23907 13157
rect 23982 13154 24042 13230
rect 27520 13200 28000 13230
rect 23841 13152 24042 13154
rect 23841 13096 23846 13152
rect 23902 13096 24042 13152
rect 23841 13094 24042 13096
rect 23841 13091 23907 13094
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 15929 13018 15995 13021
rect 18781 13018 18847 13021
rect 20897 13018 20963 13021
rect 15929 13016 20963 13018
rect 15929 12960 15934 13016
rect 15990 12960 18786 13016
rect 18842 12960 20902 13016
rect 20958 12960 20963 13016
rect 15929 12958 20963 12960
rect 15929 12955 15995 12958
rect 18781 12955 18847 12958
rect 20897 12955 20963 12958
rect 21725 13018 21791 13021
rect 22277 13018 22343 13021
rect 21725 13016 22343 13018
rect 21725 12960 21730 13016
rect 21786 12960 22282 13016
rect 22338 12960 22343 13016
rect 21725 12958 22343 12960
rect 21725 12955 21791 12958
rect 22277 12955 22343 12958
rect 6729 12880 15762 12882
rect 6729 12824 6734 12880
rect 6790 12824 15762 12880
rect 6729 12822 15762 12824
rect 18505 12882 18571 12885
rect 22553 12882 22619 12885
rect 18505 12880 22619 12882
rect 18505 12824 18510 12880
rect 18566 12824 22558 12880
rect 22614 12824 22619 12880
rect 18505 12822 22619 12824
rect 6729 12819 6795 12822
rect 18505 12819 18571 12822
rect 22553 12819 22619 12822
rect 2037 12746 2103 12749
rect 4981 12746 5047 12749
rect 23473 12746 23539 12749
rect 2037 12744 23539 12746
rect 2037 12688 2042 12744
rect 2098 12688 4986 12744
rect 5042 12688 23478 12744
rect 23534 12688 23539 12744
rect 2037 12686 23539 12688
rect 2037 12683 2103 12686
rect 4981 12683 5047 12686
rect 0 12610 480 12640
rect 3417 12610 3483 12613
rect 8661 12610 8727 12613
rect 0 12608 3483 12610
rect 0 12552 3422 12608
rect 3478 12552 3483 12608
rect 0 12550 3483 12552
rect 0 12520 480 12550
rect 3417 12547 3483 12550
rect 8342 12608 8727 12610
rect 8342 12552 8666 12608
rect 8722 12552 8727 12608
rect 8342 12550 8727 12552
rect 2221 12474 2287 12477
rect 8342 12474 8402 12550
rect 8661 12547 8727 12550
rect 10961 12610 11027 12613
rect 13077 12610 13143 12613
rect 10961 12608 13143 12610
rect 10961 12552 10966 12608
rect 11022 12552 13082 12608
rect 13138 12552 13143 12608
rect 10961 12550 13143 12552
rect 18462 12610 18522 12686
rect 23473 12683 23539 12686
rect 18597 12610 18663 12613
rect 18462 12608 18663 12610
rect 18462 12552 18602 12608
rect 18658 12552 18663 12608
rect 18462 12550 18663 12552
rect 10961 12547 11027 12550
rect 13077 12547 13143 12550
rect 18597 12547 18663 12550
rect 24945 12610 25011 12613
rect 27520 12610 28000 12640
rect 24945 12608 28000 12610
rect 24945 12552 24950 12608
rect 25006 12552 28000 12608
rect 24945 12550 28000 12552
rect 24945 12547 25011 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 27520 12520 28000 12550
rect 19610 12479 19930 12480
rect 2221 12472 8402 12474
rect 2221 12416 2226 12472
rect 2282 12416 8402 12472
rect 2221 12414 8402 12416
rect 8569 12474 8635 12477
rect 13721 12474 13787 12477
rect 8569 12472 10196 12474
rect 8569 12416 8574 12472
rect 8630 12416 10196 12472
rect 8569 12414 10196 12416
rect 2221 12411 2287 12414
rect 8569 12411 8635 12414
rect 7741 12338 7807 12341
rect 9765 12338 9831 12341
rect 7741 12336 9831 12338
rect 7741 12280 7746 12336
rect 7802 12280 9770 12336
rect 9826 12280 9831 12336
rect 7741 12278 9831 12280
rect 10136 12338 10196 12414
rect 10688 12472 13787 12474
rect 10688 12416 13726 12472
rect 13782 12416 13787 12472
rect 10688 12414 13787 12416
rect 10688 12338 10748 12414
rect 13721 12411 13787 12414
rect 10136 12278 10748 12338
rect 11053 12338 11119 12341
rect 15377 12338 15443 12341
rect 11053 12336 15443 12338
rect 11053 12280 11058 12336
rect 11114 12280 15382 12336
rect 15438 12280 15443 12336
rect 11053 12278 15443 12280
rect 7741 12275 7807 12278
rect 9765 12275 9831 12278
rect 11053 12275 11119 12278
rect 15377 12275 15443 12278
rect 15929 12338 15995 12341
rect 18965 12338 19031 12341
rect 15929 12336 19031 12338
rect 15929 12280 15934 12336
rect 15990 12280 18970 12336
rect 19026 12280 19031 12336
rect 15929 12278 19031 12280
rect 15929 12275 15995 12278
rect 18965 12275 19031 12278
rect 20345 12338 20411 12341
rect 25037 12338 25103 12341
rect 20345 12336 25103 12338
rect 20345 12280 20350 12336
rect 20406 12280 25042 12336
rect 25098 12280 25103 12336
rect 20345 12278 25103 12280
rect 20345 12275 20411 12278
rect 25037 12275 25103 12278
rect 9806 12140 9812 12204
rect 9876 12202 9882 12204
rect 12157 12202 12223 12205
rect 9876 12200 12223 12202
rect 9876 12144 12162 12200
rect 12218 12144 12223 12200
rect 9876 12142 12223 12144
rect 9876 12140 9882 12142
rect 12157 12139 12223 12142
rect 13077 12202 13143 12205
rect 13302 12202 13308 12204
rect 13077 12200 13308 12202
rect 13077 12144 13082 12200
rect 13138 12144 13308 12200
rect 13077 12142 13308 12144
rect 13077 12139 13143 12142
rect 13302 12140 13308 12142
rect 13372 12140 13378 12204
rect 13445 12202 13511 12205
rect 19517 12202 19583 12205
rect 13445 12200 19583 12202
rect 13445 12144 13450 12200
rect 13506 12144 19522 12200
rect 19578 12144 19583 12200
rect 13445 12142 19583 12144
rect 13445 12139 13511 12142
rect 19517 12139 19583 12142
rect 9489 12066 9555 12069
rect 10685 12066 10751 12069
rect 9489 12064 10751 12066
rect 9489 12008 9494 12064
rect 9550 12008 10690 12064
rect 10746 12008 10751 12064
rect 9489 12006 10751 12008
rect 9489 12003 9555 12006
rect 10685 12003 10751 12006
rect 10961 12066 11027 12069
rect 15377 12066 15443 12069
rect 16849 12066 16915 12069
rect 20069 12066 20135 12069
rect 10961 12064 12082 12066
rect 10961 12008 10966 12064
rect 11022 12008 12082 12064
rect 10961 12006 12082 12008
rect 10961 12003 11027 12006
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 9581 11930 9647 11933
rect 11789 11930 11855 11933
rect 0 11870 5044 11930
rect 0 11840 480 11870
rect 4984 11794 5044 11870
rect 9581 11928 11855 11930
rect 9581 11872 9586 11928
rect 9642 11872 11794 11928
rect 11850 11872 11855 11928
rect 9581 11870 11855 11872
rect 12022 11930 12082 12006
rect 15377 12064 20135 12066
rect 15377 12008 15382 12064
rect 15438 12008 16854 12064
rect 16910 12008 20074 12064
rect 20130 12008 20135 12064
rect 15377 12006 20135 12008
rect 15377 12003 15443 12006
rect 16849 12003 16915 12006
rect 20069 12003 20135 12006
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 13169 11930 13235 11933
rect 27520 11930 28000 11960
rect 12022 11928 13235 11930
rect 12022 11872 13174 11928
rect 13230 11872 13235 11928
rect 12022 11870 13235 11872
rect 9581 11867 9647 11870
rect 11789 11867 11855 11870
rect 13169 11867 13235 11870
rect 24902 11870 28000 11930
rect 8385 11794 8451 11797
rect 4984 11792 8451 11794
rect 4984 11736 8390 11792
rect 8446 11736 8451 11792
rect 4984 11734 8451 11736
rect 8385 11731 8451 11734
rect 13169 11794 13235 11797
rect 19333 11794 19399 11797
rect 20161 11794 20227 11797
rect 13169 11792 19399 11794
rect 13169 11736 13174 11792
rect 13230 11736 19338 11792
rect 19394 11736 19399 11792
rect 13169 11734 19399 11736
rect 13169 11731 13235 11734
rect 19333 11731 19399 11734
rect 19566 11792 20227 11794
rect 19566 11736 20166 11792
rect 20222 11736 20227 11792
rect 19566 11734 20227 11736
rect 2681 11658 2747 11661
rect 9254 11658 9260 11660
rect 2681 11656 9260 11658
rect 2681 11600 2686 11656
rect 2742 11600 9260 11656
rect 2681 11598 9260 11600
rect 2681 11595 2747 11598
rect 9254 11596 9260 11598
rect 9324 11596 9330 11660
rect 9489 11658 9555 11661
rect 11973 11658 12039 11661
rect 9489 11656 12039 11658
rect 9489 11600 9494 11656
rect 9550 11600 11978 11656
rect 12034 11600 12039 11656
rect 9489 11598 12039 11600
rect 9489 11595 9555 11598
rect 11973 11595 12039 11598
rect 13077 11658 13143 11661
rect 18045 11658 18111 11661
rect 13077 11656 18111 11658
rect 13077 11600 13082 11656
rect 13138 11600 18050 11656
rect 18106 11600 18111 11656
rect 13077 11598 18111 11600
rect 13077 11595 13143 11598
rect 18045 11595 18111 11598
rect 19333 11658 19399 11661
rect 19566 11658 19626 11734
rect 20161 11731 20227 11734
rect 21817 11794 21883 11797
rect 24902 11794 24962 11870
rect 27520 11840 28000 11870
rect 21817 11792 24962 11794
rect 21817 11736 21822 11792
rect 21878 11736 24962 11792
rect 21817 11734 24962 11736
rect 21817 11731 21883 11734
rect 19333 11656 19626 11658
rect 19333 11600 19338 11656
rect 19394 11600 19626 11656
rect 19333 11598 19626 11600
rect 19333 11595 19399 11598
rect 2589 11522 2655 11525
rect 5533 11522 5599 11525
rect 2589 11520 5599 11522
rect 2589 11464 2594 11520
rect 2650 11464 5538 11520
rect 5594 11464 5599 11520
rect 2589 11462 5599 11464
rect 2589 11459 2655 11462
rect 5533 11459 5599 11462
rect 6177 11522 6243 11525
rect 9213 11522 9279 11525
rect 15561 11522 15627 11525
rect 6177 11520 9279 11522
rect 6177 11464 6182 11520
rect 6238 11464 9218 11520
rect 9274 11464 9279 11520
rect 6177 11462 9279 11464
rect 6177 11459 6243 11462
rect 9213 11459 9279 11462
rect 10688 11520 15627 11522
rect 10688 11464 15566 11520
rect 15622 11464 15627 11520
rect 10688 11462 15627 11464
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 0 11250 480 11280
rect 0 11216 2744 11250
rect 0 11190 2836 11216
rect 0 11160 480 11190
rect 2684 11156 2836 11190
rect 9622 11188 9628 11252
rect 9692 11250 9698 11252
rect 10688 11250 10748 11462
rect 15561 11459 15627 11462
rect 21081 11522 21147 11525
rect 21081 11520 21650 11522
rect 21081 11464 21086 11520
rect 21142 11464 21650 11520
rect 21081 11462 21650 11464
rect 21081 11459 21147 11462
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 12341 11386 12407 11389
rect 14273 11386 14339 11389
rect 12341 11384 14339 11386
rect 12341 11328 12346 11384
rect 12402 11328 14278 11384
rect 14334 11328 14339 11384
rect 12341 11326 14339 11328
rect 12341 11323 12407 11326
rect 14273 11323 14339 11326
rect 9692 11190 10748 11250
rect 10869 11250 10935 11253
rect 13629 11250 13695 11253
rect 10869 11248 13695 11250
rect 10869 11192 10874 11248
rect 10930 11192 13634 11248
rect 13690 11192 13695 11248
rect 10869 11190 13695 11192
rect 9692 11188 9698 11190
rect 10869 11187 10935 11190
rect 13629 11187 13695 11190
rect 13813 11250 13879 11253
rect 17769 11250 17835 11253
rect 20345 11250 20411 11253
rect 13813 11248 20411 11250
rect 13813 11192 13818 11248
rect 13874 11192 17774 11248
rect 17830 11192 20350 11248
rect 20406 11192 20411 11248
rect 13813 11190 20411 11192
rect 21590 11250 21650 11462
rect 21725 11250 21791 11253
rect 21590 11248 21791 11250
rect 21590 11192 21730 11248
rect 21786 11192 21791 11248
rect 21590 11190 21791 11192
rect 13813 11187 13879 11190
rect 17769 11187 17835 11190
rect 20345 11187 20411 11190
rect 21725 11187 21791 11190
rect 23473 11250 23539 11253
rect 27520 11250 28000 11280
rect 23473 11248 28000 11250
rect 23473 11192 23478 11248
rect 23534 11192 28000 11248
rect 23473 11190 28000 11192
rect 23473 11187 23539 11190
rect 27520 11160 28000 11190
rect 2776 11114 2836 11156
rect 12617 11114 12683 11117
rect 21909 11114 21975 11117
rect 24577 11114 24643 11117
rect 2776 11054 12450 11114
rect 6085 10978 6151 10981
rect 9305 10978 9371 10981
rect 6085 10976 9371 10978
rect 6085 10920 6090 10976
rect 6146 10920 9310 10976
rect 9366 10920 9371 10976
rect 6085 10918 9371 10920
rect 6085 10915 6151 10918
rect 9305 10915 9371 10918
rect 10225 10978 10291 10981
rect 12390 10978 12450 11054
rect 12617 11112 24643 11114
rect 12617 11056 12622 11112
rect 12678 11056 21914 11112
rect 21970 11056 24582 11112
rect 24638 11056 24643 11112
rect 12617 11054 24643 11056
rect 12617 11051 12683 11054
rect 21909 11051 21975 11054
rect 24577 11051 24643 11054
rect 13813 10978 13879 10981
rect 10225 10976 12266 10978
rect 10225 10920 10230 10976
rect 10286 10920 12266 10976
rect 10225 10918 12266 10920
rect 12390 10976 13879 10978
rect 12390 10920 13818 10976
rect 13874 10920 13879 10976
rect 12390 10918 13879 10920
rect 10225 10915 10291 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 7557 10842 7623 10845
rect 12065 10842 12131 10845
rect 7557 10840 12131 10842
rect 7557 10784 7562 10840
rect 7618 10784 12070 10840
rect 12126 10784 12131 10840
rect 7557 10782 12131 10784
rect 12206 10842 12266 10918
rect 13813 10915 13879 10918
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 13261 10842 13327 10845
rect 12206 10840 13327 10842
rect 12206 10784 13266 10840
rect 13322 10784 13327 10840
rect 12206 10782 13327 10784
rect 7557 10779 7623 10782
rect 12065 10779 12131 10782
rect 13261 10779 13327 10782
rect 2037 10706 2103 10709
rect 4061 10706 4127 10709
rect 11697 10706 11763 10709
rect 2037 10704 3986 10706
rect 2037 10648 2042 10704
rect 2098 10648 3986 10704
rect 2037 10646 3986 10648
rect 2037 10643 2103 10646
rect 0 10570 480 10600
rect 3693 10570 3759 10573
rect 0 10568 3759 10570
rect 0 10512 3698 10568
rect 3754 10512 3759 10568
rect 0 10510 3759 10512
rect 0 10480 480 10510
rect 3693 10507 3759 10510
rect 3926 10434 3986 10646
rect 4061 10704 11763 10706
rect 4061 10648 4066 10704
rect 4122 10648 11702 10704
rect 11758 10648 11763 10704
rect 4061 10646 11763 10648
rect 4061 10643 4127 10646
rect 11697 10643 11763 10646
rect 13169 10706 13235 10709
rect 16389 10706 16455 10709
rect 13169 10704 16455 10706
rect 13169 10648 13174 10704
rect 13230 10648 16394 10704
rect 16450 10648 16455 10704
rect 13169 10646 16455 10648
rect 13169 10643 13235 10646
rect 16389 10643 16455 10646
rect 24669 10706 24735 10709
rect 24669 10704 25698 10706
rect 24669 10648 24674 10704
rect 24730 10648 25698 10704
rect 24669 10646 25698 10648
rect 24669 10643 24735 10646
rect 5533 10570 5599 10573
rect 17401 10570 17467 10573
rect 25638 10570 25698 10646
rect 27520 10570 28000 10600
rect 5533 10568 25514 10570
rect 5533 10512 5538 10568
rect 5594 10512 17406 10568
rect 17462 10512 25514 10568
rect 5533 10510 25514 10512
rect 25638 10510 28000 10570
rect 5533 10507 5599 10510
rect 17401 10507 17467 10510
rect 8753 10434 8819 10437
rect 3926 10432 8819 10434
rect 3926 10376 8758 10432
rect 8814 10376 8819 10432
rect 3926 10374 8819 10376
rect 8753 10371 8819 10374
rect 11145 10434 11211 10437
rect 19333 10434 19399 10437
rect 11145 10432 19399 10434
rect 11145 10376 11150 10432
rect 11206 10376 19338 10432
rect 19394 10376 19399 10432
rect 11145 10374 19399 10376
rect 11145 10371 11211 10374
rect 19333 10371 19399 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 2405 10298 2471 10301
rect 4521 10298 4587 10301
rect 2405 10296 4587 10298
rect 2405 10240 2410 10296
rect 2466 10240 4526 10296
rect 4582 10240 4587 10296
rect 2405 10238 4587 10240
rect 2405 10235 2471 10238
rect 4521 10235 4587 10238
rect 9438 10236 9444 10300
rect 9508 10298 9514 10300
rect 9857 10298 9923 10301
rect 9508 10296 9923 10298
rect 9508 10240 9862 10296
rect 9918 10240 9923 10296
rect 9508 10238 9923 10240
rect 9508 10236 9514 10238
rect 9857 10235 9923 10238
rect 10685 10298 10751 10301
rect 15929 10298 15995 10301
rect 17309 10298 17375 10301
rect 10685 10296 17418 10298
rect 10685 10240 10690 10296
rect 10746 10240 15934 10296
rect 15990 10240 17314 10296
rect 17370 10240 17418 10296
rect 10685 10238 17418 10240
rect 10685 10235 10751 10238
rect 15929 10235 15995 10238
rect 17309 10235 17418 10238
rect 2773 10162 2839 10165
rect 5257 10162 5323 10165
rect 8937 10162 9003 10165
rect 2773 10160 9003 10162
rect 2773 10104 2778 10160
rect 2834 10104 5262 10160
rect 5318 10104 8942 10160
rect 8998 10104 9003 10160
rect 2773 10102 9003 10104
rect 2773 10099 2839 10102
rect 5257 10099 5323 10102
rect 8937 10099 9003 10102
rect 9581 10162 9647 10165
rect 12893 10162 12959 10165
rect 9581 10160 12959 10162
rect 9581 10104 9586 10160
rect 9642 10104 12898 10160
rect 12954 10104 12959 10160
rect 9581 10102 12959 10104
rect 17358 10162 17418 10235
rect 25221 10162 25287 10165
rect 17358 10160 25287 10162
rect 17358 10104 25226 10160
rect 25282 10104 25287 10160
rect 17358 10102 25287 10104
rect 9581 10099 9647 10102
rect 12893 10099 12959 10102
rect 25221 10099 25287 10102
rect 10685 10026 10751 10029
rect 2776 10024 10751 10026
rect 2776 9968 10690 10024
rect 10746 9968 10751 10024
rect 2776 9966 10751 9968
rect 2776 9924 2836 9966
rect 10685 9963 10751 9966
rect 12893 10026 12959 10029
rect 16665 10026 16731 10029
rect 12893 10024 16731 10026
rect 12893 9968 12898 10024
rect 12954 9968 16670 10024
rect 16726 9968 16731 10024
rect 12893 9966 16731 9968
rect 12893 9963 12959 9966
rect 16665 9963 16731 9966
rect 19977 10026 20043 10029
rect 25221 10026 25287 10029
rect 19977 10024 25287 10026
rect 19977 9968 19982 10024
rect 20038 9968 25226 10024
rect 25282 9968 25287 10024
rect 19977 9966 25287 9968
rect 19977 9963 20043 9966
rect 25221 9963 25287 9966
rect 0 9890 480 9920
rect 2684 9890 2836 9924
rect 0 9864 2836 9890
rect 7189 9890 7255 9893
rect 9857 9890 9923 9893
rect 7189 9888 9923 9890
rect 0 9830 2744 9864
rect 7189 9832 7194 9888
rect 7250 9832 9862 9888
rect 9918 9832 9923 9888
rect 7189 9830 9923 9832
rect 0 9800 480 9830
rect 7189 9827 7255 9830
rect 9857 9827 9923 9830
rect 12157 9890 12223 9893
rect 13077 9890 13143 9893
rect 12157 9888 13143 9890
rect 12157 9832 12162 9888
rect 12218 9832 13082 9888
rect 13138 9832 13143 9888
rect 12157 9830 13143 9832
rect 25454 9890 25514 10510
rect 27520 10480 28000 10510
rect 27520 9890 28000 9920
rect 25454 9830 28000 9890
rect 12157 9827 12223 9830
rect 13077 9827 13143 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 27520 9800 28000 9830
rect 24277 9759 24597 9760
rect 9397 9754 9463 9757
rect 11697 9754 11763 9757
rect 9397 9752 11763 9754
rect 9397 9696 9402 9752
rect 9458 9696 11702 9752
rect 11758 9696 11763 9752
rect 9397 9694 11763 9696
rect 9397 9691 9463 9694
rect 11697 9691 11763 9694
rect 3417 9618 3483 9621
rect 12157 9618 12223 9621
rect 3417 9616 12223 9618
rect 3417 9560 3422 9616
rect 3478 9560 12162 9616
rect 12218 9560 12223 9616
rect 3417 9558 12223 9560
rect 3417 9555 3483 9558
rect 12157 9555 12223 9558
rect 12617 9618 12683 9621
rect 22461 9618 22527 9621
rect 12617 9616 22527 9618
rect 12617 9560 12622 9616
rect 12678 9560 22466 9616
rect 22522 9560 22527 9616
rect 12617 9558 22527 9560
rect 12617 9555 12683 9558
rect 22461 9555 22527 9558
rect 10133 9482 10199 9485
rect 12433 9482 12499 9485
rect 10133 9480 12499 9482
rect 10133 9424 10138 9480
rect 10194 9424 12438 9480
rect 12494 9424 12499 9480
rect 10133 9422 12499 9424
rect 10133 9419 10199 9422
rect 12433 9419 12499 9422
rect 12893 9482 12959 9485
rect 23749 9482 23815 9485
rect 12893 9480 23815 9482
rect 12893 9424 12898 9480
rect 12954 9424 23754 9480
rect 23810 9424 23815 9480
rect 12893 9422 23815 9424
rect 12893 9419 12959 9422
rect 23749 9419 23815 9422
rect 8201 9346 8267 9349
rect 3144 9344 8267 9346
rect 3144 9288 8206 9344
rect 8262 9288 8267 9344
rect 3144 9286 8267 9288
rect 0 9210 480 9240
rect 3144 9210 3204 9286
rect 8201 9283 8267 9286
rect 9990 9284 9996 9348
rect 10060 9346 10066 9348
rect 10133 9346 10199 9349
rect 10060 9344 10199 9346
rect 10060 9288 10138 9344
rect 10194 9288 10199 9344
rect 10060 9286 10199 9288
rect 10060 9284 10066 9286
rect 10133 9283 10199 9286
rect 11421 9346 11487 9349
rect 14365 9346 14431 9349
rect 11421 9344 14431 9346
rect 11421 9288 11426 9344
rect 11482 9288 14370 9344
rect 14426 9288 14431 9344
rect 11421 9286 14431 9288
rect 11421 9283 11487 9286
rect 14365 9283 14431 9286
rect 15694 9284 15700 9348
rect 15764 9346 15770 9348
rect 15837 9346 15903 9349
rect 15764 9344 15903 9346
rect 15764 9288 15842 9344
rect 15898 9288 15903 9344
rect 15764 9286 15903 9288
rect 15764 9284 15770 9286
rect 15837 9283 15903 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 21357 9212 21423 9213
rect 21357 9210 21404 9212
rect 0 9150 3204 9210
rect 21312 9208 21404 9210
rect 21312 9152 21362 9208
rect 21312 9150 21404 9152
rect 0 9120 480 9150
rect 21357 9148 21404 9150
rect 21468 9148 21474 9212
rect 24117 9210 24183 9213
rect 27520 9210 28000 9240
rect 24117 9208 28000 9210
rect 24117 9152 24122 9208
rect 24178 9152 28000 9208
rect 24117 9150 28000 9152
rect 21357 9147 21423 9148
rect 24117 9147 24183 9150
rect 27520 9120 28000 9150
rect 13077 9074 13143 9077
rect 21909 9074 21975 9077
rect 13077 9072 21975 9074
rect 13077 9016 13082 9072
rect 13138 9016 21914 9072
rect 21970 9016 21975 9072
rect 13077 9014 21975 9016
rect 13077 9011 13143 9014
rect 21909 9011 21975 9014
rect 8201 8938 8267 8941
rect 9492 8938 9690 8972
rect 10409 8938 10475 8941
rect 8201 8936 10475 8938
rect 8201 8880 8206 8936
rect 8262 8912 10414 8936
rect 8262 8880 9552 8912
rect 8201 8878 9552 8880
rect 9630 8880 10414 8912
rect 10470 8880 10475 8936
rect 9630 8878 10475 8880
rect 8201 8875 8267 8878
rect 10409 8875 10475 8878
rect 10685 8940 10751 8941
rect 10685 8936 10732 8940
rect 10796 8938 10802 8940
rect 10961 8938 11027 8941
rect 20621 8938 20687 8941
rect 10685 8880 10690 8936
rect 10685 8876 10732 8880
rect 10796 8878 10842 8938
rect 10961 8936 20687 8938
rect 10961 8880 10966 8936
rect 11022 8880 20626 8936
rect 20682 8880 20687 8936
rect 10961 8878 20687 8880
rect 10796 8876 10802 8878
rect 10685 8875 10751 8876
rect 10961 8875 11027 8878
rect 20621 8875 20687 8878
rect 9581 8802 9647 8805
rect 13813 8802 13879 8805
rect 9581 8800 13879 8802
rect 9581 8744 9586 8800
rect 9642 8744 13818 8800
rect 13874 8744 13879 8800
rect 9581 8742 13879 8744
rect 9581 8739 9647 8742
rect 13813 8739 13879 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 9397 8666 9463 8669
rect 9765 8666 9831 8669
rect 9397 8664 9831 8666
rect 9397 8608 9402 8664
rect 9458 8608 9770 8664
rect 9826 8608 9831 8664
rect 9397 8606 9831 8608
rect 9397 8603 9463 8606
rect 9765 8603 9831 8606
rect 16297 8666 16363 8669
rect 16941 8666 17007 8669
rect 16297 8664 17007 8666
rect 16297 8608 16302 8664
rect 16358 8608 16946 8664
rect 17002 8608 17007 8664
rect 16297 8606 17007 8608
rect 16297 8603 16363 8606
rect 16941 8603 17007 8606
rect 0 8530 480 8560
rect 3049 8530 3115 8533
rect 11513 8530 11579 8533
rect 12617 8530 12683 8533
rect 0 8528 3115 8530
rect 0 8472 3054 8528
rect 3110 8472 3115 8528
rect 0 8470 3115 8472
rect 0 8440 480 8470
rect 3049 8467 3115 8470
rect 9492 8528 12683 8530
rect 9492 8472 11518 8528
rect 11574 8472 12622 8528
rect 12678 8472 12683 8528
rect 9492 8470 12683 8472
rect 2497 8394 2563 8397
rect 3509 8394 3575 8397
rect 2497 8392 3575 8394
rect 2497 8336 2502 8392
rect 2558 8336 3514 8392
rect 3570 8336 3575 8392
rect 2497 8334 3575 8336
rect 2497 8331 2563 8334
rect 3509 8331 3575 8334
rect 7557 8394 7623 8397
rect 9492 8394 9552 8470
rect 11513 8467 11579 8470
rect 12617 8467 12683 8470
rect 13629 8530 13695 8533
rect 14641 8530 14707 8533
rect 13629 8528 14707 8530
rect 13629 8472 13634 8528
rect 13690 8472 14646 8528
rect 14702 8472 14707 8528
rect 13629 8470 14707 8472
rect 13629 8467 13695 8470
rect 14641 8467 14707 8470
rect 19241 8530 19307 8533
rect 21725 8530 21791 8533
rect 19241 8528 21791 8530
rect 19241 8472 19246 8528
rect 19302 8472 21730 8528
rect 21786 8472 21791 8528
rect 19241 8470 21791 8472
rect 19241 8467 19307 8470
rect 21725 8467 21791 8470
rect 24025 8530 24091 8533
rect 27520 8530 28000 8560
rect 24025 8528 28000 8530
rect 24025 8472 24030 8528
rect 24086 8472 28000 8528
rect 24025 8470 28000 8472
rect 24025 8467 24091 8470
rect 27520 8440 28000 8470
rect 11145 8394 11211 8397
rect 19425 8394 19491 8397
rect 7557 8392 9552 8394
rect 7557 8336 7562 8392
rect 7618 8336 9552 8392
rect 7557 8334 9552 8336
rect 10136 8334 10978 8394
rect 7557 8331 7623 8334
rect 3693 8258 3759 8261
rect 8109 8258 8175 8261
rect 10136 8258 10196 8334
rect 3693 8256 4906 8258
rect 3693 8200 3698 8256
rect 3754 8200 4906 8256
rect 3693 8198 4906 8200
rect 3693 8195 3759 8198
rect 2313 8122 2379 8125
rect 4705 8122 4771 8125
rect 2313 8120 4771 8122
rect 2313 8064 2318 8120
rect 2374 8064 4710 8120
rect 4766 8064 4771 8120
rect 2313 8062 4771 8064
rect 4846 8122 4906 8198
rect 8109 8256 10196 8258
rect 8109 8200 8114 8256
rect 8170 8200 10196 8256
rect 8109 8198 10196 8200
rect 8109 8195 8175 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 9397 8122 9463 8125
rect 4846 8120 9463 8122
rect 4846 8064 9402 8120
rect 9458 8064 9463 8120
rect 4846 8062 9463 8064
rect 10918 8122 10978 8334
rect 11145 8392 19491 8394
rect 11145 8336 11150 8392
rect 11206 8336 19430 8392
rect 19486 8336 19491 8392
rect 11145 8334 19491 8336
rect 11145 8331 11211 8334
rect 19425 8331 19491 8334
rect 20621 8394 20687 8397
rect 23013 8394 23079 8397
rect 23657 8394 23723 8397
rect 20621 8392 20914 8394
rect 20621 8336 20626 8392
rect 20682 8336 20914 8392
rect 20621 8334 20914 8336
rect 20621 8331 20687 8334
rect 20854 8261 20914 8334
rect 23013 8392 23723 8394
rect 23013 8336 23018 8392
rect 23074 8336 23662 8392
rect 23718 8336 23723 8392
rect 23013 8334 23723 8336
rect 23013 8331 23079 8334
rect 23657 8331 23723 8334
rect 14273 8258 14339 8261
rect 16389 8258 16455 8261
rect 14273 8256 16455 8258
rect 14273 8200 14278 8256
rect 14334 8200 16394 8256
rect 16450 8200 16455 8256
rect 14273 8198 16455 8200
rect 20854 8256 20963 8261
rect 20854 8200 20902 8256
rect 20958 8200 20963 8256
rect 20854 8198 20963 8200
rect 14273 8195 14339 8198
rect 16389 8195 16455 8198
rect 20897 8195 20963 8198
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 14733 8122 14799 8125
rect 10918 8120 14799 8122
rect 10918 8064 14738 8120
rect 14794 8064 14799 8120
rect 10918 8062 14799 8064
rect 2313 8059 2379 8062
rect 4705 8059 4771 8062
rect 9397 8059 9463 8062
rect 14733 8059 14799 8062
rect 2221 7986 2287 7989
rect 2957 7986 3023 7989
rect 10501 7986 10567 7989
rect 15929 7986 15995 7989
rect 25405 7986 25471 7989
rect 2221 7984 5090 7986
rect 2221 7928 2226 7984
rect 2282 7928 2962 7984
rect 3018 7928 5090 7984
rect 2221 7926 5090 7928
rect 2221 7923 2287 7926
rect 2957 7923 3023 7926
rect 0 7850 480 7880
rect 4245 7850 4311 7853
rect 0 7848 4311 7850
rect 0 7792 4250 7848
rect 4306 7792 4311 7848
rect 0 7790 4311 7792
rect 5030 7850 5090 7926
rect 10501 7984 25471 7986
rect 10501 7928 10506 7984
rect 10562 7928 15934 7984
rect 15990 7928 25410 7984
rect 25466 7928 25471 7984
rect 10501 7926 25471 7928
rect 10501 7923 10567 7926
rect 15929 7923 15995 7926
rect 25405 7923 25471 7926
rect 12433 7850 12499 7853
rect 14181 7850 14247 7853
rect 5030 7848 14247 7850
rect 5030 7792 12438 7848
rect 12494 7792 14186 7848
rect 14242 7792 14247 7848
rect 5030 7790 14247 7792
rect 0 7760 480 7790
rect 4245 7787 4311 7790
rect 12433 7787 12499 7790
rect 14181 7787 14247 7790
rect 14365 7850 14431 7853
rect 15837 7850 15903 7853
rect 14365 7848 15903 7850
rect 14365 7792 14370 7848
rect 14426 7792 15842 7848
rect 15898 7792 15903 7848
rect 14365 7790 15903 7792
rect 14365 7787 14431 7790
rect 15837 7787 15903 7790
rect 24761 7850 24827 7853
rect 27520 7850 28000 7880
rect 24761 7848 28000 7850
rect 24761 7792 24766 7848
rect 24822 7792 28000 7848
rect 24761 7790 28000 7792
rect 24761 7787 24827 7790
rect 27520 7760 28000 7790
rect 1853 7714 1919 7717
rect 5165 7714 5231 7717
rect 1853 7712 5231 7714
rect 1853 7656 1858 7712
rect 1914 7656 5170 7712
rect 5226 7656 5231 7712
rect 1853 7654 5231 7656
rect 1853 7651 1919 7654
rect 5165 7651 5231 7654
rect 7741 7714 7807 7717
rect 11789 7714 11855 7717
rect 18965 7714 19031 7717
rect 20713 7714 20779 7717
rect 7741 7712 14842 7714
rect 7741 7656 7746 7712
rect 7802 7656 11794 7712
rect 11850 7656 14842 7712
rect 7741 7654 14842 7656
rect 7741 7651 7807 7654
rect 11789 7651 11855 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 9213 7578 9279 7581
rect 14365 7578 14431 7581
rect 9213 7576 14431 7578
rect 9213 7520 9218 7576
rect 9274 7520 14370 7576
rect 14426 7520 14431 7576
rect 9213 7518 14431 7520
rect 9213 7515 9279 7518
rect 14365 7515 14431 7518
rect 4429 7442 4495 7445
rect 4889 7442 4955 7445
rect 6913 7442 6979 7445
rect 4429 7440 6979 7442
rect 4429 7384 4434 7440
rect 4490 7384 4894 7440
rect 4950 7384 6918 7440
rect 6974 7384 6979 7440
rect 4429 7382 6979 7384
rect 4429 7379 4495 7382
rect 4889 7379 4955 7382
rect 6913 7379 6979 7382
rect 8017 7442 8083 7445
rect 12617 7442 12683 7445
rect 8017 7440 12683 7442
rect 8017 7384 8022 7440
rect 8078 7384 12622 7440
rect 12678 7384 12683 7440
rect 8017 7382 12683 7384
rect 8017 7379 8083 7382
rect 12617 7379 12683 7382
rect 13261 7442 13327 7445
rect 13486 7442 13492 7444
rect 13261 7440 13492 7442
rect 13261 7384 13266 7440
rect 13322 7384 13492 7440
rect 13261 7382 13492 7384
rect 13261 7379 13327 7382
rect 13486 7380 13492 7382
rect 13556 7380 13562 7444
rect 14782 7442 14842 7654
rect 18965 7712 20779 7714
rect 18965 7656 18970 7712
rect 19026 7656 20718 7712
rect 20774 7656 20779 7712
rect 18965 7654 20779 7656
rect 18965 7651 19031 7654
rect 20713 7651 20779 7654
rect 21173 7714 21239 7717
rect 24117 7714 24183 7717
rect 21173 7712 24183 7714
rect 21173 7656 21178 7712
rect 21234 7656 24122 7712
rect 24178 7656 24183 7712
rect 21173 7654 24183 7656
rect 21173 7651 21239 7654
rect 24117 7651 24183 7654
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 18830 7518 24042 7578
rect 18689 7442 18755 7445
rect 18830 7442 18890 7518
rect 14782 7440 18890 7442
rect 14782 7384 18694 7440
rect 18750 7384 18890 7440
rect 14782 7382 18890 7384
rect 18965 7442 19031 7445
rect 23473 7442 23539 7445
rect 18965 7440 23539 7442
rect 18965 7384 18970 7440
rect 19026 7384 23478 7440
rect 23534 7384 23539 7440
rect 18965 7382 23539 7384
rect 23982 7442 24042 7518
rect 25221 7442 25287 7445
rect 23982 7440 25287 7442
rect 23982 7384 25226 7440
rect 25282 7384 25287 7440
rect 23982 7382 25287 7384
rect 18689 7379 18755 7382
rect 18965 7379 19031 7382
rect 23473 7379 23539 7382
rect 25221 7379 25287 7382
rect 4705 7306 4771 7309
rect 19885 7306 19951 7309
rect 4705 7304 19951 7306
rect 4705 7248 4710 7304
rect 4766 7248 19890 7304
rect 19946 7248 19951 7304
rect 4705 7246 19951 7248
rect 4705 7243 4771 7246
rect 19885 7243 19951 7246
rect 21541 7306 21607 7309
rect 23473 7306 23539 7309
rect 21541 7304 23539 7306
rect 21541 7248 21546 7304
rect 21602 7248 23478 7304
rect 23534 7248 23539 7304
rect 21541 7246 23539 7248
rect 21541 7243 21607 7246
rect 23473 7243 23539 7246
rect 0 7170 480 7200
rect 7741 7170 7807 7173
rect 9765 7170 9831 7173
rect 0 7168 7807 7170
rect 0 7112 7746 7168
rect 7802 7112 7807 7168
rect 0 7110 7807 7112
rect 0 7080 480 7110
rect 7741 7107 7807 7110
rect 7928 7168 9831 7170
rect 7928 7112 9770 7168
rect 9826 7112 9831 7168
rect 7928 7110 9831 7112
rect 7928 7034 7988 7110
rect 9765 7107 9831 7110
rect 13813 7170 13879 7173
rect 16389 7170 16455 7173
rect 13813 7168 16455 7170
rect 13813 7112 13818 7168
rect 13874 7112 16394 7168
rect 16450 7112 16455 7168
rect 13813 7110 16455 7112
rect 13813 7107 13879 7110
rect 16389 7107 16455 7110
rect 22001 7170 22067 7173
rect 27520 7170 28000 7200
rect 22001 7168 28000 7170
rect 22001 7112 22006 7168
rect 22062 7112 28000 7168
rect 22001 7110 28000 7112
rect 22001 7107 22067 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 27520 7080 28000 7110
rect 19610 7039 19930 7040
rect 1396 6974 7988 7034
rect 8109 7034 8175 7037
rect 9857 7034 9923 7037
rect 8109 7032 9923 7034
rect 8109 6976 8114 7032
rect 8170 6976 9862 7032
rect 9918 6976 9923 7032
rect 8109 6974 9923 6976
rect 0 6490 480 6520
rect 1396 6490 1456 6974
rect 8109 6971 8175 6974
rect 9857 6971 9923 6974
rect 10961 7034 11027 7037
rect 13169 7034 13235 7037
rect 10961 7032 13235 7034
rect 10961 6976 10966 7032
rect 11022 6976 13174 7032
rect 13230 6976 13235 7032
rect 10961 6974 13235 6976
rect 10961 6971 11027 6974
rect 13169 6971 13235 6974
rect 13537 7034 13603 7037
rect 18965 7034 19031 7037
rect 13537 7032 19031 7034
rect 13537 6976 13542 7032
rect 13598 6976 18970 7032
rect 19026 6976 19031 7032
rect 13537 6974 19031 6976
rect 13537 6971 13603 6974
rect 18965 6971 19031 6974
rect 3693 6898 3759 6901
rect 9673 6898 9739 6901
rect 3693 6896 9739 6898
rect 3693 6840 3698 6896
rect 3754 6840 9678 6896
rect 9734 6840 9739 6896
rect 3693 6838 9739 6840
rect 3693 6835 3759 6838
rect 9673 6835 9739 6838
rect 10041 6898 10107 6901
rect 13169 6898 13235 6901
rect 10041 6896 13235 6898
rect 10041 6840 10046 6896
rect 10102 6840 13174 6896
rect 13230 6840 13235 6896
rect 10041 6838 13235 6840
rect 10041 6835 10107 6838
rect 13169 6835 13235 6838
rect 13302 6836 13308 6900
rect 13372 6898 13378 6900
rect 23657 6898 23723 6901
rect 13372 6896 23723 6898
rect 13372 6840 23662 6896
rect 23718 6840 23723 6896
rect 13372 6838 23723 6840
rect 13372 6836 13378 6838
rect 23657 6835 23723 6838
rect 1577 6762 1643 6765
rect 9765 6762 9831 6765
rect 18873 6762 18939 6765
rect 1577 6760 9690 6762
rect 1577 6704 1582 6760
rect 1638 6704 9690 6760
rect 1577 6702 9690 6704
rect 1577 6699 1643 6702
rect 7005 6626 7071 6629
rect 9438 6626 9444 6628
rect 7005 6624 9444 6626
rect 7005 6568 7010 6624
rect 7066 6568 9444 6624
rect 7005 6566 9444 6568
rect 7005 6563 7071 6566
rect 9438 6564 9444 6566
rect 9508 6564 9514 6628
rect 9630 6626 9690 6702
rect 9765 6760 18939 6762
rect 9765 6704 9770 6760
rect 9826 6704 18878 6760
rect 18934 6704 18939 6760
rect 9765 6702 18939 6704
rect 9765 6699 9831 6702
rect 18873 6699 18939 6702
rect 12157 6626 12223 6629
rect 9630 6624 12223 6626
rect 9630 6568 12162 6624
rect 12218 6568 12223 6624
rect 9630 6566 12223 6568
rect 12157 6563 12223 6566
rect 16481 6626 16547 6629
rect 22001 6626 22067 6629
rect 16481 6624 22067 6626
rect 16481 6568 16486 6624
rect 16542 6568 22006 6624
rect 22062 6568 22067 6624
rect 16481 6566 22067 6568
rect 16481 6563 16547 6566
rect 22001 6563 22067 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 0 6430 1456 6490
rect 9397 6490 9463 6493
rect 13353 6490 13419 6493
rect 27520 6490 28000 6520
rect 9397 6488 13419 6490
rect 9397 6432 9402 6488
rect 9458 6432 13358 6488
rect 13414 6432 13419 6488
rect 9397 6430 13419 6432
rect 0 6400 480 6430
rect 9397 6427 9463 6430
rect 13353 6427 13419 6430
rect 24902 6430 28000 6490
rect 8385 6354 8451 6357
rect 13629 6354 13695 6357
rect 8385 6352 13695 6354
rect 8385 6296 8390 6352
rect 8446 6296 13634 6352
rect 13690 6296 13695 6352
rect 8385 6294 13695 6296
rect 8385 6291 8451 6294
rect 13629 6291 13695 6294
rect 16849 6354 16915 6357
rect 24902 6354 24962 6430
rect 27520 6400 28000 6430
rect 16849 6352 24962 6354
rect 16849 6296 16854 6352
rect 16910 6296 24962 6352
rect 16849 6294 24962 6296
rect 16849 6291 16915 6294
rect 2497 6218 2563 6221
rect 16573 6218 16639 6221
rect 16849 6218 16915 6221
rect 24209 6218 24275 6221
rect 2497 6216 24275 6218
rect 2497 6160 2502 6216
rect 2558 6160 16578 6216
rect 16634 6160 16854 6216
rect 16910 6160 24214 6216
rect 24270 6160 24275 6216
rect 2497 6158 24275 6160
rect 2497 6155 2563 6158
rect 16573 6155 16639 6158
rect 16849 6155 16915 6158
rect 24209 6155 24275 6158
rect 6085 6082 6151 6085
rect 9765 6082 9831 6085
rect 10041 6084 10107 6085
rect 9990 6082 9996 6084
rect 6085 6080 9831 6082
rect 6085 6024 6090 6080
rect 6146 6024 9770 6080
rect 9826 6024 9831 6080
rect 6085 6022 9831 6024
rect 9950 6022 9996 6082
rect 10060 6080 10107 6084
rect 10102 6024 10107 6080
rect 6085 6019 6151 6022
rect 9765 6019 9831 6022
rect 9990 6020 9996 6022
rect 10060 6020 10107 6024
rect 10041 6019 10107 6020
rect 10777 6082 10843 6085
rect 14549 6082 14615 6085
rect 10777 6080 19258 6082
rect 10777 6024 10782 6080
rect 10838 6024 14554 6080
rect 14610 6024 19258 6080
rect 10777 6022 19258 6024
rect 10777 6019 10843 6022
rect 14549 6019 14615 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 1393 5946 1459 5949
rect 1393 5944 7666 5946
rect 1393 5888 1398 5944
rect 1454 5888 7666 5944
rect 1393 5886 7666 5888
rect 1393 5883 1459 5886
rect 0 5810 480 5840
rect 7465 5810 7531 5813
rect 0 5808 7531 5810
rect 0 5752 7470 5808
rect 7526 5752 7531 5808
rect 0 5750 7531 5752
rect 7606 5810 7666 5886
rect 15377 5810 15443 5813
rect 7606 5808 15443 5810
rect 7606 5752 15382 5808
rect 15438 5752 15443 5808
rect 7606 5750 15443 5752
rect 19198 5810 19258 6022
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 21357 5810 21423 5813
rect 19198 5808 21423 5810
rect 19198 5752 21362 5808
rect 21418 5752 21423 5808
rect 19198 5750 21423 5752
rect 0 5720 480 5750
rect 7465 5747 7531 5750
rect 15377 5747 15443 5750
rect 21357 5747 21423 5750
rect 23657 5810 23723 5813
rect 27520 5810 28000 5840
rect 23657 5808 28000 5810
rect 23657 5752 23662 5808
rect 23718 5752 28000 5808
rect 23657 5750 28000 5752
rect 23657 5747 23723 5750
rect 27520 5720 28000 5750
rect 2037 5674 2103 5677
rect 4521 5674 4587 5677
rect 2037 5672 4587 5674
rect 2037 5616 2042 5672
rect 2098 5616 4526 5672
rect 4582 5616 4587 5672
rect 2037 5614 4587 5616
rect 2037 5611 2103 5614
rect 4521 5611 4587 5614
rect 6821 5674 6887 5677
rect 9213 5674 9279 5677
rect 6821 5672 9279 5674
rect 6821 5616 6826 5672
rect 6882 5616 9218 5672
rect 9274 5616 9279 5672
rect 6821 5614 9279 5616
rect 6821 5611 6887 5614
rect 9213 5611 9279 5614
rect 13537 5674 13603 5677
rect 19425 5674 19491 5677
rect 13537 5672 19491 5674
rect 13537 5616 13542 5672
rect 13598 5616 19430 5672
rect 19486 5616 19491 5672
rect 13537 5614 19491 5616
rect 13537 5611 13603 5614
rect 19425 5611 19491 5614
rect 13353 5540 13419 5541
rect 13302 5476 13308 5540
rect 13372 5538 13419 5540
rect 13372 5536 13464 5538
rect 13414 5480 13464 5536
rect 13372 5478 13464 5480
rect 13372 5476 13419 5478
rect 13353 5475 13419 5476
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 6361 5402 6427 5405
rect 11421 5402 11487 5405
rect 24025 5402 24091 5405
rect 6361 5400 11487 5402
rect 6361 5344 6366 5400
rect 6422 5344 11426 5400
rect 11482 5344 11487 5400
rect 6361 5342 11487 5344
rect 6361 5339 6427 5342
rect 11421 5339 11487 5342
rect 20486 5400 24091 5402
rect 20486 5344 24030 5400
rect 24086 5344 24091 5400
rect 20486 5342 24091 5344
rect 20486 5269 20546 5342
rect 24025 5339 24091 5342
rect 6545 5266 6611 5269
rect 9029 5266 9095 5269
rect 6545 5264 9095 5266
rect 6545 5208 6550 5264
rect 6606 5208 9034 5264
rect 9090 5208 9095 5264
rect 6545 5206 9095 5208
rect 6545 5203 6611 5206
rect 9029 5203 9095 5206
rect 9213 5266 9279 5269
rect 20437 5266 20546 5269
rect 9213 5264 20546 5266
rect 9213 5208 9218 5264
rect 9274 5208 20442 5264
rect 20498 5208 20546 5264
rect 9213 5206 20546 5208
rect 9213 5203 9279 5206
rect 20437 5203 20503 5206
rect 0 5130 480 5160
rect 1485 5130 1551 5133
rect 0 5128 1551 5130
rect 0 5072 1490 5128
rect 1546 5072 1551 5128
rect 0 5070 1551 5072
rect 0 5040 480 5070
rect 1485 5067 1551 5070
rect 4061 5130 4127 5133
rect 18781 5130 18847 5133
rect 4061 5128 18847 5130
rect 4061 5072 4066 5128
rect 4122 5072 18786 5128
rect 18842 5072 18847 5128
rect 4061 5070 18847 5072
rect 4061 5067 4127 5070
rect 18781 5067 18847 5070
rect 20161 5130 20227 5133
rect 23473 5130 23539 5133
rect 27520 5130 28000 5160
rect 20161 5128 23306 5130
rect 20161 5072 20166 5128
rect 20222 5072 23306 5128
rect 20161 5070 23306 5072
rect 20161 5067 20227 5070
rect 6637 4994 6703 4997
rect 9121 4994 9187 4997
rect 6637 4992 9187 4994
rect 6637 4936 6642 4992
rect 6698 4936 9126 4992
rect 9182 4936 9187 4992
rect 6637 4934 9187 4936
rect 6637 4931 6703 4934
rect 9121 4931 9187 4934
rect 10777 4994 10843 4997
rect 16481 4994 16547 4997
rect 10777 4992 16547 4994
rect 10777 4936 10782 4992
rect 10838 4936 16486 4992
rect 16542 4936 16547 4992
rect 10777 4934 16547 4936
rect 23246 4994 23306 5070
rect 23473 5128 28000 5130
rect 23473 5072 23478 5128
rect 23534 5072 28000 5128
rect 23473 5070 28000 5072
rect 23473 5067 23539 5070
rect 27520 5040 28000 5070
rect 24945 4994 25011 4997
rect 23246 4992 25011 4994
rect 23246 4936 24950 4992
rect 25006 4936 25011 4992
rect 23246 4934 25011 4936
rect 10777 4931 10843 4934
rect 16481 4931 16547 4934
rect 24945 4931 25011 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 5993 4858 6059 4861
rect 7925 4858 7991 4861
rect 16113 4858 16179 4861
rect 5993 4856 7991 4858
rect 5993 4800 5998 4856
rect 6054 4800 7930 4856
rect 7986 4800 7991 4856
rect 5993 4798 7991 4800
rect 5993 4795 6059 4798
rect 7925 4795 7991 4798
rect 10688 4856 16179 4858
rect 10688 4800 16118 4856
rect 16174 4800 16179 4856
rect 10688 4798 16179 4800
rect 1669 4722 1735 4725
rect 8293 4722 8359 4725
rect 10688 4722 10748 4798
rect 16113 4795 16179 4798
rect 1669 4720 7666 4722
rect 1669 4664 1674 4720
rect 1730 4664 7666 4720
rect 1669 4662 7666 4664
rect 1669 4659 1735 4662
rect 0 4450 480 4480
rect 5441 4450 5507 4453
rect 0 4448 5507 4450
rect 0 4392 5446 4448
rect 5502 4392 5507 4448
rect 0 4390 5507 4392
rect 0 4360 480 4390
rect 5441 4387 5507 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 7606 4178 7666 4662
rect 8293 4720 10748 4722
rect 8293 4664 8298 4720
rect 8354 4664 10748 4720
rect 8293 4662 10748 4664
rect 11421 4722 11487 4725
rect 11421 4720 24962 4722
rect 11421 4664 11426 4720
rect 11482 4664 24962 4720
rect 11421 4662 24962 4664
rect 8293 4659 8359 4662
rect 11421 4659 11487 4662
rect 7925 4586 7991 4589
rect 8937 4586 9003 4589
rect 20253 4586 20319 4589
rect 7925 4584 20319 4586
rect 7925 4528 7930 4584
rect 7986 4528 8942 4584
rect 8998 4528 20258 4584
rect 20314 4528 20319 4584
rect 7925 4526 20319 4528
rect 7925 4523 7991 4526
rect 8937 4523 9003 4526
rect 20253 4523 20319 4526
rect 8017 4450 8083 4453
rect 11421 4450 11487 4453
rect 8017 4448 11487 4450
rect 8017 4392 8022 4448
rect 8078 4392 11426 4448
rect 11482 4392 11487 4448
rect 8017 4390 11487 4392
rect 24902 4450 24962 4662
rect 27520 4450 28000 4480
rect 24902 4390 28000 4450
rect 8017 4387 8083 4390
rect 11421 4387 11487 4390
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 27520 4360 28000 4390
rect 24277 4319 24597 4320
rect 18781 4314 18847 4317
rect 20713 4314 20779 4317
rect 23749 4314 23815 4317
rect 18781 4312 23815 4314
rect 18781 4256 18786 4312
rect 18842 4256 20718 4312
rect 20774 4256 23754 4312
rect 23810 4256 23815 4312
rect 18781 4254 23815 4256
rect 18781 4251 18847 4254
rect 20713 4251 20779 4254
rect 23749 4251 23815 4254
rect 15285 4178 15351 4181
rect 7606 4176 15351 4178
rect 7606 4120 15290 4176
rect 15346 4120 15351 4176
rect 7606 4118 15351 4120
rect 15285 4115 15351 4118
rect 22645 4178 22711 4181
rect 25313 4178 25379 4181
rect 22645 4176 25379 4178
rect 22645 4120 22650 4176
rect 22706 4120 25318 4176
rect 25374 4120 25379 4176
rect 22645 4118 25379 4120
rect 22645 4115 22711 4118
rect 25313 4115 25379 4118
rect 7373 4042 7439 4045
rect 9765 4042 9831 4045
rect 7373 4040 9831 4042
rect 7373 3984 7378 4040
rect 7434 3984 9770 4040
rect 9826 3984 9831 4040
rect 7373 3982 9831 3984
rect 7373 3979 7439 3982
rect 9765 3979 9831 3982
rect 13721 4042 13787 4045
rect 15285 4042 15351 4045
rect 13721 4040 15351 4042
rect 13721 3984 13726 4040
rect 13782 3984 15290 4040
rect 15346 3984 15351 4040
rect 13721 3982 15351 3984
rect 13721 3979 13787 3982
rect 15285 3979 15351 3982
rect 15929 4042 15995 4045
rect 17125 4042 17191 4045
rect 15929 4040 17191 4042
rect 15929 3984 15934 4040
rect 15990 3984 17130 4040
rect 17186 3984 17191 4040
rect 15929 3982 17191 3984
rect 15929 3979 15995 3982
rect 17125 3979 17191 3982
rect 17309 4042 17375 4045
rect 27613 4042 27679 4045
rect 17309 4040 27679 4042
rect 17309 3984 17314 4040
rect 17370 3984 27618 4040
rect 27674 3984 27679 4040
rect 17309 3982 27679 3984
rect 17309 3979 17375 3982
rect 27613 3979 27679 3982
rect 5073 3906 5139 3909
rect 6729 3906 6795 3909
rect 5073 3904 6795 3906
rect 5073 3848 5078 3904
rect 5134 3848 6734 3904
rect 6790 3848 6795 3904
rect 5073 3846 6795 3848
rect 5073 3843 5139 3846
rect 6729 3843 6795 3846
rect 7925 3906 7991 3909
rect 9622 3906 9628 3908
rect 7925 3904 9628 3906
rect 7925 3848 7930 3904
rect 7986 3848 9628 3904
rect 7925 3846 9628 3848
rect 7925 3843 7991 3846
rect 9622 3844 9628 3846
rect 9692 3844 9698 3908
rect 11421 3906 11487 3909
rect 13261 3906 13327 3909
rect 11421 3904 13327 3906
rect 11421 3848 11426 3904
rect 11482 3848 13266 3904
rect 13322 3848 13327 3904
rect 11421 3846 13327 3848
rect 11421 3843 11487 3846
rect 13261 3843 13327 3846
rect 13537 3906 13603 3909
rect 18229 3906 18295 3909
rect 13537 3904 18295 3906
rect 13537 3848 13542 3904
rect 13598 3848 18234 3904
rect 18290 3848 18295 3904
rect 13537 3846 18295 3848
rect 13537 3843 13603 3846
rect 18229 3843 18295 3846
rect 21173 3906 21239 3909
rect 23657 3906 23723 3909
rect 24117 3906 24183 3909
rect 21173 3904 23723 3906
rect 21173 3848 21178 3904
rect 21234 3848 23662 3904
rect 23718 3848 23723 3904
rect 21173 3846 23723 3848
rect 21173 3843 21239 3846
rect 23657 3843 23723 3846
rect 23798 3904 24183 3906
rect 23798 3848 24122 3904
rect 24178 3848 24183 3904
rect 23798 3846 24183 3848
rect 10277 3840 10597 3841
rect 0 3770 480 3800
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 2773 3770 2839 3773
rect 0 3768 2839 3770
rect 0 3712 2778 3768
rect 2834 3712 2839 3768
rect 0 3710 2839 3712
rect 0 3680 480 3710
rect 2773 3707 2839 3710
rect 3141 3770 3207 3773
rect 6085 3770 6151 3773
rect 7189 3770 7255 3773
rect 8661 3770 8727 3773
rect 12157 3770 12223 3773
rect 15653 3770 15719 3773
rect 3141 3768 8727 3770
rect 3141 3712 3146 3768
rect 3202 3712 6090 3768
rect 6146 3712 7194 3768
rect 7250 3712 8666 3768
rect 8722 3712 8727 3768
rect 3141 3710 8727 3712
rect 3141 3707 3207 3710
rect 6085 3707 6151 3710
rect 7189 3707 7255 3710
rect 8661 3707 8727 3710
rect 10688 3768 15719 3770
rect 10688 3712 12162 3768
rect 12218 3712 15658 3768
rect 15714 3712 15719 3768
rect 10688 3710 15719 3712
rect 9029 3634 9095 3637
rect 10688 3634 10748 3710
rect 12157 3707 12223 3710
rect 15653 3707 15719 3710
rect 21449 3770 21515 3773
rect 23798 3770 23858 3846
rect 24117 3843 24183 3846
rect 21449 3768 23858 3770
rect 21449 3712 21454 3768
rect 21510 3712 23858 3768
rect 21449 3710 23858 3712
rect 23933 3770 23999 3773
rect 27520 3770 28000 3800
rect 23933 3768 28000 3770
rect 23933 3712 23938 3768
rect 23994 3712 28000 3768
rect 23933 3710 28000 3712
rect 21449 3707 21515 3710
rect 23933 3707 23999 3710
rect 27520 3680 28000 3710
rect 9029 3632 10748 3634
rect 9029 3576 9034 3632
rect 9090 3576 10748 3632
rect 9029 3574 10748 3576
rect 11145 3634 11211 3637
rect 12709 3634 12775 3637
rect 11145 3632 12775 3634
rect 11145 3576 11150 3632
rect 11206 3576 12714 3632
rect 12770 3576 12775 3632
rect 11145 3574 12775 3576
rect 9029 3571 9095 3574
rect 11145 3571 11211 3574
rect 12709 3571 12775 3574
rect 12985 3634 13051 3637
rect 20621 3634 20687 3637
rect 12985 3632 20687 3634
rect 12985 3576 12990 3632
rect 13046 3576 20626 3632
rect 20682 3576 20687 3632
rect 12985 3574 20687 3576
rect 12985 3571 13051 3574
rect 20621 3571 20687 3574
rect 21357 3634 21423 3637
rect 26049 3634 26115 3637
rect 21357 3632 26115 3634
rect 21357 3576 21362 3632
rect 21418 3576 26054 3632
rect 26110 3576 26115 3632
rect 21357 3574 26115 3576
rect 21357 3571 21423 3574
rect 26049 3571 26115 3574
rect 7649 3498 7715 3501
rect 9121 3498 9187 3501
rect 10225 3498 10291 3501
rect 13813 3498 13879 3501
rect 7649 3496 13879 3498
rect 7649 3440 7654 3496
rect 7710 3440 9126 3496
rect 9182 3440 10230 3496
rect 10286 3440 13818 3496
rect 13874 3440 13879 3496
rect 7649 3438 13879 3440
rect 7649 3435 7715 3438
rect 9121 3435 9187 3438
rect 10225 3435 10291 3438
rect 13813 3435 13879 3438
rect 18137 3498 18203 3501
rect 21449 3498 21515 3501
rect 18137 3496 21515 3498
rect 18137 3440 18142 3496
rect 18198 3440 21454 3496
rect 21510 3440 21515 3496
rect 18137 3438 21515 3440
rect 18137 3435 18203 3438
rect 21449 3435 21515 3438
rect 22645 3498 22711 3501
rect 25865 3498 25931 3501
rect 22645 3496 25931 3498
rect 22645 3440 22650 3496
rect 22706 3440 25870 3496
rect 25926 3440 25931 3496
rect 22645 3438 25931 3440
rect 22645 3435 22711 3438
rect 25865 3435 25931 3438
rect 9673 3362 9739 3365
rect 10041 3362 10107 3365
rect 9673 3360 10107 3362
rect 9673 3304 9678 3360
rect 9734 3304 10046 3360
rect 10102 3304 10107 3360
rect 9673 3302 10107 3304
rect 9673 3299 9739 3302
rect 10041 3299 10107 3302
rect 13486 3300 13492 3364
rect 13556 3362 13562 3364
rect 13721 3362 13787 3365
rect 13556 3360 13787 3362
rect 13556 3304 13726 3360
rect 13782 3304 13787 3360
rect 13556 3302 13787 3304
rect 13556 3300 13562 3302
rect 13721 3299 13787 3302
rect 16297 3362 16363 3365
rect 20529 3362 20595 3365
rect 16297 3360 20595 3362
rect 16297 3304 16302 3360
rect 16358 3304 20534 3360
rect 20590 3304 20595 3360
rect 16297 3302 20595 3304
rect 16297 3299 16363 3302
rect 20529 3299 20595 3302
rect 21817 3362 21883 3365
rect 22369 3362 22435 3365
rect 21817 3360 22435 3362
rect 21817 3304 21822 3360
rect 21878 3304 22374 3360
rect 22430 3304 22435 3360
rect 21817 3302 22435 3304
rect 21817 3299 21883 3302
rect 22369 3299 22435 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 8385 3226 8451 3229
rect 11789 3226 11855 3229
rect 8385 3224 11855 3226
rect 8385 3168 8390 3224
rect 8446 3168 11794 3224
rect 11850 3168 11855 3224
rect 8385 3166 11855 3168
rect 8385 3163 8451 3166
rect 11789 3163 11855 3166
rect 20713 3226 20779 3229
rect 24025 3226 24091 3229
rect 20713 3224 24091 3226
rect 20713 3168 20718 3224
rect 20774 3168 24030 3224
rect 24086 3168 24091 3224
rect 20713 3166 24091 3168
rect 20713 3163 20779 3166
rect 24025 3163 24091 3166
rect 0 3090 480 3120
rect 3417 3090 3483 3093
rect 0 3088 3483 3090
rect 0 3032 3422 3088
rect 3478 3032 3483 3088
rect 0 3030 3483 3032
rect 0 3000 480 3030
rect 3417 3027 3483 3030
rect 5349 3090 5415 3093
rect 8201 3090 8267 3093
rect 5349 3088 8267 3090
rect 5349 3032 5354 3088
rect 5410 3032 8206 3088
rect 8262 3032 8267 3088
rect 5349 3030 8267 3032
rect 5349 3027 5415 3030
rect 8201 3027 8267 3030
rect 9673 3090 9739 3093
rect 12433 3090 12499 3093
rect 9673 3088 12499 3090
rect 9673 3032 9678 3088
rect 9734 3032 12438 3088
rect 12494 3032 12499 3088
rect 9673 3030 12499 3032
rect 9673 3027 9739 3030
rect 12433 3027 12499 3030
rect 18413 3090 18479 3093
rect 21817 3090 21883 3093
rect 18413 3088 21883 3090
rect 18413 3032 18418 3088
rect 18474 3032 21822 3088
rect 21878 3032 21883 3088
rect 18413 3030 21883 3032
rect 18413 3027 18479 3030
rect 21817 3027 21883 3030
rect 24025 3090 24091 3093
rect 27520 3090 28000 3120
rect 24025 3088 28000 3090
rect 24025 3032 24030 3088
rect 24086 3032 28000 3088
rect 24025 3030 28000 3032
rect 24025 3027 24091 3030
rect 27520 3000 28000 3030
rect 1853 2954 1919 2957
rect 3049 2954 3115 2957
rect 5625 2954 5691 2957
rect 1853 2952 5691 2954
rect 1853 2896 1858 2952
rect 1914 2896 3054 2952
rect 3110 2896 5630 2952
rect 5686 2896 5691 2952
rect 1853 2894 5691 2896
rect 1853 2891 1919 2894
rect 3049 2891 3115 2894
rect 5625 2891 5691 2894
rect 9213 2954 9279 2957
rect 11421 2954 11487 2957
rect 17769 2954 17835 2957
rect 9213 2952 10794 2954
rect 9213 2896 9218 2952
rect 9274 2896 10794 2952
rect 9213 2894 10794 2896
rect 9213 2891 9279 2894
rect 841 2818 907 2821
rect 5349 2818 5415 2821
rect 841 2816 5415 2818
rect 841 2760 846 2816
rect 902 2760 5354 2816
rect 5410 2760 5415 2816
rect 841 2758 5415 2760
rect 841 2755 907 2758
rect 5349 2755 5415 2758
rect 5533 2818 5599 2821
rect 6177 2818 6243 2821
rect 5533 2816 6243 2818
rect 5533 2760 5538 2816
rect 5594 2760 6182 2816
rect 6238 2760 6243 2816
rect 5533 2758 6243 2760
rect 5533 2755 5599 2758
rect 6177 2755 6243 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 2313 2682 2379 2685
rect 6913 2682 6979 2685
rect 2313 2680 6979 2682
rect 2313 2624 2318 2680
rect 2374 2624 6918 2680
rect 6974 2624 6979 2680
rect 2313 2622 6979 2624
rect 10734 2682 10794 2894
rect 11421 2952 17835 2954
rect 11421 2896 11426 2952
rect 11482 2896 17774 2952
rect 17830 2896 17835 2952
rect 11421 2894 17835 2896
rect 11421 2891 11487 2894
rect 17769 2891 17835 2894
rect 19885 2954 19951 2957
rect 24577 2954 24643 2957
rect 19885 2952 24643 2954
rect 19885 2896 19890 2952
rect 19946 2896 24582 2952
rect 24638 2896 24643 2952
rect 19885 2894 24643 2896
rect 19885 2891 19951 2894
rect 24577 2891 24643 2894
rect 11973 2818 12039 2821
rect 13997 2818 14063 2821
rect 15561 2818 15627 2821
rect 11973 2816 15627 2818
rect 11973 2760 11978 2816
rect 12034 2760 14002 2816
rect 14058 2760 15566 2816
rect 15622 2760 15627 2816
rect 11973 2758 15627 2760
rect 11973 2755 12039 2758
rect 13997 2755 14063 2758
rect 15561 2755 15627 2758
rect 20345 2818 20411 2821
rect 22645 2818 22711 2821
rect 26509 2818 26575 2821
rect 20345 2816 22570 2818
rect 20345 2760 20350 2816
rect 20406 2760 22570 2816
rect 20345 2758 22570 2760
rect 20345 2755 20411 2758
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 14733 2682 14799 2685
rect 10734 2680 14799 2682
rect 10734 2624 14738 2680
rect 14794 2624 14799 2680
rect 10734 2622 14799 2624
rect 2313 2619 2379 2622
rect 6913 2619 6979 2622
rect 14733 2619 14799 2622
rect 15009 2682 15075 2685
rect 16849 2682 16915 2685
rect 15009 2680 16915 2682
rect 15009 2624 15014 2680
rect 15070 2624 16854 2680
rect 16910 2624 16915 2680
rect 15009 2622 16915 2624
rect 22510 2682 22570 2758
rect 22645 2816 26575 2818
rect 22645 2760 22650 2816
rect 22706 2760 26514 2816
rect 26570 2760 26575 2816
rect 22645 2758 26575 2760
rect 22645 2755 22711 2758
rect 26509 2755 26575 2758
rect 23013 2682 23079 2685
rect 22510 2680 23079 2682
rect 22510 2624 23018 2680
rect 23074 2624 23079 2680
rect 22510 2622 23079 2624
rect 15009 2619 15075 2622
rect 16849 2619 16915 2622
rect 23013 2619 23079 2622
rect 1945 2546 2011 2549
rect 11237 2546 11303 2549
rect 17677 2546 17743 2549
rect 1945 2544 11303 2546
rect 1945 2488 1950 2544
rect 2006 2488 11242 2544
rect 11298 2488 11303 2544
rect 1945 2486 11303 2488
rect 1945 2483 2011 2486
rect 11237 2483 11303 2486
rect 11424 2544 17743 2546
rect 11424 2488 17682 2544
rect 17738 2488 17743 2544
rect 11424 2486 17743 2488
rect 0 2410 480 2440
rect 7465 2410 7531 2413
rect 11424 2410 11484 2486
rect 17677 2483 17743 2486
rect 0 2350 6562 2410
rect 0 2320 480 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 6502 2138 6562 2350
rect 7465 2408 11484 2410
rect 7465 2352 7470 2408
rect 7526 2352 11484 2408
rect 7465 2350 11484 2352
rect 11697 2410 11763 2413
rect 24485 2410 24551 2413
rect 27520 2410 28000 2440
rect 11697 2408 17234 2410
rect 11697 2352 11702 2408
rect 11758 2352 17234 2408
rect 11697 2350 17234 2352
rect 7465 2347 7531 2350
rect 11697 2347 11763 2350
rect 6729 2274 6795 2277
rect 9765 2274 9831 2277
rect 6729 2272 9831 2274
rect 6729 2216 6734 2272
rect 6790 2216 9770 2272
rect 9826 2216 9831 2272
rect 6729 2214 9831 2216
rect 17174 2274 17234 2350
rect 24485 2408 28000 2410
rect 24485 2352 24490 2408
rect 24546 2352 28000 2408
rect 24485 2350 28000 2352
rect 24485 2347 24551 2350
rect 27520 2320 28000 2350
rect 23933 2274 23999 2277
rect 17174 2272 23999 2274
rect 17174 2216 23938 2272
rect 23994 2216 23999 2272
rect 17174 2214 23999 2216
rect 6729 2211 6795 2214
rect 9765 2211 9831 2214
rect 23933 2211 23999 2214
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 8661 2138 8727 2141
rect 14365 2138 14431 2141
rect 23473 2138 23539 2141
rect 6502 2078 8586 2138
rect 4613 2002 4679 2005
rect 8293 2002 8359 2005
rect 4613 2000 8359 2002
rect 4613 1944 4618 2000
rect 4674 1944 8298 2000
rect 8354 1944 8359 2000
rect 4613 1942 8359 1944
rect 8526 2002 8586 2078
rect 8661 2136 14431 2138
rect 8661 2080 8666 2136
rect 8722 2080 14370 2136
rect 14426 2080 14431 2136
rect 8661 2078 14431 2080
rect 8661 2075 8727 2078
rect 14365 2075 14431 2078
rect 20302 2136 23539 2138
rect 20302 2080 23478 2136
rect 23534 2080 23539 2136
rect 20302 2078 23539 2080
rect 10869 2002 10935 2005
rect 8526 2000 10935 2002
rect 8526 1944 10874 2000
rect 10930 1944 10935 2000
rect 8526 1942 10935 1944
rect 4613 1939 4679 1942
rect 8293 1939 8359 1942
rect 10869 1939 10935 1942
rect 14733 2002 14799 2005
rect 17309 2002 17375 2005
rect 14733 2000 17375 2002
rect 14733 1944 14738 2000
rect 14794 1944 17314 2000
rect 17370 1944 17375 2000
rect 14733 1942 17375 1944
rect 14733 1939 14799 1942
rect 17309 1939 17375 1942
rect 9857 1866 9923 1869
rect 20069 1866 20135 1869
rect 9857 1864 20135 1866
rect 9857 1808 9862 1864
rect 9918 1808 20074 1864
rect 20130 1808 20135 1864
rect 9857 1806 20135 1808
rect 9857 1803 9923 1806
rect 20069 1803 20135 1806
rect 0 1730 480 1760
rect 3918 1730 3924 1732
rect 0 1670 3924 1730
rect 0 1640 480 1670
rect 3918 1668 3924 1670
rect 3988 1668 3994 1732
rect 10685 1730 10751 1733
rect 18321 1730 18387 1733
rect 10685 1728 18387 1730
rect 10685 1672 10690 1728
rect 10746 1672 18326 1728
rect 18382 1672 18387 1728
rect 10685 1670 18387 1672
rect 10685 1667 10751 1670
rect 18321 1667 18387 1670
rect 3417 1594 3483 1597
rect 11421 1594 11487 1597
rect 3417 1592 11487 1594
rect 3417 1536 3422 1592
rect 3478 1536 11426 1592
rect 11482 1536 11487 1592
rect 3417 1534 11487 1536
rect 3417 1531 3483 1534
rect 11421 1531 11487 1534
rect 11605 1594 11671 1597
rect 16573 1594 16639 1597
rect 20302 1594 20362 2078
rect 23473 2075 23539 2078
rect 27520 1730 28000 1760
rect 11605 1592 16639 1594
rect 11605 1536 11610 1592
rect 11666 1536 16578 1592
rect 16634 1536 16639 1592
rect 11605 1534 16639 1536
rect 11605 1531 11671 1534
rect 16573 1531 16639 1534
rect 17174 1534 20362 1594
rect 27478 1640 28000 1730
rect 9397 1458 9463 1461
rect 17174 1458 17234 1534
rect 9397 1456 17234 1458
rect 9397 1400 9402 1456
rect 9458 1400 17234 1456
rect 9397 1398 17234 1400
rect 17309 1458 17375 1461
rect 27478 1458 27538 1640
rect 17309 1456 27538 1458
rect 17309 1400 17314 1456
rect 17370 1400 27538 1456
rect 17309 1398 27538 1400
rect 9397 1395 9463 1398
rect 17309 1395 17375 1398
rect 3693 1322 3759 1325
rect 14549 1322 14615 1325
rect 3693 1320 14615 1322
rect 3693 1264 3698 1320
rect 3754 1264 14554 1320
rect 14610 1264 14615 1320
rect 3693 1262 14615 1264
rect 3693 1259 3759 1262
rect 14549 1259 14615 1262
rect 10685 1188 10751 1189
rect 10685 1186 10732 1188
rect 10640 1184 10732 1186
rect 10640 1128 10690 1184
rect 10640 1126 10732 1128
rect 10685 1124 10732 1126
rect 10796 1124 10802 1188
rect 10685 1123 10751 1124
rect 0 1050 480 1080
rect 2957 1050 3023 1053
rect 0 1048 3023 1050
rect 0 992 2962 1048
rect 3018 992 3023 1048
rect 0 990 3023 992
rect 0 960 480 990
rect 2957 987 3023 990
rect 23657 1050 23723 1053
rect 27520 1050 28000 1080
rect 23657 1048 28000 1050
rect 23657 992 23662 1048
rect 23718 992 28000 1048
rect 23657 990 28000 992
rect 23657 987 23723 990
rect 27520 960 28000 990
rect 0 370 480 400
rect 3693 370 3759 373
rect 0 368 3759 370
rect 0 312 3698 368
rect 3754 312 3759 368
rect 0 310 3759 312
rect 0 280 480 310
rect 3693 307 3759 310
rect 18781 370 18847 373
rect 27520 370 28000 400
rect 18781 368 28000 370
rect 18781 312 18786 368
rect 18842 312 28000 368
rect 18781 310 28000 312
rect 18781 307 18847 310
rect 27520 280 28000 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 21404 19892 21468 19956
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 21404 14996 21468 15060
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 9812 12140 9876 12204
rect 13308 12140 13372 12204
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 9260 11596 9324 11660
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 9628 11188 9692 11252
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 9444 10236 9508 10300
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 9996 9284 10060 9348
rect 15700 9284 15764 9348
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 21404 9208 21468 9212
rect 21404 9152 21418 9208
rect 21418 9152 21468 9208
rect 21404 9148 21468 9152
rect 10732 8936 10796 8940
rect 10732 8880 10746 8936
rect 10746 8880 10796 8936
rect 10732 8876 10796 8880
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 13492 7380 13556 7444
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 13308 6836 13372 6900
rect 9444 6564 9508 6628
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 9996 6080 10060 6084
rect 9996 6024 10046 6080
rect 10046 6024 10060 6080
rect 9996 6020 10060 6024
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 13308 5536 13372 5540
rect 13308 5480 13358 5536
rect 13358 5480 13372 5536
rect 13308 5476 13372 5480
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 9628 3844 9692 3908
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 13492 3300 13556 3364
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 3924 1668 3988 1732
rect 10732 1184 10796 1188
rect 10732 1128 10746 1184
rect 10746 1128 10796 1184
rect 10732 1124 10796 1128
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 9262 12550 9874 12610
rect 9262 11661 9322 12550
rect 9814 12205 9874 12550
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 9811 12204 9877 12205
rect 9811 12140 9812 12204
rect 9876 12140 9877 12204
rect 9811 12139 9877 12140
rect 9259 11660 9325 11661
rect 9259 11596 9260 11660
rect 9324 11596 9325 11660
rect 9259 11595 9325 11596
rect 10277 11456 10597 12480
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 13307 12204 13373 12205
rect 13307 12140 13308 12204
rect 13372 12140 13373 12204
rect 13307 12139 13373 12140
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 9627 11252 9693 11253
rect 9627 11188 9628 11252
rect 9692 11188 9693 11252
rect 9627 11187 9693 11188
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 9443 10300 9509 10301
rect 9443 10236 9444 10300
rect 9508 10236 9509 10300
rect 9443 10235 9509 10236
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 9446 6629 9506 10235
rect 9443 6628 9509 6629
rect 9443 6564 9444 6628
rect 9508 6564 9509 6628
rect 9443 6563 9509 6564
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 9630 3909 9690 11187
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 9995 9348 10061 9349
rect 9995 9284 9996 9348
rect 10060 9284 10061 9348
rect 9995 9283 10061 9284
rect 9998 6085 10058 9283
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10731 8940 10797 8941
rect 10731 8876 10732 8940
rect 10796 8876 10797 8940
rect 10731 8875 10797 8876
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 9995 6084 10061 6085
rect 9995 6020 9996 6084
rect 10060 6020 10061 6084
rect 9995 6019 10061 6020
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 9627 3908 9693 3909
rect 9627 3844 9628 3908
rect 9692 3844 9693 3908
rect 9627 3843 9693 3844
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 3926 1733 3986 2262
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 3923 1732 3989 1733
rect 3923 1668 3924 1732
rect 3988 1668 3989 1732
rect 3923 1667 3989 1668
rect 10734 1189 10794 8875
rect 13310 6901 13370 12139
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 21403 19956 21469 19957
rect 21403 19892 21404 19956
rect 21468 19892 21469 19956
rect 21403 19891 21469 19892
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 21406 15061 21466 19891
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 21403 15060 21469 15061
rect 21403 14996 21404 15060
rect 21468 14996 21469 15060
rect 21403 14995 21469 14996
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 15699 9348 15765 9349
rect 15699 9284 15700 9348
rect 15764 9284 15765 9348
rect 15699 9283 15765 9284
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 13491 7444 13557 7445
rect 13491 7380 13492 7444
rect 13556 7380 13557 7444
rect 13491 7379 13557 7380
rect 13307 6900 13373 6901
rect 13307 6836 13308 6900
rect 13372 6836 13373 6900
rect 13307 6835 13373 6836
rect 13310 5541 13370 6835
rect 13307 5540 13373 5541
rect 13307 5476 13308 5540
rect 13372 5476 13373 5540
rect 13307 5475 13373 5476
rect 13494 3365 13554 7379
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 13491 3364 13557 3365
rect 13491 3300 13492 3364
rect 13556 3300 13557 3364
rect 13491 3299 13557 3300
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 15702 2498 15762 9283
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 21406 9213 21466 14995
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 21403 9212 21469 9213
rect 21403 9148 21404 9212
rect 21468 9148 21469 9212
rect 21403 9147 21469 9148
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 2128 19930 2688
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 10731 1188 10797 1189
rect 10731 1124 10732 1188
rect 10796 1124 10797 1188
rect 10731 1123 10797 1124
<< via4 >>
rect 3838 2262 4074 2498
rect 15614 2262 15850 2498
<< metal5 >>
rect 3796 2498 15892 2540
rect 3796 2262 3838 2498
rect 4074 2262 15614 2498
rect 15850 2262 15892 2498
rect 3796 2220 15892 2262
use sky130_fd_sc_hd__fill_2  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3
timestamp 1604666999
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604666999
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1840 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17
timestamp 1604666999
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1564 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_24 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3312 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604666999
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21
timestamp 1604666999
transform 1 0 3036 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_30
timestamp 1604666999
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 1604666999
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4232 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 4324 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 6532 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1604666999
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58
timestamp 1604666999
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604666999
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604666999
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp 1604666999
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1604666999
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604666999
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604666999
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604666999
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_79
timestamp 1604666999
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_75
timestamp 1604666999
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_71
timestamp 1604666999
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 7176 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 8740 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604666999
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604666999
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604666999
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604666999
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_102
timestamp 1604666999
transform 1 0 10488 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1604666999
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_107
timestamp 1604666999
transform 1 0 10948 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_107
timestamp 1604666999
transform 1 0 10948 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1604666999
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _127_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1604666999
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604666999
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604666999
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604666999
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604666999
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604666999
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604666999
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_136
timestamp 1604666999
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1604666999
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12604 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1604666999
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_140
timestamp 1604666999
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148
timestamp 1604666999
transform 1 0 14720 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_144
timestamp 1604666999
transform 1 0 14352 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_39.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604666999
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_39.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_39.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604666999
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_39.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 14720 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_39.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 15456 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_37.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_39.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_39.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1604666999
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_167
timestamp 1604666999
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_171
timestamp 1604666999
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_175
timestamp 1604666999
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_179
timestamp 1604666999
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1604666999
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_179
timestamp 1604666999
transform 1 0 17572 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_37.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_37.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_37.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604666999
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604666999
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_37.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18308 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_37.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18032 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_207
timestamp 1604666999
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_203
timestamp 1604666999
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1604666999
transform 1 0 20056 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_35.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1604666999
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_210
timestamp 1604666999
transform 1 0 20424 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_35.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_35.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_35.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604666999
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_35.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 21160 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_35.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 20516 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_35.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1604666999
transform 1 0 22908 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_230
timestamp 1604666999
transform 1 0 22264 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_234
timestamp 1604666999
transform 1 0 22632 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_245
timestamp 1604666999
transform 1 0 23644 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_240
timestamp 1604666999
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_244
timestamp 1604666999
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_241
timestamp 1604666999
transform 1 0 23276 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604666999
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_249
timestamp 1604666999
transform 1 0 24012 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 23920 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604666999
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1604666999
transform 1 0 24196 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 24104 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604666999
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604666999
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_35.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 26036 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_260
timestamp 1604666999
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_264 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 25392 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_276
timestamp 1604666999
transform 1 0 26496 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_269
timestamp 1604666999
transform 1 0 25852 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_273
timestamp 1604666999
transform 1 0 26220 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604666999
transform 1 0 2024 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604666999
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1604666999
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_7
timestamp 1604666999
transform 1 0 1748 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_19
timestamp 1604666999
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4048 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604666999
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 3036 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604666999
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604666999
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604666999
transform 1 0 6532 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 6348 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_51
timestamp 1604666999
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_55
timestamp 1604666999
transform 1 0 6164 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7912 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_68
timestamp 1604666999
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_72
timestamp 1604666999
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_76
timestamp 1604666999
transform 1 0 8096 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 8556 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1604666999
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604666999
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1604666999
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1604666999
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1604666999
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_97
timestamp 1604666999
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 10764 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1604666999
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1604666999
transform 1 0 13248 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_124
timestamp 1604666999
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_128
timestamp 1604666999
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_39.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604666999
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_39.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_39.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14260 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1604666999
transform 1 0 14076 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_145
timestamp 1604666999
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1604666999
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604666999
transform 1 0 16836 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 17388 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1604666999
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_167
timestamp 1604666999
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_175
timestamp 1604666999
transform 1 0 17204 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_37.mux_l2_in_0_
timestamp 1604666999
transform 1 0 18032 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_37.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_37.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_179
timestamp 1604666999
transform 1 0 17572 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_193
timestamp 1604666999
transform 1 0 18860 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1604666999
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604666999
transform 1 0 19688 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_35.mux_l2_in_0_
timestamp 1604666999
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604666999
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604666999
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_31.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_201
timestamp 1604666999
transform 1 0 19596 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_206
timestamp 1604666999
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_210
timestamp 1604666999
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604666999
transform 1 0 22448 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_35.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604666999
transform 1 0 23000 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604666999
transform 1 0 22264 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_224
timestamp 1604666999
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_228
timestamp 1604666999
transform 1 0 22080 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_236
timestamp 1604666999
transform 1 0 22816 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 23552 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 23368 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_240
timestamp 1604666999
transform 1 0 23184 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604666999
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604666999
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604666999
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604666999
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 2024 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604666999
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1604666999
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1604666999
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_29
timestamp 1604666999
transform 1 0 3772 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_34
timestamp 1604666999
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_38
timestamp 1604666999
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_42
timestamp 1604666999
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_53
timestamp 1604666999
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1604666999
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604666999
transform 1 0 8372 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1604666999
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604666999
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_71
timestamp 1604666999
transform 1 0 7636 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_76
timestamp 1604666999
transform 1 0 8096 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604666999
transform 1 0 9936 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_88
timestamp 1604666999
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1604666999
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11500 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_105
timestamp 1604666999
transform 1 0 10764 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_111
timestamp 1604666999
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1604666999
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_119
timestamp 1604666999
transform 1 0 12052 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13064 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604666999
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604666999
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1604666999
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_127
timestamp 1604666999
transform 1 0 12788 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_39.mux_l1_in_0_
timestamp 1604666999
transform 1 0 14628 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_39.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_139
timestamp 1604666999
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_143
timestamp 1604666999
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_156
timestamp 1604666999
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604666999
transform 1 0 16192 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_160
timestamp 1604666999
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_173
timestamp 1604666999
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_177
timestamp 1604666999
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_37.mux_l1_in_0_
timestamp 1604666999
transform 1 0 18216 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604666999
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_37.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 1604666999
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_195
timestamp 1604666999
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_35.mux_l1_in_0_
timestamp 1604666999
transform 1 0 20700 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_35.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_35.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_35.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_199
timestamp 1604666999
transform 1 0 19412 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_205
timestamp 1604666999
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_209
timestamp 1604666999
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604666999
transform 1 0 22448 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_31.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_31.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_31.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 22080 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1604666999
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_226
timestamp 1604666999
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_230
timestamp 1604666999
transform 1 0 22264 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_236
timestamp 1604666999
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1604666999
transform 1 0 24104 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604666999
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 23920 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_31.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_240
timestamp 1604666999
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_245
timestamp 1604666999
transform 1 0 23644 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604666999
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 25116 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 25484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604666999
transform 1 0 25852 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_259
timestamp 1604666999
transform 1 0 24932 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_263
timestamp 1604666999
transform 1 0 25300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_267
timestamp 1604666999
transform 1 0 25668 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_271 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 26036 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2024 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604666999
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1604666999
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_7
timestamp 1604666999
transform 1 0 1748 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_19
timestamp 1604666999
transform 1 0 2852 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1604666999
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1604666999
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604666999
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1604666999
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_36
timestamp 1604666999
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1604666999
transform 1 0 4784 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1604666999
transform 1 0 6348 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_49
timestamp 1604666999
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_53
timestamp 1604666999
transform 1 0 5980 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1604666999
transform 1 0 7912 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7728 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1604666999
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_70
timestamp 1604666999
transform 1 0 7544 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1604666999
transform 1 0 10028 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604666999
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9292 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_83
timestamp 1604666999
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_87
timestamp 1604666999
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1604666999
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1604666999
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 11132 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 10580 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 10948 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_101
timestamp 1604666999
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_105
timestamp 1604666999
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_37.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_128
timestamp 1604666999
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_132
timestamp 1604666999
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604666999
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_39.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1604666999
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1604666999
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1604666999
transform 1 0 16836 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_163
timestamp 1604666999
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_167
timestamp 1604666999
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1604666999
transform 1 0 19136 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_37.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 18952 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_37.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 18584 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_180
timestamp 1604666999
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_184
timestamp 1604666999
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_188
timestamp 1604666999
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_192
timestamp 1604666999
transform 1 0 18768 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_31.mux_l2_in_0_
timestamp 1604666999
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604666999
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 20516 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 20148 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_205
timestamp 1604666999
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_209
timestamp 1604666999
transform 1 0 20332 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1604666999
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_31.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 22448 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_31.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_224
timestamp 1604666999
transform 1 0 21712 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_230
timestamp 1604666999
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 24380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 24748 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_251
timestamp 1604666999
transform 1 0 24196 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_255
timestamp 1604666999
transform 1 0 24564 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604666999
transform 1 0 24932 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604666999
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604666999
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1604666999
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604666999
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1604666999
transform 1 0 1380 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604666999
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_12
timestamp 1604666999
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_16
timestamp 1604666999
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604666999
transform 1 0 3220 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 4232 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 3680 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_20
timestamp 1604666999
transform 1 0 2944 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_26
timestamp 1604666999
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_30
timestamp 1604666999
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1604666999
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604666999
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 6808 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604666999
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9292 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_81
timestamp 1604666999
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_85
timestamp 1604666999
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_39.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_108
timestamp 1604666999
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_112
timestamp 1604666999
transform 1 0 11408 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604666999
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1604666999
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604666999
transform 1 0 13524 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604666999
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 1604666999
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_131
timestamp 1604666999
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 15088 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_144
timestamp 1604666999
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_148
timestamp 1604666999
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_171
timestamp 1604666999
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1604666999
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18032 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604666999
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1604666999
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1604666999
transform 1 0 20516 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_203
timestamp 1604666999
transform 1 0 19780 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_207
timestamp 1604666999
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604666999
transform 1 0 22448 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_31.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 22080 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 21528 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604666999
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_220
timestamp 1604666999
transform 1 0 21344 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_224
timestamp 1604666999
transform 1 0 21712 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_230
timestamp 1604666999
transform 1 0 22264 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_236
timestamp 1604666999
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1604666999
transform 1 0 24380 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604666999
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 24196 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 23828 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_240
timestamp 1604666999
transform 1 0 23184 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_245
timestamp 1604666999
transform 1 0 23644 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_249
timestamp 1604666999
transform 1 0 24012 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604666999
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 25392 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_262
timestamp 1604666999
transform 1 0 25208 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_266 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 25576 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_274
timestamp 1604666999
transform 1 0 26312 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_6
timestamp 1604666999
transform 1 0 1656 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_7
timestamp 1604666999
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1604666999
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604666999
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604666999
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604666999
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_16
timestamp 1604666999
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_12
timestamp 1604666999
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1604666999
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2760 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604666999
transform 1 0 2300 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_27
timestamp 1604666999
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_26
timestamp 1604666999
transform 1 0 3496 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_22
timestamp 1604666999
transform 1 0 3128 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 3312 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_31
timestamp 1604666999
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604666999
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604666999
transform 1 0 4324 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_3_
timestamp 1604666999
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_48
timestamp 1604666999
transform 1 0 5520 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_44
timestamp 1604666999
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_45
timestamp 1604666999
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_41
timestamp 1604666999
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 5336 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_2_
timestamp 1604666999
transform 1 0 5612 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1604666999
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1604666999
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1604666999
transform 1 0 6440 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_69
timestamp 1604666999
transform 1 0 7452 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_65
timestamp 1604666999
transform 1 0 7084 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_68
timestamp 1604666999
transform 1 0 7360 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_64
timestamp 1604666999
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604666999
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604666999
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_72
timestamp 1604666999
transform 1 0 7728 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_72
timestamp 1604666999
transform 1 0 7728 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 8096 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604666999
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604666999
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9292 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_84
timestamp 1604666999
transform 1 0 8832 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_88
timestamp 1604666999
transform 1 0 9200 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1604666999
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_95
timestamp 1604666999
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_99
timestamp 1604666999
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_107
timestamp 1604666999
transform 1 0 10948 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_102
timestamp 1604666999
transform 1 0 10488 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1604666999
transform 1 0 10580 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_116
timestamp 1604666999
transform 1 0 11776 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_112
timestamp 1604666999
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_118
timestamp 1604666999
transform 1 0 11960 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_112
timestamp 1604666999
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1604666999
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1604666999
transform 1 0 11592 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1604666999
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_125
timestamp 1604666999
transform 1 0 12604 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_122
timestamp 1604666999
transform 1 0 12328 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1604666999
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1604666999
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604666999
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1604666999
transform 1 0 12604 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_135
timestamp 1604666999
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_129
timestamp 1604666999
transform 1 0 12972 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 13340 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 13708 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12696 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _126_
timestamp 1604666999
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604666999
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1604666999
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_145
timestamp 1604666999
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_149
timestamp 1604666999
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_158
timestamp 1604666999
transform 1 0 15640 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_156
timestamp 1604666999
transform 1 0 15456 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_162
timestamp 1604666999
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_168
timestamp 1604666999
transform 1 0 16560 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_164
timestamp 1604666999
transform 1 0 16192 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 16008 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16376 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1604666999
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 16744 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_7_184
timestamp 1604666999
transform 1 0 18032 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604666999
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604666999
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604666999
transform 1 0 18124 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1604666999
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_189
timestamp 1604666999
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_193
timestamp 1604666999
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_189
timestamp 1604666999
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 18676 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_1_
timestamp 1604666999
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 19228 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604666999
transform 1 0 20976 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604666999
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1604666999
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_206
timestamp 1604666999
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_210
timestamp 1604666999
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_215
timestamp 1604666999
transform 1 0 20884 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_216
timestamp 1604666999
transform 1 0 20976 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_223
timestamp 1604666999
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_220
timestamp 1604666999
transform 1 0 21344 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_224
timestamp 1604666999
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_220
timestamp 1604666999
transform 1 0 21344 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604666999
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 21528 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_31.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_31.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_31.mux_l1_in_0_
timestamp 1604666999
transform 1 0 21988 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_236
timestamp 1604666999
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_31.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 22080 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_7_245
timestamp 1604666999
transform 1 0 23644 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_240
timestamp 1604666999
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_247
timestamp 1604666999
transform 1 0 23828 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604666999
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_251
timestamp 1604666999
transform 1 0 24196 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 24012 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 24380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 23920 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1604666999
transform 1 0 24564 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 24104 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604666999
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604666999
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604666999
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_264
timestamp 1604666999
transform 1 0 25392 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_272
timestamp 1604666999
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604666999
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1604666999
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_39.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604666999
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604666999
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_6
timestamp 1604666999
transform 1 0 1656 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_10
timestamp 1604666999
transform 1 0 2024 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_13
timestamp 1604666999
transform 1 0 2300 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604666999
transform 1 0 4324 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604666999
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_23
timestamp 1604666999
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1604666999
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_32
timestamp 1604666999
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604666999
transform 1 0 5888 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_44
timestamp 1604666999
transform 1 0 5152 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_50
timestamp 1604666999
transform 1 0 5704 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 7820 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_61
timestamp 1604666999
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_65
timestamp 1604666999
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_69
timestamp 1604666999
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1604666999
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_86
timestamp 1604666999
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1604666999
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_93
timestamp 1604666999
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604666999
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1604666999
transform 1 0 9752 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_97
timestamp 1604666999
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1604666999
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 10764 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 10580 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_101
timestamp 1604666999
transform 1 0 10396 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604666999
transform 1 0 13340 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_124
timestamp 1604666999
transform 1 0 12512 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_129
timestamp 1604666999
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604666999
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 14720 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_142
timestamp 1604666999
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_146
timestamp 1604666999
transform 1 0 14536 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp 1604666999
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_154
timestamp 1604666999
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_158
timestamp 1604666999
transform 1 0 15640 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 16008 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18492 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_181
timestamp 1604666999
transform 1 0 17756 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_186
timestamp 1604666999
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_198
timestamp 1604666999
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 20884 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604666999
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 19504 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_202
timestamp 1604666999
transform 1 0 19688 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp 1604666999
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_210
timestamp 1604666999
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_31.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 22816 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_234
timestamp 1604666999
transform 1 0 22632 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_238
timestamp 1604666999
transform 1 0 23000 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 23736 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 23552 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604666999
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604666999
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_265
timestamp 1604666999
transform 1 0 25484 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_273
timestamp 1604666999
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604666999
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 2116 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604666999
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1604666999
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_7
timestamp 1604666999
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1604666999
transform 1 0 3864 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_34
timestamp 1604666999
transform 1 0 4232 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_37
timestamp 1604666999
transform 1 0 4508 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_41
timestamp 1604666999
transform 1 0 4876 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1604666999
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604666999
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 6808 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604666999
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604666999
transform 1 0 9752 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_81
timestamp 1604666999
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_85
timestamp 1604666999
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_89
timestamp 1604666999
transform 1 0 9292 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_97
timestamp 1604666999
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1604666999
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604666999
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604666999
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1604666999
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604666999
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1604666999
transform 1 0 12788 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_134
timestamp 1604666999
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_130
timestamp 1604666999
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13800 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_9_157
timestamp 1604666999
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16284 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_161
timestamp 1604666999
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_174
timestamp 1604666999
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_178
timestamp 1604666999
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604666999
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_193
timestamp 1604666999
transform 1 0 18860 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604666999
transform 1 0 19596 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604666999
transform 1 0 20700 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 20516 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 20148 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_199
timestamp 1604666999
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_205
timestamp 1604666999
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_209
timestamp 1604666999
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604666999
transform 1 0 22264 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 21712 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 22080 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1604666999
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_226
timestamp 1604666999
transform 1 0 21896 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_234
timestamp 1604666999
transform 1 0 22632 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1604666999
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604666999
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_240
timestamp 1604666999
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_254
timestamp 1604666999
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604666999
transform 1 0 25208 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604666999
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604666999
transform 1 0 25760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_258
timestamp 1604666999
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_266
timestamp 1604666999
transform 1 0 25576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_270
timestamp 1604666999
transform 1 0 25944 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_276
timestamp 1604666999
transform 1 0 26496 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604666999
transform 1 0 2300 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604666999
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 2116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_39.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1604666999
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1604666999
transform 1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_22
timestamp 1604666999
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1604666999
transform 1 0 3496 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 3680 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1604666999
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604666999
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604666999
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_39
timestamp 1604666999
transform 1 0 4692 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_35
timestamp 1604666999
transform 1 0 4324 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 4508 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 5520 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_43
timestamp 1604666999
transform 1 0 5060 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_46
timestamp 1604666999
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604666999
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_67
timestamp 1604666999
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_71
timestamp 1604666999
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604666999
transform 1 0 10120 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604666999
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 9936 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1604666999
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_88
timestamp 1604666999
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_93
timestamp 1604666999
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1604666999
transform 1 0 11684 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1604666999
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_107
timestamp 1604666999
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_111
timestamp 1604666999
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l3_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_124
timestamp 1604666999
transform 1 0 12512 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_128
timestamp 1604666999
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_132
timestamp 1604666999
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604666999
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 15456 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_145
timestamp 1604666999
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_149
timestamp 1604666999
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_154
timestamp 1604666999
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_158
timestamp 1604666999
transform 1 0 15640 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16100 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 17112 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 17480 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_172
timestamp 1604666999
transform 1 0 16928 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_176
timestamp 1604666999
transform 1 0 17296 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604666999
transform 1 0 19228 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1604666999
transform 1 0 17664 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_189
timestamp 1604666999
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_193
timestamp 1604666999
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 20884 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604666999
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1604666999
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_206
timestamp 1604666999
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_210
timestamp 1604666999
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604666999
transform 1 0 22816 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_234
timestamp 1604666999
transform 1 0 22632 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_238
timestamp 1604666999
transform 1 0 23000 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 23920 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 23736 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604666999
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604666999
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_267
timestamp 1604666999
transform 1 0 25668 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604666999
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 2208 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604666999
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1604666999
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_8
timestamp 1604666999
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_31
timestamp 1604666999
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_35
timestamp 1604666999
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_39
timestamp 1604666999
transform 1 0 4692 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604666999
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1604666999
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604666999
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604666999
transform 1 0 7176 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604666999
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1604666999
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_75
timestamp 1604666999
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_79
timestamp 1604666999
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 8740 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604666999
transform 1 0 11224 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_102
timestamp 1604666999
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_106
timestamp 1604666999
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp 1604666999
transform 1 0 11500 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1604666999
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12420 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604666999
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 14996 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 14812 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14444 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_142
timestamp 1604666999
transform 1 0 14168 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_147
timestamp 1604666999
transform 1 0 14628 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_170
timestamp 1604666999
transform 1 0 16744 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp 1604666999
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18032 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604666999
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1604666999
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 20608 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 20056 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_203
timestamp 1604666999
transform 1 0 19780 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_208
timestamp 1604666999
transform 1 0 20240 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 22540 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_231
timestamp 1604666999
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_235
timestamp 1604666999
transform 1 0 22724 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1604666999
transform 1 0 23828 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604666999
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_240
timestamp 1604666999
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_245
timestamp 1604666999
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_256
timestamp 1604666999
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604666999
transform 1 0 25392 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604666999
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604666999
transform 1 0 25944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 25208 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_260
timestamp 1604666999
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_268
timestamp 1604666999
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_272
timestamp 1604666999
transform 1 0 26128 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_276
timestamp 1604666999
transform 1 0 26496 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604666999
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604666999
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_6
timestamp 1604666999
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_10
timestamp 1604666999
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4048 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604666999
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1604666999
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1604666999
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_51
timestamp 1604666999
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_55
timestamp 1604666999
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_59
timestamp 1604666999
transform 1 0 6532 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604666999
transform 1 0 7176 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_63
timestamp 1604666999
transform 1 0 6900 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_75
timestamp 1604666999
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_79
timestamp 1604666999
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_87
timestamp 1604666999
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_83
timestamp 1604666999
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9292 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_97
timestamp 1604666999
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1604666999
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1604666999
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604666999
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 10212 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_12_118
timestamp 1604666999
transform 1 0 11960 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 12696 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_122
timestamp 1604666999
transform 1 0 12328 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_125
timestamp 1604666999
transform 1 0 12604 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 15272 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604666999
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_145
timestamp 1604666999
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_149
timestamp 1604666999
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 17480 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_173
timestamp 1604666999
transform 1 0 17020 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_177
timestamp 1604666999
transform 1 0 17388 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1604666999
transform 1 0 18032 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_180
timestamp 1604666999
transform 1 0 17664 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_193
timestamp 1604666999
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1604666999
transform 1 0 19228 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1604666999
transform 1 0 19688 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604666999
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604666999
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1604666999
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 19412 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_201
timestamp 1604666999
transform 1 0 19596 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_206
timestamp 1604666999
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_210
timestamp 1604666999
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604666999
transform 1 0 22724 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 21988 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_224
timestamp 1604666999
transform 1 0 21712 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_229
timestamp 1604666999
transform 1 0 22172 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_12_238
timestamp 1604666999
transform 1 0 23000 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 23736 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 23276 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_243
timestamp 1604666999
transform 1 0 23460 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604666999
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604666999
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_265
timestamp 1604666999
transform 1 0 25484 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_273
timestamp 1604666999
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604666999
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_6
timestamp 1604666999
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_7
timestamp 1604666999
transform 1 0 1748 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604666999
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604666999
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604666999
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_10
timestamp 1604666999
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_14
timestamp 1604666999
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_11
timestamp 1604666999
transform 1 0 2116 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 2760 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1604666999
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604666999
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_27
timestamp 1604666999
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604666999
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_32
timestamp 1604666999
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_31
timestamp 1604666999
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 4324 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 4140 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604666999
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604666999
transform 1 0 4324 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 4508 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_13_44
timestamp 1604666999
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_48
timestamp 1604666999
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_52
timestamp 1604666999
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_56
timestamp 1604666999
transform 1 0 6256 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_56
timestamp 1604666999
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 6440 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_64
timestamp 1604666999
transform 1 0 6992 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_60
timestamp 1604666999
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_69
timestamp 1604666999
transform 1 0 7452 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_65
timestamp 1604666999
transform 1 0 7084 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604666999
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604666999
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_79
timestamp 1604666999
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_72
timestamp 1604666999
transform 1 0 7728 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604666999
transform 1 0 7544 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 7912 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_83
timestamp 1604666999
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_87
timestamp 1604666999
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 9292 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_93
timestamp 1604666999
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1604666999
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_93
timestamp 1604666999
transform 1 0 9660 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604666999
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_98
timestamp 1604666999
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9936 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604666999
transform 1 0 10120 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_105
timestamp 1604666999
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_101
timestamp 1604666999
transform 1 0 10396 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10580 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10488 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604666999
transform 1 0 11132 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_118
timestamp 1604666999
transform 1 0 11960 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1604666999
transform 1 0 11684 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_111
timestamp 1604666999
transform 1 0 11316 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1604666999
transform 1 0 12052 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_125
timestamp 1604666999
transform 1 0 12604 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_122
timestamp 1604666999
transform 1 0 12328 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604666999
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604666999
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12696 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_135
timestamp 1604666999
transform 1 0 13524 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_136
timestamp 1604666999
transform 1 0 13616 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1604666999
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_147
timestamp 1604666999
transform 1 0 14628 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_143
timestamp 1604666999
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_139
timestamp 1604666999
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_141
timestamp 1604666999
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_1_
timestamp 1604666999
transform 1 0 14444 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_158
timestamp 1604666999
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_154
timestamp 1604666999
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604666999
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_167
timestamp 1604666999
transform 1 0 16468 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_163
timestamp 1604666999
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1604666999
transform 1 0 16008 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_177
timestamp 1604666999
transform 1 0 17388 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_171
timestamp 1604666999
transform 1 0 16836 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1604666999
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_171
timestamp 1604666999
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1604666999
transform 1 0 17112 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18032 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18124 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604666999
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 17940 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 17572 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1604666999
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_181
timestamp 1604666999
transform 1 0 17756 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_194
timestamp 1604666999
transform 1 0 18952 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_206
timestamp 1604666999
transform 1 0 20056 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_202
timestamp 1604666999
transform 1 0 19688 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_207
timestamp 1604666999
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_203
timestamp 1604666999
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 19780 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604666999
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_210
timestamp 1604666999
transform 1 0 20424 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_215
timestamp 1604666999
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1604666999
transform 1 0 20516 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 20332 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604666999
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_1_
timestamp 1604666999
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604666999
transform 1 0 20516 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_224
timestamp 1604666999
transform 1 0 21712 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_223
timestamp 1604666999
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_219
timestamp 1604666999
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 21988 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604666999
transform 1 0 21988 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_237
timestamp 1604666999
transform 1 0 22908 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_229
timestamp 1604666999
transform 1 0 22172 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_236
timestamp 1604666999
transform 1 0 22816 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 22724 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 23276 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604666999
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604666999
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 23276 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 23092 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_240
timestamp 1604666999
transform 1 0 23184 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 1604666999
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_254
timestamp 1604666999
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_266
timestamp 1604666999
transform 1 0 25576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_258
timestamp 1604666999
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604666999
transform 1 0 25208 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604666999
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_272
timestamp 1604666999
transform 1 0 26128 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_276
timestamp 1604666999
transform 1 0 26496 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_270
timestamp 1604666999
transform 1 0 25944 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604666999
transform 1 0 25760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604666999
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604666999
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604666999
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_260
timestamp 1604666999
transform 1 0 25024 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604666999
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 2576 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604666999
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604666999
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604666999
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_7
timestamp 1604666999
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_11
timestamp 1604666999
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_15
timestamp 1604666999
transform 1 0 2484 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_35
timestamp 1604666999
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_39
timestamp 1604666999
transform 1 0 4692 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604666999
transform 1 0 5060 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 4876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 6440 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_52
timestamp 1604666999
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_56
timestamp 1604666999
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 7544 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604666999
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1604666999
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1604666999
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_66
timestamp 1604666999
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1604666999
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_93
timestamp 1604666999
transform 1 0 9660 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_97
timestamp 1604666999
transform 1 0 10028 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10304 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_109
timestamp 1604666999
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_113
timestamp 1604666999
transform 1 0 11500 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1604666999
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604666999
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1604666999
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1604666999
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604666999
transform 1 0 14444 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 15456 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_140
timestamp 1604666999
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_144
timestamp 1604666999
transform 1 0 14352 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_148
timestamp 1604666999
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_152
timestamp 1604666999
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1604666999
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1604666999
transform 1 0 18216 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604666999
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604666999
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1604666999
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_195
timestamp 1604666999
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1604666999
transform 1 0 20608 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_199
timestamp 1604666999
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_203
timestamp 1604666999
transform 1 0 19780 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_208
timestamp 1604666999
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604666999
transform 1 0 22448 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604666999
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1604666999
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_225
timestamp 1604666999
transform 1 0 21804 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_229
timestamp 1604666999
transform 1 0 22172 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_236
timestamp 1604666999
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604666999
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604666999
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604666999
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_254
timestamp 1604666999
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604666999
transform 1 0 25208 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604666999
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604666999
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604666999
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_258
timestamp 1604666999
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_266
timestamp 1604666999
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_270
timestamp 1604666999
transform 1 0 25944 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_276
timestamp 1604666999
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604666999
transform 1 0 2484 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604666999
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604666999
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_7
timestamp 1604666999
transform 1 0 1748 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_11
timestamp 1604666999
transform 1 0 2116 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_14
timestamp 1604666999
transform 1 0 2392 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_19
timestamp 1604666999
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604666999
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604666999
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604666999
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604666999
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1604666999
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604666999
transform 1 0 5612 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 1604666999
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_45
timestamp 1604666999
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_58
timestamp 1604666999
transform 1 0 6440 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1604666999
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_62
timestamp 1604666999
transform 1 0 6808 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_65
timestamp 1604666999
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_69
timestamp 1604666999
transform 1 0 7452 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_74
timestamp 1604666999
transform 1 0 7912 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604666999
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604666999
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 10120 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_84
timestamp 1604666999
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_88
timestamp 1604666999
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_96
timestamp 1604666999
transform 1 0 9936 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 10672 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_100
timestamp 1604666999
transform 1 0 10304 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604666999
transform 1 0 13156 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_123
timestamp 1604666999
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_127
timestamp 1604666999
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 15272 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604666999
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_140
timestamp 1604666999
transform 1 0 13984 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_144
timestamp 1604666999
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_148
timestamp 1604666999
transform 1 0 14720 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 17204 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_173
timestamp 1604666999
transform 1 0 17020 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_177
timestamp 1604666999
transform 1 0 17388 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18032 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 17848 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_181
timestamp 1604666999
transform 1 0 17756 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 20884 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604666999
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_203
timestamp 1604666999
transform 1 0 19780 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_207
timestamp 1604666999
transform 1 0 20148 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_210
timestamp 1604666999
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 22908 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_234
timestamp 1604666999
transform 1 0 22632 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604666999
transform 1 0 23460 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604666999
transform 1 0 24564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 23276 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_239
timestamp 1604666999
transform 1 0 23092 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_252
timestamp 1604666999
transform 1 0 24288 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_257
timestamp 1604666999
transform 1 0 24748 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604666999
transform 1 0 25024 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604666999
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604666999
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_264
timestamp 1604666999
transform 1 0 25392 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_272
timestamp 1604666999
transform 1 0 26128 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604666999
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604666999
transform 1 0 2208 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604666999
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 1656 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1604666999
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_8
timestamp 1604666999
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 3772 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_21
timestamp 1604666999
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_25
timestamp 1604666999
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_48
timestamp 1604666999
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_52
timestamp 1604666999
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_56
timestamp 1604666999
transform 1 0 6256 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 7268 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604666999
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1604666999
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_62
timestamp 1604666999
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1604666999
transform 1 0 9752 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_86
timestamp 1604666999
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_90
timestamp 1604666999
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604666999
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_103
timestamp 1604666999
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_107
timestamp 1604666999
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1604666999
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604666999
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604666999
transform 1 0 12604 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 13616 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604666999
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1604666999
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_128
timestamp 1604666999
transform 1 0 12880 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_133
timestamp 1604666999
transform 1 0 13340 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1604666999
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604666999
transform 1 0 16100 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_159
timestamp 1604666999
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_172
timestamp 1604666999
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_176
timestamp 1604666999
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1604666999
transform 1 0 18124 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 19320 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604666999
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 19136 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 18768 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1604666999
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_184
timestamp 1604666999
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_188
timestamp 1604666999
transform 1 0 18400 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_194
timestamp 1604666999
transform 1 0 18952 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1604666999
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1604666999
transform 1 0 21804 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1604666999
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_234
timestamp 1604666999
transform 1 0 22632 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_238
timestamp 1604666999
transform 1 0 23000 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 23644 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604666999
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604666999
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_264
timestamp 1604666999
transform 1 0 25392 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_276
timestamp 1604666999
transform 1 0 26496 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1604666999
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604666999
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_6
timestamp 1604666999
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_10
timestamp 1604666999
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604666999
transform 1 0 4232 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604666999
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 4692 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604666999
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604666999
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1604666999
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_37
timestamp 1604666999
transform 1 0 4508 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1604666999
transform 1 0 5244 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1604666999
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_54
timestamp 1604666999
transform 1 0 6072 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_58
timestamp 1604666999
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604666999
transform 1 0 7728 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_62
timestamp 1604666999
transform 1 0 6808 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_67
timestamp 1604666999
transform 1 0 7268 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_81
timestamp 1604666999
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp 1604666999
transform 1 0 9292 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1604666999
transform 1 0 8924 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1604666999
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604666999
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_97
timestamp 1604666999
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 10212 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 10396 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13156 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_120
timestamp 1604666999
transform 1 0 12144 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_124
timestamp 1604666999
transform 1 0 12512 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_128
timestamp 1604666999
transform 1 0 12880 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_140
timestamp 1604666999
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_144
timestamp 1604666999
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_148
timestamp 1604666999
transform 1 0 14720 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14904 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1604666999
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604666999
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604666999
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_157
timestamp 1604666999
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 16560 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 15732 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_161
timestamp 1604666999
transform 1 0 15916 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_165
timestamp 1604666999
transform 1 0 16284 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604666999
transform 1 0 19044 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_187
timestamp 1604666999
transform 1 0 18308 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_191
timestamp 1604666999
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1604666999
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604666999
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_204
timestamp 1604666999
transform 1 0 19872 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_208
timestamp 1604666999
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1604666999
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_218
timestamp 1604666999
transform 1 0 21160 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 21988 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 21804 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 21436 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_223
timestamp 1604666999
transform 1 0 21620 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604666999
transform 1 0 24564 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 23920 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_246
timestamp 1604666999
transform 1 0 23736 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_250
timestamp 1604666999
transform 1 0 24104 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_254
timestamp 1604666999
transform 1 0 24472 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604666999
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604666999
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_259
timestamp 1604666999
transform 1 0 24932 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_271
timestamp 1604666999
transform 1 0 26036 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604666999
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604666999
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604666999
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604666999
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604666999
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_7
timestamp 1604666999
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1604666999
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604666999
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604666999
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1604666999
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1604666999
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 2300 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_19
timestamp 1604666999
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_15
timestamp 1604666999
transform 1 0 2484 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604666999
transform 1 0 2484 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1604666999
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1604666999
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604666999
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604666999
transform 1 0 3036 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1604666999
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_34
timestamp 1604666999
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_30
timestamp 1604666999
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604666999
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604666999
transform 1 0 4600 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 4232 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_47
timestamp 1604666999
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604666999
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_53
timestamp 1604666999
transform 1 0 5980 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_68
timestamp 1604666999
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_64
timestamp 1604666999
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_61
timestamp 1604666999
transform 1 0 6716 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_68
timestamp 1604666999
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_62
timestamp 1604666999
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604666999
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 7084 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_79
timestamp 1604666999
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_72
timestamp 1604666999
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1604666999
transform 1 0 7544 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1604666999
transform 1 0 8096 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_89
timestamp 1604666999
transform 1 0 9292 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_83
timestamp 1604666999
transform 1 0 8740 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_89
timestamp 1604666999
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_85
timestamp 1604666999
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604666999
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604666999
transform 1 0 9660 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_106
timestamp 1604666999
transform 1 0 10856 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1604666999
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_106
timestamp 1604666999
transform 1 0 10856 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_102
timestamp 1604666999
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_113
timestamp 1604666999
transform 1 0 11500 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_110
timestamp 1604666999
transform 1 0 11224 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_114
timestamp 1604666999
transform 1 0 11592 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 11684 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 11316 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604666999
transform 1 0 11868 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_119
timestamp 1604666999
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_126
timestamp 1604666999
transform 1 0 12696 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1604666999
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1604666999
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604666999
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 12604 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_132
timestamp 1604666999
transform 1 0 13248 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1604666999
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 13064 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13524 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604666999
transform 1 0 13616 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_148
timestamp 1604666999
transform 1 0 14720 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_144
timestamp 1604666999
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_145
timestamp 1604666999
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_158
timestamp 1604666999
transform 1 0 15640 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1604666999
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_149
timestamp 1604666999
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604666999
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604666999
transform 1 0 15180 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 16008 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16744 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 15824 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_162
timestamp 1604666999
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1604666999
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_173
timestamp 1604666999
transform 1 0 17020 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_186
timestamp 1604666999
transform 1 0 18216 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_181
timestamp 1604666999
transform 1 0 17756 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604666999
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604666999
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_198
timestamp 1604666999
transform 1 0 19320 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_197
timestamp 1604666999
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_193
timestamp 1604666999
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604666999
transform 1 0 18492 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_207
timestamp 1604666999
transform 1 0 20148 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_203
timestamp 1604666999
transform 1 0 19780 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 19964 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 19596 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1604666999
transform 1 0 19596 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1604666999
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_214
timestamp 1604666999
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_210
timestamp 1604666999
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 20976 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604666999
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1604666999
transform 1 0 21160 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604666999
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_218
timestamp 1604666999
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1604666999
transform 1 0 22540 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 22540 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_221
timestamp 1604666999
transform 1 0 21436 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1604666999
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_230
timestamp 1604666999
transform 1 0 22264 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_236
timestamp 1604666999
transform 1 0 22816 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_245
timestamp 1604666999
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_240
timestamp 1604666999
transform 1 0 23184 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604666999
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 23552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_247
timestamp 1604666999
transform 1 0 23828 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_249
timestamp 1604666999
transform 1 0 24012 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23828 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604666999
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604666999
transform 1 0 24564 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604666999
transform 1 0 24564 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_259
timestamp 1604666999
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604666999
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604666999
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_271
timestamp 1604666999
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_275
timestamp 1604666999
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604666999
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604666999
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604666999
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_259
timestamp 1604666999
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_263
timestamp 1604666999
transform 1 0 25300 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604666999
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 2484 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604666999
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604666999
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604666999
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_7
timestamp 1604666999
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1604666999
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_18
timestamp 1604666999
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 4232 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_22
timestamp 1604666999
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_26
timestamp 1604666999
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_30
timestamp 1604666999
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1604666999
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604666999
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 7176 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604666999
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1604666999
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_85
timestamp 1604666999
transform 1 0 8924 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_91
timestamp 1604666999
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_95
timestamp 1604666999
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_99
timestamp 1604666999
transform 1 0 10212 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10488 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_111
timestamp 1604666999
transform 1 0 11316 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_115
timestamp 1604666999
transform 1 0 11684 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604666999
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 13064 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604666999
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1604666999
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_127
timestamp 1604666999
transform 1 0 12788 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_149
timestamp 1604666999
transform 1 0 14812 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_153
timestamp 1604666999
transform 1 0 15180 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_156
timestamp 1604666999
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604666999
transform 1 0 16100 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 17480 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_160
timestamp 1604666999
transform 1 0 15824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_172
timestamp 1604666999
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_176
timestamp 1604666999
transform 1 0 17296 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604666999
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604666999
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_180
timestamp 1604666999
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_193
timestamp 1604666999
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_197
timestamp 1604666999
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604666999
transform 1 0 19596 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 20976 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604666999
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_204
timestamp 1604666999
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_208
timestamp 1604666999
transform 1 0 20240 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 22540 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_219
timestamp 1604666999
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_223
timestamp 1604666999
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_227
timestamp 1604666999
transform 1 0 21988 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_236
timestamp 1604666999
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604666999
transform 1 0 24564 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604666999
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23828 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604666999
transform 1 0 24380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604666999
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_245
timestamp 1604666999
transform 1 0 23644 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_249
timestamp 1604666999
transform 1 0 24012 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604666999
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604666999
transform 1 0 25116 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_259
timestamp 1604666999
transform 1 0 24932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_263
timestamp 1604666999
transform 1 0 25300 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_275
timestamp 1604666999
transform 1 0 26404 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604666999
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 2484 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604666999
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1932 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2300 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1604666999
transform 1 0 1748 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_11
timestamp 1604666999
transform 1 0 2116 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_18
timestamp 1604666999
transform 1 0 2760 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604666999
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604666999
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604666999
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604666999
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 5612 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_41
timestamp 1604666999
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_45
timestamp 1604666999
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604666999
transform 1 0 8188 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 7912 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_68
timestamp 1604666999
transform 1 0 7360 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_76
timestamp 1604666999
transform 1 0 8096 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9660 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604666999
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_80
timestamp 1604666999
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_84
timestamp 1604666999
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 11960 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_112
timestamp 1604666999
transform 1 0 11408 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1604666999
transform 1 0 11776 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604666999
transform 1 0 12144 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13616 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_129
timestamp 1604666999
transform 1 0 12972 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_133
timestamp 1604666999
transform 1 0 13340 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1604666999
transform 1 0 13800 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 14168 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604666999
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1604666999
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1604666999
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604666999
transform 1 0 16836 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_163
timestamp 1604666999
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_167
timestamp 1604666999
transform 1 0 16468 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604666999
transform 1 0 18400 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 18952 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_180
timestamp 1604666999
transform 1 0 17664 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_186
timestamp 1604666999
transform 1 0 18216 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_192
timestamp 1604666999
transform 1 0 18768 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_196
timestamp 1604666999
transform 1 0 19136 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 19504 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604666999
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_203
timestamp 1604666999
transform 1 0 19780 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_211
timestamp 1604666999
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_218
timestamp 1604666999
transform 1 0 21160 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 22540 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_230
timestamp 1604666999
transform 1 0 22264 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_236
timestamp 1604666999
transform 1 0 22816 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604666999
transform 1 0 24564 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 23552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_247
timestamp 1604666999
transform 1 0 23828 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604666999
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604666999
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_259
timestamp 1604666999
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1604666999
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604666999
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604666999
transform 1 0 1840 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604666999
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604666999
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604666999
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1604666999
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1604666999
transform 1 0 1748 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_12
timestamp 1604666999
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_16
timestamp 1604666999
transform 1 0 2576 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604666999
transform 1 0 3864 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_26
timestamp 1604666999
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604666999
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604666999
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604666999
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1604666999
transform 1 0 6900 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 7912 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604666999
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 7360 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_62
timestamp 1604666999
transform 1 0 6808 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_66
timestamp 1604666999
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_70
timestamp 1604666999
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_93
timestamp 1604666999
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_97
timestamp 1604666999
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1604666999
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1604666999
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604666999
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604666999
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604666999
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1604666999
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_136
timestamp 1604666999
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13984 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_23_159
timestamp 1604666999
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_163
timestamp 1604666999
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_170
timestamp 1604666999
transform 1 0 16744 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16468 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_174
timestamp 1604666999
transform 1 0 17112 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 16928 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_178
timestamp 1604666999
transform 1 0 17480 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604666999
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 19136 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604666999
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 18492 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 17664 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1604666999
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_187
timestamp 1604666999
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_191
timestamp 1604666999
transform 1 0 18676 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_195
timestamp 1604666999
transform 1 0 19044 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 20332 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 20792 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 19964 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_199
timestamp 1604666999
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_203
timestamp 1604666999
transform 1 0 19780 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_207
timestamp 1604666999
transform 1 0 20148 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_212
timestamp 1604666999
transform 1 0 20608 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_216
timestamp 1604666999
transform 1 0 20976 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1604666999
transform 1 0 21528 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 22540 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_225
timestamp 1604666999
transform 1 0 21804 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1604666999
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604666999
transform 1 0 24564 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604666999
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604666999
transform 1 0 24380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23828 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_240
timestamp 1604666999
transform 1 0 23184 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_245
timestamp 1604666999
transform 1 0 23644 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_249
timestamp 1604666999
transform 1 0 24012 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604666999
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604666999
transform 1 0 25116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_259
timestamp 1604666999
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_263
timestamp 1604666999
transform 1 0 25300 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_275
timestamp 1604666999
transform 1 0 26404 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604666999
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604666999
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_7
timestamp 1604666999
transform 1 0 1748 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_19
timestamp 1604666999
transform 1 0 2852 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604666999
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1604666999
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_36
timestamp 1604666999
transform 1 0 4416 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_48
timestamp 1604666999
transform 1 0 5520 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604666999
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_60
timestamp 1604666999
transform 1 0 6624 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_72
timestamp 1604666999
transform 1 0 7728 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604666999
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604666999
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_84
timestamp 1604666999
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_96
timestamp 1604666999
transform 1 0 9936 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 10672 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_123
timestamp 1604666999
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_127
timestamp 1604666999
transform 1 0 12788 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_131
timestamp 1604666999
transform 1 0 13156 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_134
timestamp 1604666999
transform 1 0 13432 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604666999
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604666999
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_145
timestamp 1604666999
transform 1 0 14444 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1604666999
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 16836 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 16652 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_163
timestamp 1604666999
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_167
timestamp 1604666999
transform 1 0 16468 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 18400 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_180
timestamp 1604666999
transform 1 0 17664 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_191
timestamp 1604666999
transform 1 0 18676 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 19412 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604666999
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1604666999
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604666999
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1604666999
transform 1 0 22540 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_227
timestamp 1604666999
transform 1 0 21988 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_236
timestamp 1604666999
transform 1 0 22816 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604666999
transform 1 0 24564 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 23552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_247
timestamp 1604666999
transform 1 0 23828 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604666999
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604666999
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_259
timestamp 1604666999
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_271
timestamp 1604666999
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604666999
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604666999
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 2484 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604666999
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604666999
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604666999
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1604666999
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1604666999
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_18
timestamp 1604666999
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_22
timestamp 1604666999
transform 1 0 3128 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_34
timestamp 1604666999
transform 1 0 4232 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_46
timestamp 1604666999
transform 1 0 5336 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_58
timestamp 1604666999
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604666999
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604666999
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_74
timestamp 1604666999
transform 1 0 7912 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_78
timestamp 1604666999
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1604666999
transform 1 0 10212 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1604666999
transform 1 0 8648 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_91
timestamp 1604666999
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_95
timestamp 1604666999
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_108
timestamp 1604666999
transform 1 0 11040 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_112
timestamp 1604666999
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_116
timestamp 1604666999
transform 1 0 11776 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 13248 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604666999
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1604666999
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_127
timestamp 1604666999
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp 1604666999
transform 1 0 13156 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 14812 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_141
timestamp 1604666999
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_145
timestamp 1604666999
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16744 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_168
timestamp 1604666999
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1604666999
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_176
timestamp 1604666999
transform 1 0 17296 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604666999
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1604666999
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_187
timestamp 1604666999
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_191
timestamp 1604666999
transform 1 0 18676 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_203
timestamp 1604666999
transform 1 0 19780 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_215
timestamp 1604666999
transform 1 0 20884 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_227
timestamp 1604666999
transform 1 0 21988 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1604666999
transform 1 0 24196 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604666999
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604666999
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23828 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_239
timestamp 1604666999
transform 1 0 23092 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_243
timestamp 1604666999
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_245
timestamp 1604666999
transform 1 0 23644 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_249
timestamp 1604666999
transform 1 0 24012 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_254
timestamp 1604666999
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604666999
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_258
timestamp 1604666999
transform 1 0 24840 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_270
timestamp 1604666999
transform 1 0 25944 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_276
timestamp 1604666999
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1604666999
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604666999
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604666999
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604666999
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604666999
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604666999
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1604666999
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604666999
transform 1 0 2300 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604666999
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_19
timestamp 1604666999
transform 1 0 2852 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_7
timestamp 1604666999
transform 1 0 1748 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604666999
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604666999
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604666999
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604666999
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604666999
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604666999
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604666999
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604666999
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604666999
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604666999
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604666999
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604666999
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_86
timestamp 1604666999
transform 1 0 9016 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_84
timestamp 1604666999
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_80
timestamp 1604666999
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_96
timestamp 1604666999
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_93
timestamp 1604666999
transform 1 0 9660 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604666999
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 10212 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 10488 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604666999
transform 1 0 10672 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_101
timestamp 1604666999
transform 1 0 10396 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_100
timestamp 1604666999
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1604666999
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_117
timestamp 1604666999
transform 1 0 11868 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_125
timestamp 1604666999
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_121
timestamp 1604666999
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604666999
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_137
timestamp 1604666999
transform 1 0 13708 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_132
timestamp 1604666999
transform 1 0 13248 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1604666999
transform 1 0 13800 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12972 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_141
timestamp 1604666999
transform 1 0 14076 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_146
timestamp 1604666999
transform 1 0 14536 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_142
timestamp 1604666999
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_150
timestamp 1604666999
transform 1 0 14904 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604666999
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 14352 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16836 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_163
timestamp 1604666999
transform 1 0 16100 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_174
timestamp 1604666999
transform 1 0 17112 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_163
timestamp 1604666999
transform 1 0 16100 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_175
timestamp 1604666999
transform 1 0 17204 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604666999
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_186
timestamp 1604666999
transform 1 0 18216 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_198
timestamp 1604666999
transform 1 0 19320 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604666999
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604666999
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604666999
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1604666999
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604666999
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604666999
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604666999
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604666999
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604666999
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604666999
transform 1 0 24564 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604666999
transform 1 0 24564 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 23552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604666999
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604666999
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_239
timestamp 1604666999
transform 1 0 23092 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_243
timestamp 1604666999
transform 1 0 23460 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_247
timestamp 1604666999
transform 1 0 23828 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_245
timestamp 1604666999
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_259
timestamp 1604666999
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604666999
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_275
timestamp 1604666999
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604666999
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1604666999
transform 1 0 26036 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604666999
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604666999
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604666999
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_263
timestamp 1604666999
transform 1 0 25300 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_259
timestamp 1604666999
transform 1 0 24932 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604666999
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604666999
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_7
timestamp 1604666999
transform 1 0 1748 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_19
timestamp 1604666999
transform 1 0 2852 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604666999
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604666999
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604666999
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604666999
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604666999
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604666999
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604666999
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_93
timestamp 1604666999
transform 1 0 9660 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 11040 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_101
timestamp 1604666999
transform 1 0 10396 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_106
timestamp 1604666999
transform 1 0 10856 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1604666999
transform 1 0 13524 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13340 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_127
timestamp 1604666999
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_131
timestamp 1604666999
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604666999
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604666999
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_144
timestamp 1604666999
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_148
timestamp 1604666999
transform 1 0 14720 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1604666999
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_157
timestamp 1604666999
transform 1 0 15548 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_169
timestamp 1604666999
transform 1 0 16652 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_181
timestamp 1604666999
transform 1 0 17756 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_193
timestamp 1604666999
transform 1 0 18860 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604666999
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_205
timestamp 1604666999
transform 1 0 19964 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1604666999
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604666999
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604666999
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604666999
transform 1 0 24564 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604666999
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_251
timestamp 1604666999
transform 1 0 24196 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604666999
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604666999
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_259
timestamp 1604666999
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1604666999
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604666999
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604666999
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604666999
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604666999
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_7
timestamp 1604666999
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1604666999
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604666999
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604666999
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604666999
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604666999
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604666999
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604666999
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604666999
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604666999
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1604666999
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1604666999
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1604666999
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604666999
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604666999
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12420 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604666999
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_142
timestamp 1604666999
transform 1 0 14168 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_154
timestamp 1604666999
transform 1 0 15272 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_166
timestamp 1604666999
transform 1 0 16376 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_178
timestamp 1604666999
transform 1 0 17480 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604666999
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1604666999
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604666999
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604666999
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604666999
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604666999
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604666999
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604666999
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1604666999
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604666999
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604666999
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1604666999
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1564 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604666999
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1604666999
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_8
timestamp 1604666999
transform 1 0 1840 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604666999
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_20
timestamp 1604666999
transform 1 0 2944 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_28
timestamp 1604666999
transform 1 0 3680 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604666999
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604666999
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604666999
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1604666999
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604666999
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604666999
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1604666999
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1604666999
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_117
timestamp 1604666999
transform 1 0 11868 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1604666999
transform 1 0 12420 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 13524 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 12236 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_132
timestamp 1604666999
transform 1 0 13248 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_137
timestamp 1604666999
transform 1 0 13708 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604666999
transform 1 0 13984 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604666999
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_143
timestamp 1604666999
transform 1 0 14260 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1604666999
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604666999
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1604666999
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1604666999
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1604666999
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604666999
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1604666999
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604666999
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604666999
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604666999
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604666999
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604666999
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604666999
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604666999
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604666999
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604666999
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604666999
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604666999
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604666999
transform 1 0 2300 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1604666999
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1604666999
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604666999
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604666999
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604666999
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604666999
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604666999
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604666999
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604666999
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604666999
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604666999
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604666999
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604666999
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 13524 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604666999
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 13340 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_123
timestamp 1604666999
transform 1 0 12420 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_131
timestamp 1604666999
transform 1 0 13156 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_154
timestamp 1604666999
transform 1 0 15272 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_166
timestamp 1604666999
transform 1 0 16376 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_178
timestamp 1604666999
transform 1 0 17480 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604666999
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1604666999
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604666999
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604666999
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604666999
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604666999
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604666999
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604666999
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604666999
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604666999
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604666999
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1604666999
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604666999
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604666999
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_7
timestamp 1604666999
transform 1 0 1748 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_19
timestamp 1604666999
transform 1 0 2852 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604666999
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604666999
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604666999
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604666999
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604666999
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604666999
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604666999
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604666999
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604666999
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604666999
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13340 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_129
timestamp 1604666999
transform 1 0 12972 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_135
timestamp 1604666999
transform 1 0 13524 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604666999
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_147
timestamp 1604666999
transform 1 0 14628 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604666999
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1604666999
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1604666999
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1604666999
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604666999
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1604666999
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604666999
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604666999
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1604666999
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1604666999
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604666999
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604666999
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1604666999
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604666999
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1604666999
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1604666999
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604666999
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604666999
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604666999
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1564 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604666999
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_11
timestamp 1604666999
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_8
timestamp 1604666999
transform 1 0 1840 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604666999
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604666999
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604666999
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604666999
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_20
timestamp 1604666999
transform 1 0 2944 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_28
timestamp 1604666999
transform 1 0 3680 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604666999
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604666999
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604666999
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604666999
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604666999
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604666999
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604666999
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1604666999
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604666999
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604666999
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1604666999
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1604666999
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604666999
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604666999
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1604666999
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604666999
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604666999
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13340 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604666999
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 13156 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_123
timestamp 1604666999
transform 1 0 12420 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604666999
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604666999
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_152
timestamp 1604666999
transform 1 0 15088 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604666999
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604666999
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_164
timestamp 1604666999
transform 1 0 16192 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_176
timestamp 1604666999
transform 1 0 17296 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604666999
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604666999
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604666999
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_182
timestamp 1604666999
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604666999
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604666999
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604666999
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604666999
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604666999
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604666999
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604666999
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604666999
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1604666999
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604666999
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604666999
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604666999
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1604666999
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604666999
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604666999
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604666999
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604666999
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604666999
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1604666999
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604666999
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604666999
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604666999
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604666999
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604666999
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1604666999
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1604666999
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1604666999
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604666999
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604666999
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604666999
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1604666999
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_86
timestamp 1604666999
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_98
timestamp 1604666999
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_110
timestamp 1604666999
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604666999
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1604666999
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_135
timestamp 1604666999
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_147
timestamp 1604666999
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_159
timestamp 1604666999
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_171
timestamp 1604666999
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604666999
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604666999
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604666999
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604666999
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604666999
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1604666999
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604666999
transform 1 0 24564 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604666999
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604666999
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23828 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_245
timestamp 1604666999
transform 1 0 23644 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_249
timestamp 1604666999
transform 1 0 24012 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604666999
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604666999
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_259
timestamp 1604666999
transform 1 0 24932 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_263
timestamp 1604666999
transform 1 0 25300 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_275
timestamp 1604666999
transform 1 0 26404 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604666999
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604666999
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604666999
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604666999
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604666999
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604666999
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1604666999
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1604666999
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1604666999
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604666999
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1604666999
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1604666999
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1604666999
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_117
timestamp 1604666999
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1604666999
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604666999
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1604666999
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1604666999
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_166
timestamp 1604666999
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_178
timestamp 1604666999
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_190
timestamp 1604666999
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604666999
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_202
timestamp 1604666999
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604666999
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604666999
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604666999
transform 1 0 24564 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 23552 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_239
timestamp 1604666999
transform 1 0 23092 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_243
timestamp 1604666999
transform 1 0 23460 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_247
timestamp 1604666999
transform 1 0 23828 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604666999
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604666999
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_259
timestamp 1604666999
transform 1 0 24932 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_271
timestamp 1604666999
transform 1 0 26036 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604666999
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604666999
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604666999
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604666999
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_7
timestamp 1604666999
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_11
timestamp 1604666999
transform 1 0 2116 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_23
timestamp 1604666999
transform 1 0 3220 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_35
timestamp 1604666999
transform 1 0 4324 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_47
timestamp 1604666999
transform 1 0 5428 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1604666999
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604666999
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1604666999
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1604666999
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1604666999
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_98
timestamp 1604666999
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_110
timestamp 1604666999
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604666999
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1604666999
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_135
timestamp 1604666999
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_147
timestamp 1604666999
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_159
timestamp 1604666999
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_171
timestamp 1604666999
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604666999
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1604666999
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1604666999
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1604666999
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_220
timestamp 1604666999
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_232
timestamp 1604666999
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604666999
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604666999
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_245
timestamp 1604666999
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_253
timestamp 1604666999
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1604666999
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604666999
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1604666999
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604666999
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604666999
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604666999
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604666999
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604666999
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604666999
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604666999
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604666999
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1604666999
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604666999
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1604666999
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1604666999
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1604666999
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_117
timestamp 1604666999
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_129
timestamp 1604666999
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604666999
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1604666999
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1604666999
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1604666999
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_178
timestamp 1604666999
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_190
timestamp 1604666999
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604666999
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_202
timestamp 1604666999
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1604666999
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1604666999
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604666999
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1604666999
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_251
timestamp 1604666999
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604666999
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604666999
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_259
timestamp 1604666999
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_271
timestamp 1604666999
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604666999
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604666999
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604666999
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604666999
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604666999
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604666999
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604666999
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604666999
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604666999
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1604666999
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604666999
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604666999
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1604666999
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1604666999
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604666999
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604666999
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604666999
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604666999
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1604666999
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1604666999
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604666999
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1604666999
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_98
timestamp 1604666999
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604666999
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604666999
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_110
timestamp 1604666999
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1604666999
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_117
timestamp 1604666999
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604666999
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1604666999
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_135
timestamp 1604666999
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1604666999
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604666999
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_147
timestamp 1604666999
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1604666999
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1604666999
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_159
timestamp 1604666999
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_171
timestamp 1604666999
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_166
timestamp 1604666999
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1604666999
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604666999
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1604666999
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1604666999
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_190
timestamp 1604666999
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604666999
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1604666999
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_202
timestamp 1604666999
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1604666999
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_220
timestamp 1604666999
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_232
timestamp 1604666999
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1604666999
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604666999
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1604666999
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_257
timestamp 1604666999
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1604666999
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_251
timestamp 1604666999
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604666999
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604666999
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604666999
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1604666999
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_263
timestamp 1604666999
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604666999
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604666999
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604666999
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604666999
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604666999
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1604666999
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1604666999
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604666999
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604666999
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604666999
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604666999
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604666999
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604666999
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1604666999
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604666999
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604666999
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1604666999
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_147
timestamp 1604666999
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_159
timestamp 1604666999
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_171
timestamp 1604666999
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604666999
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604666999
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604666999
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604666999
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604666999
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604666999
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604666999
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604666999
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604666999
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604666999
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604666999
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604666999
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604666999
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604666999
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604666999
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604666999
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604666999
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604666999
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604666999
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604666999
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604666999
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604666999
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604666999
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604666999
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604666999
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604666999
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604666999
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604666999
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604666999
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604666999
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604666999
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604666999
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604666999
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604666999
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604666999
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604666999
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604666999
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604666999
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604666999
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604666999
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604666999
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604666999
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604666999
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604666999
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604666999
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604666999
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604666999
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604666999
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_34_
port 0 nsew default input
rlabel metal2 s 846 0 902 480 6 bottom_left_grid_pin_35_
port 1 nsew default input
rlabel metal2 s 1398 0 1454 480 6 bottom_left_grid_pin_36_
port 2 nsew default input
rlabel metal2 s 2042 0 2098 480 6 bottom_left_grid_pin_37_
port 3 nsew default input
rlabel metal2 s 2594 0 2650 480 6 bottom_left_grid_pin_38_
port 4 nsew default input
rlabel metal2 s 3146 0 3202 480 6 bottom_left_grid_pin_39_
port 5 nsew default input
rlabel metal2 s 3790 0 3846 480 6 bottom_left_grid_pin_40_
port 6 nsew default input
rlabel metal2 s 4342 0 4398 480 6 bottom_left_grid_pin_41_
port 7 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 ccff_head
port 8 nsew default input
rlabel metal2 s 23202 27520 23258 28000 6 ccff_tail
port 9 nsew default tristate
rlabel metal3 s 0 280 480 400 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[10]
port 11 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[11]
port 12 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[12]
port 13 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[13]
port 14 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_left_in[14]
port 15 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[15]
port 16 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_left_in[16]
port 17 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[17]
port 18 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[18]
port 19 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_in[19]
port 20 nsew default input
rlabel metal3 s 0 960 480 1080 6 chanx_left_in[1]
port 21 nsew default input
rlabel metal3 s 0 1640 480 1760 6 chanx_left_in[2]
port 22 nsew default input
rlabel metal3 s 0 2320 480 2440 6 chanx_left_in[3]
port 23 nsew default input
rlabel metal3 s 0 3000 480 3120 6 chanx_left_in[4]
port 24 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[5]
port 25 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[6]
port 26 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_left_in[7]
port 27 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[8]
port 28 nsew default input
rlabel metal3 s 0 6400 480 6520 6 chanx_left_in[9]
port 29 nsew default input
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[0]
port 30 nsew default tristate
rlabel metal3 s 0 20680 480 20800 6 chanx_left_out[10]
port 31 nsew default tristate
rlabel metal3 s 0 21360 480 21480 6 chanx_left_out[11]
port 32 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[12]
port 33 nsew default tristate
rlabel metal3 s 0 22720 480 22840 6 chanx_left_out[13]
port 34 nsew default tristate
rlabel metal3 s 0 23400 480 23520 6 chanx_left_out[14]
port 35 nsew default tristate
rlabel metal3 s 0 24080 480 24200 6 chanx_left_out[15]
port 36 nsew default tristate
rlabel metal3 s 0 24760 480 24880 6 chanx_left_out[16]
port 37 nsew default tristate
rlabel metal3 s 0 25440 480 25560 6 chanx_left_out[17]
port 38 nsew default tristate
rlabel metal3 s 0 26120 480 26240 6 chanx_left_out[18]
port 39 nsew default tristate
rlabel metal3 s 0 26800 480 26920 6 chanx_left_out[19]
port 40 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[1]
port 41 nsew default tristate
rlabel metal3 s 0 15240 480 15360 6 chanx_left_out[2]
port 42 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[3]
port 43 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[4]
port 44 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[5]
port 45 nsew default tristate
rlabel metal3 s 0 17960 480 18080 6 chanx_left_out[6]
port 46 nsew default tristate
rlabel metal3 s 0 18640 480 18760 6 chanx_left_out[7]
port 47 nsew default tristate
rlabel metal3 s 0 19320 480 19440 6 chanx_left_out[8]
port 48 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[9]
port 49 nsew default tristate
rlabel metal3 s 27520 280 28000 400 6 chanx_right_in[0]
port 50 nsew default input
rlabel metal3 s 27520 7080 28000 7200 6 chanx_right_in[10]
port 51 nsew default input
rlabel metal3 s 27520 7760 28000 7880 6 chanx_right_in[11]
port 52 nsew default input
rlabel metal3 s 27520 8440 28000 8560 6 chanx_right_in[12]
port 53 nsew default input
rlabel metal3 s 27520 9120 28000 9240 6 chanx_right_in[13]
port 54 nsew default input
rlabel metal3 s 27520 9800 28000 9920 6 chanx_right_in[14]
port 55 nsew default input
rlabel metal3 s 27520 10480 28000 10600 6 chanx_right_in[15]
port 56 nsew default input
rlabel metal3 s 27520 11160 28000 11280 6 chanx_right_in[16]
port 57 nsew default input
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_in[17]
port 58 nsew default input
rlabel metal3 s 27520 12520 28000 12640 6 chanx_right_in[18]
port 59 nsew default input
rlabel metal3 s 27520 13200 28000 13320 6 chanx_right_in[19]
port 60 nsew default input
rlabel metal3 s 27520 960 28000 1080 6 chanx_right_in[1]
port 61 nsew default input
rlabel metal3 s 27520 1640 28000 1760 6 chanx_right_in[2]
port 62 nsew default input
rlabel metal3 s 27520 2320 28000 2440 6 chanx_right_in[3]
port 63 nsew default input
rlabel metal3 s 27520 3000 28000 3120 6 chanx_right_in[4]
port 64 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 chanx_right_in[5]
port 65 nsew default input
rlabel metal3 s 27520 4360 28000 4480 6 chanx_right_in[6]
port 66 nsew default input
rlabel metal3 s 27520 5040 28000 5160 6 chanx_right_in[7]
port 67 nsew default input
rlabel metal3 s 27520 5720 28000 5840 6 chanx_right_in[8]
port 68 nsew default input
rlabel metal3 s 27520 6400 28000 6520 6 chanx_right_in[9]
port 69 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_out[0]
port 70 nsew default tristate
rlabel metal3 s 27520 20680 28000 20800 6 chanx_right_out[10]
port 71 nsew default tristate
rlabel metal3 s 27520 21360 28000 21480 6 chanx_right_out[11]
port 72 nsew default tristate
rlabel metal3 s 27520 22040 28000 22160 6 chanx_right_out[12]
port 73 nsew default tristate
rlabel metal3 s 27520 22720 28000 22840 6 chanx_right_out[13]
port 74 nsew default tristate
rlabel metal3 s 27520 23400 28000 23520 6 chanx_right_out[14]
port 75 nsew default tristate
rlabel metal3 s 27520 24080 28000 24200 6 chanx_right_out[15]
port 76 nsew default tristate
rlabel metal3 s 27520 24760 28000 24880 6 chanx_right_out[16]
port 77 nsew default tristate
rlabel metal3 s 27520 25440 28000 25560 6 chanx_right_out[17]
port 78 nsew default tristate
rlabel metal3 s 27520 26120 28000 26240 6 chanx_right_out[18]
port 79 nsew default tristate
rlabel metal3 s 27520 26800 28000 26920 6 chanx_right_out[19]
port 80 nsew default tristate
rlabel metal3 s 27520 14560 28000 14680 6 chanx_right_out[1]
port 81 nsew default tristate
rlabel metal3 s 27520 15240 28000 15360 6 chanx_right_out[2]
port 82 nsew default tristate
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_out[3]
port 83 nsew default tristate
rlabel metal3 s 27520 16600 28000 16720 6 chanx_right_out[4]
port 84 nsew default tristate
rlabel metal3 s 27520 17280 28000 17400 6 chanx_right_out[5]
port 85 nsew default tristate
rlabel metal3 s 27520 17960 28000 18080 6 chanx_right_out[6]
port 86 nsew default tristate
rlabel metal3 s 27520 18640 28000 18760 6 chanx_right_out[7]
port 87 nsew default tristate
rlabel metal3 s 27520 19320 28000 19440 6 chanx_right_out[8]
port 88 nsew default tristate
rlabel metal3 s 27520 20000 28000 20120 6 chanx_right_out[9]
port 89 nsew default tristate
rlabel metal2 s 4894 0 4950 480 6 chany_bottom_in[0]
port 90 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chany_bottom_in[10]
port 91 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[11]
port 92 nsew default input
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_in[12]
port 93 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[13]
port 94 nsew default input
rlabel metal2 s 13082 0 13138 480 6 chany_bottom_in[14]
port 95 nsew default input
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_in[15]
port 96 nsew default input
rlabel metal2 s 14278 0 14334 480 6 chany_bottom_in[16]
port 97 nsew default input
rlabel metal2 s 14830 0 14886 480 6 chany_bottom_in[17]
port 98 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[18]
port 99 nsew default input
rlabel metal2 s 16026 0 16082 480 6 chany_bottom_in[19]
port 100 nsew default input
rlabel metal2 s 5538 0 5594 480 6 chany_bottom_in[1]
port 101 nsew default input
rlabel metal2 s 6090 0 6146 480 6 chany_bottom_in[2]
port 102 nsew default input
rlabel metal2 s 6642 0 6698 480 6 chany_bottom_in[3]
port 103 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chany_bottom_in[4]
port 104 nsew default input
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_in[5]
port 105 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[6]
port 106 nsew default input
rlabel metal2 s 9034 0 9090 480 6 chany_bottom_in[7]
port 107 nsew default input
rlabel metal2 s 9586 0 9642 480 6 chany_bottom_in[8]
port 108 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[9]
port 109 nsew default input
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_out[0]
port 110 nsew default tristate
rlabel metal2 s 22374 0 22430 480 6 chany_bottom_out[10]
port 111 nsew default tristate
rlabel metal2 s 23018 0 23074 480 6 chany_bottom_out[11]
port 112 nsew default tristate
rlabel metal2 s 23570 0 23626 480 6 chany_bottom_out[12]
port 113 nsew default tristate
rlabel metal2 s 24122 0 24178 480 6 chany_bottom_out[13]
port 114 nsew default tristate
rlabel metal2 s 24766 0 24822 480 6 chany_bottom_out[14]
port 115 nsew default tristate
rlabel metal2 s 25318 0 25374 480 6 chany_bottom_out[15]
port 116 nsew default tristate
rlabel metal2 s 25870 0 25926 480 6 chany_bottom_out[16]
port 117 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[17]
port 118 nsew default tristate
rlabel metal2 s 27066 0 27122 480 6 chany_bottom_out[18]
port 119 nsew default tristate
rlabel metal2 s 27618 0 27674 480 6 chany_bottom_out[19]
port 120 nsew default tristate
rlabel metal2 s 17130 0 17186 480 6 chany_bottom_out[1]
port 121 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 chany_bottom_out[2]
port 122 nsew default tristate
rlabel metal2 s 18326 0 18382 480 6 chany_bottom_out[3]
port 123 nsew default tristate
rlabel metal2 s 18878 0 18934 480 6 chany_bottom_out[4]
port 124 nsew default tristate
rlabel metal2 s 19522 0 19578 480 6 chany_bottom_out[5]
port 125 nsew default tristate
rlabel metal2 s 20074 0 20130 480 6 chany_bottom_out[6]
port 126 nsew default tristate
rlabel metal2 s 20626 0 20682 480 6 chany_bottom_out[7]
port 127 nsew default tristate
rlabel metal2 s 21270 0 21326 480 6 chany_bottom_out[8]
port 128 nsew default tristate
rlabel metal2 s 21822 0 21878 480 6 chany_bottom_out[9]
port 129 nsew default tristate
rlabel metal3 s 0 27480 480 27600 6 left_top_grid_pin_1_
port 130 nsew default input
rlabel metal2 s 4618 27520 4674 28000 6 prog_clk
port 131 nsew default input
rlabel metal3 s 27520 27480 28000 27600 6 right_top_grid_pin_1_
port 132 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 133 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 134 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
