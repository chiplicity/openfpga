VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_3__0_
  CLASS BLOCK ;
  FOREIGN sb_3__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 137.010 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 2.400 ;
    END
  END address[5]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 2.400 2.680 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 2.400 23.080 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 2.400 28.520 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.400 33.280 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.400 38.720 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 2.400 44.160 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.400 95.840 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 2.400 106.040 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 2.400 111.480 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.400 116.240 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 2.400 121.680 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 2.400 127.120 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 2.400 131.880 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 2.400 137.320 ;
    END
  END chanx_left_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 137.600 2.670 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 137.600 7.730 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 137.600 12.790 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 137.600 17.850 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 137.600 23.370 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 137.600 28.430 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 137.600 33.490 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 137.600 38.550 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 137.600 44.070 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.310 137.600 95.590 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 137.600 100.650 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.890 137.600 106.170 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.950 137.600 111.230 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.010 137.600 116.290 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.070 137.600 121.350 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 126.590 137.600 126.870 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.650 137.600 131.930 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 136.710 137.600 136.990 140.000 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.400 80.200 ;
    END
  END left_bottom_grid_pin_11_
  PIN left_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 2.400 85.640 ;
    END
  END left_bottom_grid_pin_13_
  PIN left_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 2.400 90.400 ;
    END
  END left_bottom_grid_pin_15_
  PIN left_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 2.400 54.360 ;
    END
  END left_bottom_grid_pin_1_
  PIN left_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 2.400 59.120 ;
    END
  END left_bottom_grid_pin_3_
  PIN left_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 2.400 64.560 ;
    END
  END left_bottom_grid_pin_5_
  PIN left_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.400 70.000 ;
    END
  END left_bottom_grid_pin_7_
  PIN left_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 2.400 74.760 ;
    END
  END left_bottom_grid_pin_9_
  PIN left_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.400 48.920 ;
    END
  END left_top_grid_pin_10_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 137.600 49.130 140.000 ;
    END
  END top_left_grid_pin_13_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.670 137.600 79.950 140.000 ;
    END
  END top_right_grid_pin_11_
  PIN top_right_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.190 137.600 85.470 140.000 ;
    END
  END top_right_grid_pin_13_
  PIN top_right_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.250 137.600 90.530 140.000 ;
    END
  END top_right_grid_pin_15_
  PIN top_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.910 137.600 54.190 140.000 ;
    END
  END top_right_grid_pin_1_
  PIN top_right_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 137.600 59.250 140.000 ;
    END
  END top_right_grid_pin_3_
  PIN top_right_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.490 137.600 64.770 140.000 ;
    END
  END top_right_grid_pin_5_
  PIN top_right_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 137.600 69.830 140.000 ;
    END
  END top_right_grid_pin_7_
  PIN top_right_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 137.600 74.890 140.000 ;
    END
  END top_right_grid_pin_9_
  PIN vpwr
    USE POWER ;
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    USE GROUND ;
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.530 0.380 137.010 131.200 ;
      LAYER met2 ;
        RECT 0.550 137.320 2.110 137.770 ;
        RECT 2.950 137.320 7.170 137.770 ;
        RECT 8.010 137.320 12.230 137.770 ;
        RECT 13.070 137.320 17.290 137.770 ;
        RECT 18.130 137.320 22.810 137.770 ;
        RECT 23.650 137.320 27.870 137.770 ;
        RECT 28.710 137.320 32.930 137.770 ;
        RECT 33.770 137.320 37.990 137.770 ;
        RECT 38.830 137.320 43.510 137.770 ;
        RECT 44.350 137.320 48.570 137.770 ;
        RECT 49.410 137.320 53.630 137.770 ;
        RECT 54.470 137.320 58.690 137.770 ;
        RECT 59.530 137.320 64.210 137.770 ;
        RECT 65.050 137.320 69.270 137.770 ;
        RECT 70.110 137.320 74.330 137.770 ;
        RECT 75.170 137.320 79.390 137.770 ;
        RECT 80.230 137.320 84.910 137.770 ;
        RECT 85.750 137.320 89.970 137.770 ;
        RECT 90.810 137.320 95.030 137.770 ;
        RECT 95.870 137.320 100.090 137.770 ;
        RECT 100.930 137.320 105.610 137.770 ;
        RECT 106.450 137.320 110.670 137.770 ;
        RECT 111.510 137.320 115.730 137.770 ;
        RECT 116.570 137.320 120.790 137.770 ;
        RECT 121.630 137.320 126.310 137.770 ;
        RECT 127.150 137.320 131.370 137.770 ;
        RECT 132.210 137.320 136.430 137.770 ;
        RECT 0.550 2.680 136.980 137.320 ;
        RECT 0.550 0.270 8.550 2.680 ;
        RECT 9.390 0.270 26.030 2.680 ;
        RECT 26.870 0.270 43.510 2.680 ;
        RECT 44.350 0.270 60.990 2.680 ;
        RECT 61.830 0.270 78.470 2.680 ;
        RECT 79.310 0.270 95.950 2.680 ;
        RECT 96.790 0.270 113.430 2.680 ;
        RECT 114.270 0.270 130.910 2.680 ;
        RECT 131.750 0.270 136.980 2.680 ;
      LAYER met3 ;
        RECT 0.310 137.720 130.115 137.865 ;
        RECT 2.800 136.320 130.115 137.720 ;
        RECT 0.310 132.280 130.115 136.320 ;
        RECT 2.800 130.880 130.115 132.280 ;
        RECT 0.310 127.520 130.115 130.880 ;
        RECT 2.800 126.120 130.115 127.520 ;
        RECT 0.310 122.080 130.115 126.120 ;
        RECT 2.800 120.680 130.115 122.080 ;
        RECT 0.310 116.640 130.115 120.680 ;
        RECT 2.800 115.240 130.115 116.640 ;
        RECT 0.310 111.880 130.115 115.240 ;
        RECT 2.800 110.480 130.115 111.880 ;
        RECT 0.310 106.440 130.115 110.480 ;
        RECT 2.800 105.040 130.115 106.440 ;
        RECT 0.310 101.000 130.115 105.040 ;
        RECT 2.800 99.600 130.115 101.000 ;
        RECT 0.310 96.240 130.115 99.600 ;
        RECT 2.800 94.840 130.115 96.240 ;
        RECT 0.310 90.800 130.115 94.840 ;
        RECT 2.800 89.400 130.115 90.800 ;
        RECT 0.310 86.040 130.115 89.400 ;
        RECT 2.800 84.640 130.115 86.040 ;
        RECT 0.310 80.600 130.115 84.640 ;
        RECT 2.800 79.200 130.115 80.600 ;
        RECT 0.310 75.160 130.115 79.200 ;
        RECT 2.800 73.760 130.115 75.160 ;
        RECT 0.310 70.400 130.115 73.760 ;
        RECT 2.800 69.000 130.115 70.400 ;
        RECT 0.310 64.960 130.115 69.000 ;
        RECT 2.800 63.560 130.115 64.960 ;
        RECT 0.310 59.520 130.115 63.560 ;
        RECT 2.800 58.120 130.115 59.520 ;
        RECT 0.310 54.760 130.115 58.120 ;
        RECT 2.800 53.360 130.115 54.760 ;
        RECT 0.310 49.320 130.115 53.360 ;
        RECT 2.800 47.920 130.115 49.320 ;
        RECT 0.310 44.560 130.115 47.920 ;
        RECT 2.800 43.160 130.115 44.560 ;
        RECT 0.310 39.120 130.115 43.160 ;
        RECT 2.800 37.720 130.115 39.120 ;
        RECT 0.310 33.680 130.115 37.720 ;
        RECT 2.800 32.280 130.115 33.680 ;
        RECT 0.310 28.920 130.115 32.280 ;
        RECT 2.800 27.520 130.115 28.920 ;
        RECT 0.310 23.480 130.115 27.520 ;
        RECT 2.800 22.080 130.115 23.480 ;
        RECT 0.310 18.040 130.115 22.080 ;
        RECT 2.800 16.640 130.115 18.040 ;
        RECT 0.310 13.280 130.115 16.640 ;
        RECT 2.800 11.880 130.115 13.280 ;
        RECT 0.310 7.840 130.115 11.880 ;
        RECT 2.800 6.440 130.115 7.840 ;
        RECT 0.310 3.080 130.115 6.440 ;
        RECT 2.800 2.680 130.115 3.080 ;
      LAYER met4 ;
        RECT 14.095 128.480 122.985 137.865 ;
        RECT 14.095 10.640 27.655 128.480 ;
        RECT 30.055 10.640 50.985 128.480 ;
        RECT 53.385 10.640 122.985 128.480 ;
      LAYER met5 ;
        RECT 30.020 109.700 95.100 114.700 ;
  END
END sb_3__0_
END LIBRARY

