* NGSPICE file created from sb_0__3_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt sb_0__3_ address[0] address[1] address[2] address[3] address[4] address[5]
+ bottom_left_grid_pin_11_ bottom_left_grid_pin_13_ bottom_left_grid_pin_15_ bottom_left_grid_pin_1_
+ bottom_left_grid_pin_3_ bottom_left_grid_pin_5_ bottom_left_grid_pin_7_ bottom_left_grid_pin_9_
+ bottom_right_grid_pin_11_ chanx_right_in[0] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4]
+ chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_out[0]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ data_in enable right_bottom_grid_pin_12_ right_top_grid_pin_11_ right_top_grid_pin_13_
+ right_top_grid_pin_15_ right_top_grid_pin_1_ right_top_grid_pin_3_ right_top_grid_pin_5_
+ right_top_grid_pin_7_ right_top_grid_pin_9_ vpwr vgnd
Xmem_right_track_12.LATCH_1_.latch data_in _184_/A _131_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_258 vgnd vpwr scs8hd_decap_4
XFILLER_27_236 vpwr vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _184_/A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XANTENNA__108__B enable vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_173 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_200_ _200_/A _200_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_228 vpwr vgnd scs8hd_fill_2
X_131_ _135_/A _131_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_86 vgnd vpwr scs8hd_decap_12
XFILLER_2_154 vpwr vgnd scs8hd_fill_2
XANTENNA__110__C _118_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_68 vpwr vgnd scs8hd_fill_2
XANTENNA__119__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_250 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _239_/A vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _191_/Y mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_213 vpwr vgnd scs8hd_fill_2
X_114_ _113_/Y _118_/B vgnd vpwr scs8hd_buf_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _221_/HI _188_/Y mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
XFILLER_37_172 vgnd vpwr scs8hd_decap_8
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XFILLER_4_238 vgnd vpwr scs8hd_decap_3
XFILLER_29_74 vgnd vpwr scs8hd_decap_12
XANTENNA__116__B _116_/B vgnd vpwr scs8hd_diode_2
XANTENNA__132__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_6_67 vgnd vpwr scs8hd_decap_3
XFILLER_6_56 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_172 vpwr vgnd scs8hd_fill_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_1_.latch data_in _180_/A _124_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_208 vpwr vgnd scs8hd_fill_2
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_15_98 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _179_/A mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _205_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _183_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
XFILLER_22_178 vgnd vpwr scs8hd_decap_4
XFILLER_22_145 vpwr vgnd scs8hd_fill_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_3
XFILLER_13_101 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XFILLER_3_46 vpwr vgnd scs8hd_fill_2
XFILLER_3_35 vgnd vpwr scs8hd_decap_4
XFILLER_3_24 vgnd vpwr scs8hd_decap_4
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XANTENNA__230__A _230_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XFILLER_18_215 vgnd vpwr scs8hd_decap_3
XANTENNA__124__B _125_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _191_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__140__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_4
X_130_ _123_/A _118_/B _100_/A _115_/D _131_/B vgnd vpwr scs8hd_or4_4
XFILLER_23_240 vpwr vgnd scs8hd_fill_2
XFILLER_23_98 vgnd vpwr scs8hd_decap_12
XFILLER_2_122 vpwr vgnd scs8hd_fill_2
XANTENNA__110__D _118_/D vgnd vpwr scs8hd_diode_2
XANTENNA__119__B _120_/B vgnd vpwr scs8hd_diode_2
XANTENNA__135__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _207_/A vgnd
+ vpwr scs8hd_diode_2
X_113_ address[2] _113_/Y vgnd vpwr scs8hd_inv_8
XFILLER_11_265 vpwr vgnd scs8hd_fill_2
XFILLER_11_254 vpwr vgnd scs8hd_fill_2
XFILLER_7_236 vgnd vpwr scs8hd_fill_1
XFILLER_7_258 vpwr vgnd scs8hd_fill_2
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _185_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _187_/A mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_8
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_29_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_162 vpwr vgnd scs8hd_fill_2
XFILLER_19_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_187 vpwr vgnd scs8hd_fill_2
XFILLER_25_110 vgnd vpwr scs8hd_decap_12
XFILLER_15_66 vgnd vpwr scs8hd_fill_1
XFILLER_31_98 vgnd vpwr scs8hd_decap_12
XANTENNA__233__A _233_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _127_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_135 vgnd vpwr scs8hd_decap_12
XFILLER_16_176 vpwr vgnd scs8hd_fill_2
XFILLER_16_154 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _193_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__143__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XFILLER_13_135 vpwr vgnd scs8hd_fill_2
XANTENNA__228__A _228_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _235_/A vgnd vpwr scs8hd_inv_1
XANTENNA__138__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XFILLER_8_150 vgnd vpwr scs8hd_fill_1
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_149 vpwr vgnd scs8hd_fill_2
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XANTENNA__140__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_208 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_230 vgnd vpwr scs8hd_decap_3
XFILLER_2_145 vpwr vgnd scs8hd_fill_2
XANTENNA__241__A _241_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_189 vpwr vgnd scs8hd_fill_2
XFILLER_0_37 vpwr vgnd scs8hd_fill_2
X_189_ _189_/A _189_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__135__B _136_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_79 vpwr vgnd scs8hd_fill_2
XANTENNA__151__A _136_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_211 vgnd vpwr scs8hd_fill_1
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
X_112_ _120_/A _112_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__236__A _236_/A vgnd vpwr scs8hd_diode_2
XANTENNA__146__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_1_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _174_/A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_56 vgnd vpwr scs8hd_decap_12
XFILLER_28_141 vgnd vpwr scs8hd_decap_12
XFILLER_29_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_273 vgnd vpwr scs8hd_decap_4
XFILLER_3_240 vpwr vgnd scs8hd_fill_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_166 vpwr vgnd scs8hd_fill_2
XFILLER_16_144 vpwr vgnd scs8hd_fill_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_147 vgnd vpwr scs8hd_decap_12
XANTENNA__143__B _110_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_158 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_4.LATCH_1_.latch data_in _176_/A _116_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_169 vgnd vpwr scs8hd_decap_4
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _224_/HI _178_/Y mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__138__B _137_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XANTENNA__154__A _152_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_180 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_15_ mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_128 vpwr vgnd scs8hd_fill_2
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XFILLER_18_206 vpwr vgnd scs8hd_fill_2
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XANTENNA__239__A _239_/A vgnd vpwr scs8hd_diode_2
XANTENNA__140__C _139_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_187 vpwr vgnd scs8hd_fill_2
XFILLER_5_143 vpwr vgnd scs8hd_fill_2
XANTENNA__149__A address[3] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _206_/A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
X_188_ _188_/A _188_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _182_/A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__151__B _149_/X vgnd vpwr scs8hd_diode_2
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_245 vpwr vgnd scs8hd_fill_2
XFILLER_18_56 vgnd vpwr scs8hd_decap_12
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_18_78 vgnd vpwr scs8hd_decap_12
XFILLER_11_223 vpwr vgnd scs8hd_fill_2
XFILLER_11_201 vpwr vgnd scs8hd_fill_2
X_111_ _127_/A _112_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__146__B _118_/B vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_37_197 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_219 vgnd vpwr scs8hd_decap_4
XFILLER_20_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _225_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XFILLER_19_142 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _220_/HI _186_/Y mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_123 vgnd vpwr scs8hd_decap_12
XFILLER_25_178 vgnd vpwr scs8hd_decap_3
XFILLER_25_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_244 vpwr vgnd scs8hd_fill_2
XFILLER_16_189 vpwr vgnd scs8hd_fill_2
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_159 vgnd vpwr scs8hd_decap_12
XANTENNA__143__C _139_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_259 vpwr vgnd scs8hd_fill_2
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_26_56 vgnd vpwr scs8hd_decap_12
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_148 vpwr vgnd scs8hd_fill_2
XFILLER_9_119 vgnd vpwr scs8hd_decap_3
XFILLER_3_16 vgnd vpwr scs8hd_fill_1
Xmux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _177_/A mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__154__B _153_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_185 vpwr vgnd scs8hd_fill_2
XFILLER_8_174 vpwr vgnd scs8hd_fill_2
XFILLER_8_163 vpwr vgnd scs8hd_fill_2
XANTENNA__170__A _118_/D vgnd vpwr scs8hd_diode_2
XFILLER_27_207 vgnd vpwr scs8hd_fill_1
XFILLER_18_229 vgnd vpwr scs8hd_decap_8
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_273 vpwr vgnd scs8hd_fill_2
XFILLER_5_111 vpwr vgnd scs8hd_fill_2
XANTENNA__140__D _140_/D vgnd vpwr scs8hd_diode_2
XFILLER_5_177 vgnd vpwr scs8hd_decap_6
XANTENNA__149__B _118_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__165__A _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XFILLER_23_265 vpwr vgnd scs8hd_fill_2
XFILLER_23_254 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_13_ mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_169 vgnd vpwr scs8hd_decap_4
XFILLER_2_158 vpwr vgnd scs8hd_fill_2
XFILLER_0_17 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
XFILLER_9_59 vpwr vgnd scs8hd_fill_2
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
X_187_ _187_/A _187_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_180 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _181_/Y mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_224 vpwr vgnd scs8hd_fill_2
XFILLER_20_202 vgnd vpwr scs8hd_fill_1
XFILLER_18_68 vgnd vpwr scs8hd_decap_6
X_110_ _118_/A _110_/B _118_/C _118_/D _112_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _204_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XFILLER_7_239 vgnd vpwr scs8hd_decap_3
XFILLER_7_228 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd
+ vpwr scs8hd_diode_2
X_239_ _239_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__146__C _139_/X vgnd vpwr scs8hd_diode_2
XANTENNA__162__B _160_/X vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_250 vgnd vpwr scs8hd_decap_8
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
XFILLER_1_60 vgnd vpwr scs8hd_fill_1
XFILLER_28_154 vgnd vpwr scs8hd_decap_8
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_19_121 vgnd vpwr scs8hd_fill_1
XFILLER_19_110 vgnd vpwr scs8hd_decap_8
XANTENNA__157__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_19_176 vgnd vpwr scs8hd_decap_4
XANTENNA__173__A _173_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_135 vgnd vpwr scs8hd_decap_6
Xmux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _185_/A mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_113 vgnd vpwr scs8hd_decap_3
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__143__D _143_/D vgnd vpwr scs8hd_diode_2
XANTENNA__168__A _115_/D vgnd vpwr scs8hd_diode_2
XFILLER_22_149 vgnd vpwr scs8hd_decap_4
XFILLER_22_105 vgnd vpwr scs8hd_decap_12
XFILLER_38_271 vgnd vpwr scs8hd_decap_4
XFILLER_26_68 vgnd vpwr scs8hd_decap_12
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XANTENNA__170__B _170_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_263 vgnd vpwr scs8hd_decap_12
XFILLER_27_219 vpwr vgnd scs8hd_fill_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _206_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_right_track_0.LATCH_1_.latch data_in _172_/A _105_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ _189_/Y mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_5_156 vpwr vgnd scs8hd_fill_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _184_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__149__C _139_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__165__B _163_/X vgnd vpwr scs8hd_diode_2
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vpwr vgnd scs8hd_fill_2
XFILLER_23_222 vpwr vgnd scs8hd_fill_2
XFILLER_2_104 vgnd vpwr scs8hd_fill_1
XFILLER_3_6 vpwr vgnd scs8hd_fill_2
XFILLER_2_137 vpwr vgnd scs8hd_fill_2
XFILLER_0_29 vpwr vgnd scs8hd_fill_2
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
X_186_ _186_/A _186_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _177_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_258 vgnd vpwr scs8hd_decap_12
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
XFILLER_11_258 vpwr vgnd scs8hd_fill_2
XFILLER_11_236 vpwr vgnd scs8hd_fill_2
XFILLER_7_207 vgnd vpwr scs8hd_decap_4
XFILLER_1_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _192_/A vgnd
+ vpwr scs8hd_diode_2
X_169_ _115_/D _170_/B _169_/C _169_/Y vgnd vpwr scs8hd_nor3_4
X_238_ _238_/A chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
Xmux_right_track_10.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_11_ mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__146__D _140_/D vgnd vpwr scs8hd_diode_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_7.LATCH_0_.latch data_in _197_/A _156_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_155 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_210 vpwr vgnd scs8hd_fill_2
XFILLER_19_199 vpwr vgnd scs8hd_fill_2
XFILLER_19_155 vpwr vgnd scs8hd_fill_2
XANTENNA__157__C _139_/X vgnd vpwr scs8hd_diode_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XFILLER_0_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vgnd vpwr scs8hd_decap_6
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _172_/A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _170_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_128 vgnd vpwr scs8hd_decap_6
XFILLER_22_117 vgnd vpwr scs8hd_decap_8
XANTENNA__184__A _184_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_80 vgnd vpwr scs8hd_decap_12
XFILLER_12_194 vgnd vpwr scs8hd_decap_3
XFILLER_8_143 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _179_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__170__C _152_/X vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _179_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_35_253 vpwr vgnd scs8hd_fill_2
XFILLER_35_275 vpwr vgnd scs8hd_fill_2
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_109 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.tap_buf4_0_.scs8hd_inv_1 mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _228_/A vgnd vpwr scs8hd_inv_1
XFILLER_26_231 vgnd vpwr scs8hd_decap_8
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XANTENNA__149__D _143_/D vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _223_/HI _176_/Y mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_59 vpwr vgnd scs8hd_fill_2
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
XFILLER_14_201 vpwr vgnd scs8hd_fill_2
X_185_ _185_/A _185_/Y vgnd vpwr scs8hd_inv_8
XFILLER_14_267 vgnd vpwr scs8hd_decap_8
XFILLER_9_39 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_193 vgnd vpwr scs8hd_decap_4
XFILLER_1_171 vgnd vpwr scs8hd_decap_3
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _204_/A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_168_ _115_/D _170_/B _152_/X _168_/Y vgnd vpwr scs8hd_nor3_4
X_237_ _237_/A chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_24_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_230 vgnd vpwr scs8hd_decap_6
X_099_ address[4] address[5] _100_/A vgnd vpwr scs8hd_or2_4
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XFILLER_1_84 vpwr vgnd scs8hd_fill_2
XFILLER_1_62 vgnd vpwr scs8hd_decap_6
XFILLER_1_40 vpwr vgnd scs8hd_fill_2
XANTENNA__187__A _187_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XANTENNA__097__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_28_167 vgnd vpwr scs8hd_decap_12
XFILLER_28_189 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_15.LATCH_0_.latch data_in _205_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_93 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_123 vgnd vpwr scs8hd_decap_4
XANTENNA__157__D _143_/D vgnd vpwr scs8hd_diode_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_0_269 vgnd vpwr scs8hd_decap_8
XFILLER_0_258 vpwr vgnd scs8hd_fill_2
XFILLER_0_203 vpwr vgnd scs8hd_fill_2
XFILLER_16_148 vgnd vpwr scs8hd_decap_3
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_159 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__168__C _152_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_72 vgnd vpwr scs8hd_decap_3
XFILLER_7_83 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_15_ mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_6.tap_buf4_0_.scs8hd_inv_1 mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _231_/A vgnd vpwr scs8hd_inv_1
XFILLER_38_251 vgnd vpwr scs8hd_decap_4
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_151 vgnd vpwr scs8hd_decap_6
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _219_/HI _184_/Y mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_3
XFILLER_21_173 vgnd vpwr scs8hd_decap_4
XFILLER_29_240 vgnd vpwr scs8hd_decap_4
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_12_184 vgnd vpwr scs8hd_decap_8
XFILLER_8_122 vgnd vpwr scs8hd_decap_3
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XANTENNA__195__A _195_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_265 vgnd vpwr scs8hd_decap_8
XFILLER_26_221 vgnd vpwr scs8hd_fill_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _241_/A vgnd vpwr scs8hd_inv_1
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_265 vpwr vgnd scs8hd_fill_2
XFILLER_17_254 vpwr vgnd scs8hd_fill_2
XFILLER_17_232 vgnd vpwr scs8hd_fill_1
XFILLER_4_191 vpwr vgnd scs8hd_fill_2
XFILLER_4_84 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _175_/A mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
X_184_ _184_/A _184_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_205 vgnd vpwr scs8hd_decap_6
XFILLER_9_261 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_205 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_098_ address[2] _110_/B vgnd vpwr scs8hd_buf_1
X_167_ _167_/A _170_/B vgnd vpwr scs8hd_buf_1
X_236_ _236_/A chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_28_179 vgnd vpwr scs8hd_fill_1
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _179_/Y mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
XFILLER_3_245 vgnd vpwr scs8hd_decap_3
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
X_219_ _219_/HI _219_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XFILLER_25_149 vpwr vgnd scs8hd_fill_2
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_3.LATCH_0_.latch data_in _193_/A _148_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_105 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_60 vgnd vpwr scs8hd_fill_1
XFILLER_39_208 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _207_/A mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_193 vgnd vpwr scs8hd_decap_4
XFILLER_15_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _207_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_141 vgnd vpwr scs8hd_decap_12
XFILLER_7_95 vpwr vgnd scs8hd_fill_2
XFILLER_7_62 vpwr vgnd scs8hd_fill_2
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _185_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_196 vgnd vpwr scs8hd_decap_3
XFILLER_29_263 vgnd vpwr scs8hd_decap_12
XFILLER_16_93 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _183_/A mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_163 vpwr vgnd scs8hd_fill_2
XFILLER_12_152 vgnd vpwr scs8hd_fill_1
XFILLER_8_189 vpwr vgnd scs8hd_fill_2
XFILLER_8_178 vpwr vgnd scs8hd_fill_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_115 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_15.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_52 vgnd vpwr scs8hd_decap_12
XFILLER_4_41 vgnd vpwr scs8hd_decap_8
XFILLER_23_236 vpwr vgnd scs8hd_fill_2
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XFILLER_23_258 vgnd vpwr scs8hd_decap_4
XFILLER_23_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _193_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_118 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_183_ _183_/A _183_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _187_/Y mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_228 vgnd vpwr scs8hd_decap_4
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
X_235_ _235_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_24_93 vgnd vpwr scs8hd_decap_12
X_097_ address[3] _118_/A vgnd vpwr scs8hd_buf_1
X_166_ address[3] address[2] address[4] _137_/Y _167_/A vgnd vpwr scs8hd_or4_4
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
XFILLER_37_147 vgnd vpwr scs8hd_decap_8
XFILLER_1_53 vgnd vpwr scs8hd_decap_4
XFILLER_1_97 vpwr vgnd scs8hd_fill_2
XFILLER_29_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _187_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_73 vgnd vpwr scs8hd_decap_8
XFILLER_3_257 vgnd vpwr scs8hd_decap_8
XFILLER_10_84 vgnd vpwr scs8hd_decap_8
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
X_149_ address[3] _118_/B _139_/X _143_/D _149_/X vgnd vpwr scs8hd_or4_4
X_218_ _218_/HI _218_/LO vgnd vpwr scs8hd_conb_1
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _237_/A vgnd vpwr scs8hd_inv_1
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
XFILLER_0_227 vgnd vpwr scs8hd_decap_6
Xmux_right_track_2.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_track_11.LATCH_0_.latch data_in _201_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _195_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_220 vpwr vgnd scs8hd_fill_2
XFILLER_29_275 vpwr vgnd scs8hd_fill_2
XFILLER_12_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_157 vgnd vpwr scs8hd_decap_4
XFILLER_8_146 vgnd vpwr scs8hd_decap_4
XFILLER_35_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_190 vpwr vgnd scs8hd_fill_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_5_127 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XFILLER_32_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_182 vpwr vgnd scs8hd_fill_2
XFILLER_4_171 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_226 vpwr vgnd scs8hd_fill_2
XFILLER_23_204 vgnd vpwr scs8hd_decap_3
X_182_ _182_/A _182_/Y vgnd vpwr scs8hd_inv_8
XFILLER_14_226 vgnd vpwr scs8hd_decap_12
XFILLER_13_51 vgnd vpwr scs8hd_decap_8
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
XFILLER_1_152 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_11_ mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__100__A _100_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_274 vgnd vpwr scs8hd_decap_3
Xmux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _222_/HI _174_/Y mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_165_ _169_/C _163_/X _165_/Y vgnd vpwr scs8hd_nor2_4
X_234_ _234_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_10_240 vgnd vpwr scs8hd_decap_4
X_096_ _129_/A _127_/A vgnd vpwr scs8hd_buf_1
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.INVTX1_0_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_39 vgnd vpwr scs8hd_decap_12
XFILLER_3_269 vpwr vgnd scs8hd_fill_2
XFILLER_3_236 vpwr vgnd scs8hd_fill_2
XFILLER_3_225 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_159 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _202_/A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_148_ _136_/A _147_/B _148_/Y vgnd vpwr scs8hd_nor2_4
X_217_ _217_/HI _217_/LO vgnd vpwr scs8hd_conb_1
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_239 vgnd vpwr scs8hd_decap_3
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vgnd vpwr scs8hd_decap_12
XFILLER_21_51 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XFILLER_15_151 vgnd vpwr scs8hd_fill_1
XFILLER_38_210 vgnd vpwr scs8hd_decap_4
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_110 vgnd vpwr scs8hd_decap_12
XFILLER_21_132 vpwr vgnd scs8hd_fill_2
XFILLER_12_132 vgnd vpwr scs8hd_fill_1
XFILLER_8_103 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__103__A _140_/D vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _212_/HI _206_/Y mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XFILLER_26_202 vgnd vpwr scs8hd_fill_1
XFILLER_5_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_235 vpwr vgnd scs8hd_fill_2
XFILLER_17_213 vpwr vgnd scs8hd_fill_2
Xmux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _218_/HI _182_/Y mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_271 vgnd vpwr scs8hd_decap_4
XFILLER_4_32 vgnd vpwr scs8hd_decap_6
XFILLER_31_260 vpwr vgnd scs8hd_fill_2
XFILLER_14_238 vgnd vpwr scs8hd_decap_3
XFILLER_14_205 vgnd vpwr scs8hd_decap_8
X_181_ _181_/A _181_/Y vgnd vpwr scs8hd_inv_8
XFILLER_22_260 vgnd vpwr scs8hd_decap_12
XFILLER_13_74 vgnd vpwr scs8hd_decap_12
Xmem_right_track_14.LATCH_0_.latch data_in _187_/A _136_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_13_260 vpwr vgnd scs8hd_fill_2
XFILLER_11_219 vpwr vgnd scs8hd_fill_2
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ _173_/A mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_095_ address[0] _129_/A vgnd vpwr scs8hd_inv_8
X_164_ _152_/X _163_/X _164_/Y vgnd vpwr scs8hd_nor2_4
X_233_ _233_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_267 vgnd vpwr scs8hd_decap_8
XANTENNA__111__A _127_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_11.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_9_ mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_97 vgnd vpwr scs8hd_fill_1
XFILLER_19_138 vpwr vgnd scs8hd_fill_2
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
XFILLER_27_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_147_ _135_/A _147_/B _147_/Y vgnd vpwr scs8hd_nor2_4
X_216_ _216_/HI _216_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__106__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _218_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_193 vpwr vgnd scs8hd_fill_2
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.INVTX1_0_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_207 vgnd vpwr scs8hd_decap_4
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_185 vpwr vgnd scs8hd_fill_2
XFILLER_24_163 vgnd vpwr scs8hd_decap_3
XFILLER_21_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_130 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _177_/Y mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_174 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _205_/A mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_5_107 vpwr vgnd scs8hd_fill_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_269 vgnd vpwr scs8hd_decap_8
XFILLER_17_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__114__A _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_88 vpwr vgnd scs8hd_fill_2
X_180_ _180_/A _180_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _208_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_272 vgnd vpwr scs8hd_decap_3
XFILLER_13_97 vpwr vgnd scs8hd_fill_2
XFILLER_13_86 vgnd vpwr scs8hd_decap_8
XFILLER_1_176 vpwr vgnd scs8hd_fill_2
XFILLER_1_132 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A _143_/D vgnd vpwr scs8hd_diode_2
XFILLER_9_210 vpwr vgnd scs8hd_fill_2
X_232_ _232_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
X_163_ _121_/Y _113_/Y _139_/A _143_/D _163_/X vgnd vpwr scs8hd_or4_4
XANTENNA__111__B _112_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _206_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _184_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_117 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _185_/Y mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_74 vgnd vpwr scs8hd_decap_12
X_215_ _215_/HI _215_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
X_146_ address[3] _118_/B _139_/X _140_/D _147_/B vgnd vpwr scs8hd_or4_4
XANTENNA__122__A _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_172 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XANTENNA__117__A _120_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
X_129_ _129_/A _135_/A vgnd vpwr scs8hd_buf_1
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XFILLER_7_99 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _198_/A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _192_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_123 vpwr vgnd scs8hd_fill_2
XFILLER_29_245 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_7.LATCH_1_.latch data_in _196_/A _154_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_3.INVTX1_0_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_167 vgnd vpwr scs8hd_decap_4
XFILLER_12_112 vgnd vpwr scs8hd_fill_1
XFILLER_8_127 vgnd vpwr scs8hd_decap_3
XFILLER_35_259 vpwr vgnd scs8hd_fill_2
XFILLER_7_171 vpwr vgnd scs8hd_fill_2
XFILLER_26_248 vgnd vpwr scs8hd_decap_8
XFILLER_26_215 vgnd vpwr scs8hd_decap_6
XFILLER_5_119 vgnd vpwr scs8hd_fill_1
XFILLER_40_251 vgnd vpwr scs8hd_decap_4
XFILLER_27_74 vgnd vpwr scs8hd_decap_12
XANTENNA__130__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_163 vpwr vgnd scs8hd_fill_2
XFILLER_4_67 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _186_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_199 vpwr vgnd scs8hd_fill_2
XFILLER_13_273 vgnd vpwr scs8hd_decap_4
XFILLER_13_240 vpwr vgnd scs8hd_fill_2
XFILLER_9_266 vgnd vpwr scs8hd_decap_8
XANTENNA__125__A _120_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _179_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_162_ _169_/C _160_/X _162_/Y vgnd vpwr scs8hd_nor2_4
X_231_ _231_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_10_221 vgnd vpwr scs8hd_decap_4
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XFILLER_6_236 vgnd vpwr scs8hd_fill_1
Xmem_right_track_10.LATCH_0_.latch data_in _183_/A _128_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_68 vgnd vpwr scs8hd_fill_1
XFILLER_1_57 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _194_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_129 vgnd vpwr scs8hd_decap_12
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_206 vpwr vgnd scs8hd_fill_2
XFILLER_19_118 vgnd vpwr scs8hd_fill_1
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_decap_6
XFILLER_27_162 vpwr vgnd scs8hd_fill_2
XFILLER_19_86 vgnd vpwr scs8hd_decap_12
X_145_ _136_/A _144_/B _145_/Y vgnd vpwr scs8hd_nor2_4
X_214_ _214_/HI _214_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _217_/HI _172_/Y mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
XFILLER_2_250 vpwr vgnd scs8hd_fill_2
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_98 vgnd vpwr scs8hd_decap_12
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_143 vpwr vgnd scs8hd_fill_2
XFILLER_15_110 vgnd vpwr scs8hd_decap_6
X_128_ _120_/A _127_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__117__B _116_/B vgnd vpwr scs8hd_diode_2
XANTENNA__133__A _136_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_78 vgnd vpwr scs8hd_decap_3
XFILLER_7_67 vgnd vpwr scs8hd_decap_3
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _200_/A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XFILLER_21_157 vgnd vpwr scs8hd_fill_1
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_12_146 vgnd vpwr scs8hd_decap_6
XFILLER_8_139 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_15.LATCH_1_.latch data_in _204_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__128__A _120_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_271 vgnd vpwr scs8hd_decap_4
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _181_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_86 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__130__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_186 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _211_/HI _204_/Y mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_22_230 vgnd vpwr scs8hd_decap_4
XFILLER_1_156 vpwr vgnd scs8hd_fill_2
XFILLER_1_101 vpwr vgnd scs8hd_fill_2
XANTENNA__231__A _231_/A vgnd vpwr scs8hd_diode_2
Xmem_right_track_6.LATCH_0_.latch data_in _179_/A _120_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__125__B _125_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_4
XFILLER_9_223 vpwr vgnd scs8hd_fill_2
XANTENNA__141__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_171 vgnd vpwr scs8hd_decap_12
X_161_ _152_/X _160_/X _161_/Y vgnd vpwr scs8hd_nor2_4
X_230_ _230_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
XFILLER_10_244 vgnd vpwr scs8hd_fill_1
XFILLER_6_215 vpwr vgnd scs8hd_fill_2
XANTENNA__226__A _226_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_36 vpwr vgnd scs8hd_fill_2
XFILLER_1_25 vpwr vgnd scs8hd_fill_2
XFILLER_1_14 vpwr vgnd scs8hd_fill_2
XANTENNA__136__A _136_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_270 vgnd vpwr scs8hd_decap_6
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XFILLER_3_229 vpwr vgnd scs8hd_fill_2
XFILLER_19_98 vgnd vpwr scs8hd_decap_12
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
X_144_ _135_/A _144_/B _144_/Y vgnd vpwr scs8hd_nor2_4
X_213_ _213_/HI _213_/LO vgnd vpwr scs8hd_conb_1
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.tap_buf4_0_.scs8hd_inv_1 mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _233_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_163 vpwr vgnd scs8hd_fill_2
XFILLER_18_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_199 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_127_ _127_/A _127_/B _127_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__133__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _243_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_169 vpwr vgnd scs8hd_fill_2
XFILLER_21_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_225 vgnd vpwr scs8hd_decap_8
XFILLER_29_236 vpwr vgnd scs8hd_fill_2
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_12_125 vgnd vpwr scs8hd_decap_4
XFILLER_8_107 vpwr vgnd scs8hd_fill_2
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA__234__A _234_/A vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _127_/B vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_140 vgnd vpwr scs8hd_decap_3
XFILLER_7_184 vgnd vpwr scs8hd_decap_4
XFILLER_26_206 vgnd vpwr scs8hd_decap_8
Xmux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _175_/Y mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_27_98 vgnd vpwr scs8hd_decap_12
XFILLER_17_239 vgnd vpwr scs8hd_decap_3
XFILLER_17_228 vgnd vpwr scs8hd_decap_4
XANTENNA__229__A _229_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_3.LATCH_1_.latch data_in _192_/A _147_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_132 vpwr vgnd scs8hd_fill_2
XFILLER_4_121 vgnd vpwr scs8hd_decap_4
XANTENNA__130__C _100_/A vgnd vpwr scs8hd_diode_2
XANTENNA__139__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XFILLER_23_209 vpwr vgnd scs8hd_fill_2
XFILLER_31_264 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _203_/A mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_231 vgnd vpwr scs8hd_decap_3
XANTENNA__141__B _141_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_90 vpwr vgnd scs8hd_fill_2
X_160_ _121_/Y _113_/Y _139_/A _140_/D _160_/X vgnd vpwr scs8hd_or4_4
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_44 vgnd vpwr scs8hd_decap_12
XFILLER_10_267 vgnd vpwr scs8hd_decap_8
XFILLER_10_256 vgnd vpwr scs8hd_decap_8
XFILLER_10_212 vpwr vgnd scs8hd_fill_2
XANTENNA__242__A _242_/A vgnd vpwr scs8hd_diode_2
XANTENNA__136__B _136_/B vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_260 vpwr vgnd scs8hd_fill_2
XFILLER_10_68 vpwr vgnd scs8hd_fill_2
X_212_ _212_/HI _212_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_27_175 vgnd vpwr scs8hd_decap_4
XANTENNA__237__A _237_/A vgnd vpwr scs8hd_diode_2
X_143_ _118_/A _110_/B _139_/X _143_/D _144_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _207_/Y mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XFILLER_18_142 vgnd vpwr scs8hd_decap_4
XFILLER_18_131 vpwr vgnd scs8hd_fill_2
XANTENNA__147__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _219_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_189 vgnd vpwr scs8hd_decap_4
XFILLER_24_145 vgnd vpwr scs8hd_decap_8
Xmux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _183_/Y mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_178 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_126_ _123_/A _110_/B _118_/C _118_/D _127_/B vgnd vpwr scs8hd_or4_4
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_38_259 vgnd vpwr scs8hd_decap_12
XFILLER_29_259 vpwr vgnd scs8hd_fill_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_16_56 vgnd vpwr scs8hd_decap_12
XFILLER_12_115 vgnd vpwr scs8hd_fill_1
XFILLER_20_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _187_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__144__B _144_/B vgnd vpwr scs8hd_diode_2
X_109_ _143_/D _118_/D vgnd vpwr scs8hd_buf_1
XANTENNA__160__A _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_251 vgnd vpwr scs8hd_decap_4
XFILLER_25_273 vgnd vpwr scs8hd_decap_4
XFILLER_25_262 vgnd vpwr scs8hd_decap_4
XFILLER_25_240 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _196_/A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XANTENNA__130__D _115_/D vgnd vpwr scs8hd_diode_2
XANTENNA__155__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XFILLER_31_276 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_11.LATCH_1_.latch data_in _200_/A _161_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_22_243 vpwr vgnd scs8hd_fill_2
XFILLER_1_136 vgnd vpwr scs8hd_decap_3
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _213_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_265 vpwr vgnd scs8hd_fill_2
XFILLER_13_254 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _195_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_236 vgnd vpwr scs8hd_decap_6
XFILLER_39_184 vgnd vpwr scs8hd_decap_12
XFILLER_24_56 vgnd vpwr scs8hd_decap_12
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_239 vpwr vgnd scs8hd_fill_2
XFILLER_6_206 vgnd vpwr scs8hd_decap_8
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.LATCH_0_.latch data_in _175_/A _112_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XFILLER_27_110 vgnd vpwr scs8hd_decap_12
X_142_ _136_/A _141_/B _142_/Y vgnd vpwr scs8hd_nor2_4
X_211_ _211_/HI _211_/LO vgnd vpwr scs8hd_conb_1
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _189_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__147__B _147_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
XANTENNA__163__A _121_/Y vgnd vpwr scs8hd_diode_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XFILLER_24_168 vgnd vpwr scs8hd_decap_8
XFILLER_24_135 vgnd vpwr scs8hd_fill_1
XFILLER_21_57 vgnd vpwr scs8hd_fill_1
XFILLER_15_157 vpwr vgnd scs8hd_fill_2
X_125_ _120_/A _125_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_105 vgnd vpwr scs8hd_decap_12
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_90 vpwr vgnd scs8hd_fill_2
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XANTENNA__158__A _152_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_127 vgnd vpwr scs8hd_decap_3
XFILLER_14_190 vpwr vgnd scs8hd_fill_2
XFILLER_29_249 vgnd vpwr scs8hd_decap_4
XFILLER_16_68 vgnd vpwr scs8hd_decap_12
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _197_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_260 vgnd vpwr scs8hd_decap_12
X_108_ address[1] enable _143_/D vgnd vpwr scs8hd_nand2_4
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XANTENNA__160__B _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XFILLER_19_271 vgnd vpwr scs8hd_decap_6
XFILLER_19_260 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _201_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_167 vpwr vgnd scs8hd_fill_2
XFILLER_4_145 vpwr vgnd scs8hd_fill_2
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
XFILLER_16_252 vpwr vgnd scs8hd_fill_2
XANTENNA__171__A _118_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _209_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__166__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_196 vgnd vpwr scs8hd_decap_12
XFILLER_24_68 vgnd vpwr scs8hd_decap_12
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _210_/HI _202_/Y mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_240 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _199_/A mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
X_141_ _135_/A _141_/B _141_/Y vgnd vpwr scs8hd_nor2_4
X_210_ _210_/HI _210_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_254 vgnd vpwr scs8hd_decap_4
XFILLER_2_210 vpwr vgnd scs8hd_fill_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_147 vgnd vpwr scs8hd_decap_12
XANTENNA__163__B _113_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_14.LATCH_1_.latch data_in _186_/A _135_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
XFILLER_15_147 vgnd vpwr scs8hd_decap_4
X_124_ _127_/A _125_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XANTENNA__158__B _157_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XFILLER_28_272 vgnd vpwr scs8hd_decap_3
X_107_ _120_/A _104_/X _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_154 vpwr vgnd scs8hd_fill_2
XFILLER_7_132 vpwr vgnd scs8hd_fill_2
XANTENNA__160__C _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XANTENNA__169__A _115_/D vgnd vpwr scs8hd_diode_2
XFILLER_17_209 vpwr vgnd scs8hd_fill_2
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_8
XFILLER_31_256 vpwr vgnd scs8hd_fill_2
XANTENNA__171__B _170_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ _173_/Y mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_212 vpwr vgnd scs8hd_fill_2
XFILLER_9_249 vgnd vpwr scs8hd_fill_1
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XANTENNA__166__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__182__A _182_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XFILLER_6_219 vpwr vgnd scs8hd_fill_2
XFILLER_1_29 vgnd vpwr scs8hd_decap_4
XFILLER_1_18 vpwr vgnd scs8hd_fill_2
XFILLER_14_80 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _201_/A mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XANTENNA__177__A _177_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_27_123 vgnd vpwr scs8hd_decap_12
X_140_ _118_/A _110_/B _139_/X _140_/D _141_/B vgnd vpwr scs8hd_or4_4
XFILLER_18_167 vgnd vpwr scs8hd_decap_3
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_33_159 vgnd vpwr scs8hd_decap_12
XFILLER_18_189 vpwr vgnd scs8hd_fill_2
XANTENNA__163__C _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_50 vgnd vpwr scs8hd_decap_8
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_129 vgnd vpwr scs8hd_decap_12
XFILLER_15_126 vpwr vgnd scs8hd_fill_2
X_123_ _123_/A _110_/B _118_/C _115_/D _125_/B vgnd vpwr scs8hd_or4_4
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__190__A _190_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _205_/Y mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XFILLER_12_129 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_162 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_173 vpwr vgnd scs8hd_fill_2
X_106_ address[0] _120_/A vgnd vpwr scs8hd_buf_1
XANTENNA__160__D _140_/D vgnd vpwr scs8hd_diode_2
XFILLER_22_91 vgnd vpwr scs8hd_fill_1
XFILLER_11_184 vgnd vpwr scs8hd_decap_6
XANTENNA__169__B _170_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _185_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_93 vgnd vpwr scs8hd_fill_1
XANTENNA__095__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XFILLER_16_210 vpwr vgnd scs8hd_fill_2
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__171__C _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_3_180 vgnd vpwr scs8hd_fill_1
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_9_217 vgnd vpwr scs8hd_decap_4
XFILLER_9_206 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _194_/A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_9_ mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__166__C address[4] vgnd vpwr scs8hd_diode_2
XFILLER_8_250 vpwr vgnd scs8hd_fill_2
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
XFILLER_5_94 vpwr vgnd scs8hd_fill_2
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XFILLER_5_220 vpwr vgnd scs8hd_fill_2
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_135 vgnd vpwr scs8hd_decap_12
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_27_179 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _186_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_267 vgnd vpwr scs8hd_decap_8
XFILLER_18_113 vgnd vpwr scs8hd_decap_3
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
X_199_ _199_/A _199_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__163__D _143_/D vgnd vpwr scs8hd_diode_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_84 vgnd vpwr scs8hd_decap_8
XFILLER_2_73 vpwr vgnd scs8hd_fill_2
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _220_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _216_/HI _198_/Y mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_105 vgnd vpwr scs8hd_decap_12
XFILLER_21_27 vgnd vpwr scs8hd_decap_12
XANTENNA__098__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_23_193 vpwr vgnd scs8hd_fill_2
X_122_ _121_/Y _123_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_82 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_208 vgnd vpwr scs8hd_decap_12
XFILLER_37_241 vgnd vpwr scs8hd_decap_3
Xmem_right_track_10.LATCH_1_.latch data_in _182_/A _127_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_12_108 vgnd vpwr scs8hd_decap_4
XFILLER_20_185 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _194_/Y vgnd
+ vpwr scs8hd_diode_2
X_105_ _127_/A _104_/X _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_152 vpwr vgnd scs8hd_fill_2
XANTENNA__169__C _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_27_59 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_104 vpwr vgnd scs8hd_fill_2
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_247 vpwr vgnd scs8hd_fill_2
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _188_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_269 vpwr vgnd scs8hd_fill_2
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _214_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_80 vgnd vpwr scs8hd_decap_12
XANTENNA__166__D _137_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_73 vpwr vgnd scs8hd_fill_2
XFILLER_5_62 vpwr vgnd scs8hd_fill_2
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_206 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _181_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_254 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_7_ mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_158 vpwr vgnd scs8hd_fill_2
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _196_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_125 vgnd vpwr scs8hd_decap_4
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ _198_/A _198_/Y vgnd vpwr scs8hd_inv_8
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _209_/HI _200_/Y mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_96 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _200_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_117 vgnd vpwr scs8hd_decap_12
XFILLER_17_191 vgnd vpwr scs8hd_decap_3
Xmem_right_track_6.LATCH_1_.latch data_in _178_/A _119_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_39 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _197_/A mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_121_ address[3] _121_/Y vgnd vpwr scs8hd_inv_8
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XFILLER_14_172 vpwr vgnd scs8hd_fill_2
XFILLER_14_194 vpwr vgnd scs8hd_fill_2
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_253 vpwr vgnd scs8hd_fill_2
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
X_104_ _118_/A _110_/B _118_/C _115_/D _104_/X vgnd vpwr scs8hd_or4_4
XFILLER_22_93 vgnd vpwr scs8hd_decap_12
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_19_231 vpwr vgnd scs8hd_fill_2
XFILLER_8_84 vpwr vgnd scs8hd_fill_2
XFILLER_8_73 vpwr vgnd scs8hd_fill_2
XFILLER_8_62 vpwr vgnd scs8hd_fill_2
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vpwr vgnd scs8hd_fill_2
XFILLER_25_223 vpwr vgnd scs8hd_fill_2
XFILLER_40_259 vgnd vpwr scs8hd_decap_12
XFILLER_4_149 vpwr vgnd scs8hd_fill_2
XFILLER_4_127 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_256 vgnd vpwr scs8hd_decap_4
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_22_226 vpwr vgnd scs8hd_fill_2
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _210_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_263 vgnd vpwr scs8hd_decap_12
XFILLER_8_230 vpwr vgnd scs8hd_fill_2
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_266 vpwr vgnd scs8hd_fill_2
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_19_39 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.tap_buf4_0_.scs8hd_inv_1 mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _227_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _173_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_82 vgnd vpwr scs8hd_decap_3
XFILLER_18_148 vpwr vgnd scs8hd_fill_2
X_197_ _197_/A _197_/Y vgnd vpwr scs8hd_inv_8
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XFILLER_24_129 vgnd vpwr scs8hd_decap_6
XFILLER_17_170 vpwr vgnd scs8hd_fill_2
XFILLER_23_140 vpwr vgnd scs8hd_fill_2
XFILLER_15_118 vgnd vpwr scs8hd_decap_4
X_120_ _120_/A _120_/B _120_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_4.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_5_ mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
XFILLER_11_51 vgnd vpwr scs8hd_decap_8
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_221 vgnd vpwr scs8hd_decap_12
XFILLER_20_198 vgnd vpwr scs8hd_decap_4
XFILLER_28_243 vgnd vpwr scs8hd_decap_8
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
X_103_ _140_/D _115_/D vgnd vpwr scs8hd_buf_1
XFILLER_22_61 vgnd vpwr scs8hd_decap_12
XFILLER_11_165 vpwr vgnd scs8hd_fill_2
XFILLER_7_158 vpwr vgnd scs8hd_fill_2
XFILLER_7_136 vpwr vgnd scs8hd_fill_2
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_27_39 vgnd vpwr scs8hd_decap_12
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _203_/Y mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_16_235 vgnd vpwr scs8hd_decap_8
XFILLER_16_224 vpwr vgnd scs8hd_fill_2
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_172 vpwr vgnd scs8hd_fill_2
XFILLER_30_271 vgnd vpwr scs8hd_decap_4
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XFILLER_13_227 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_42 vpwr vgnd scs8hd_fill_2
XFILLER_39_135 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _230_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_212 vpwr vgnd scs8hd_fill_2
XANTENNA__101__A enable vgnd vpwr scs8hd_diode_2
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _192_/A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_226 vgnd vpwr scs8hd_decap_12
XFILLER_18_105 vgnd vpwr scs8hd_decap_8
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_26_193 vgnd vpwr scs8hd_decap_3
X_196_ _196_/A _196_/Y vgnd vpwr scs8hd_inv_8
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _240_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_43 vgnd vpwr scs8hd_fill_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_4
XFILLER_1_270 vgnd vpwr scs8hd_decap_6
XFILLER_17_182 vgnd vpwr scs8hd_fill_1
XFILLER_32_141 vgnd vpwr scs8hd_decap_12
XFILLER_23_163 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_74 vgnd vpwr scs8hd_decap_8
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_179_ _179_/A _179_/Y vgnd vpwr scs8hd_inv_8
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_233 vgnd vpwr scs8hd_decap_8
XFILLER_20_166 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.LATCH_1_.latch data_in _174_/A _111_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _215_/HI _196_/Y mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_102_ address[1] _102_/B _140_/D vgnd vpwr scs8hd_or2_4
XFILLER_22_73 vgnd vpwr scs8hd_decap_12
XFILLER_11_177 vgnd vpwr scs8hd_decap_6
Xmux_right_track_2.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_3_ mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_181 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _189_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_269 vpwr vgnd scs8hd_fill_2
XFILLER_25_258 vpwr vgnd scs8hd_fill_2
XFILLER_25_236 vpwr vgnd scs8hd_fill_2
XFILLER_17_62 vgnd vpwr scs8hd_decap_12
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_195 vpwr vgnd scs8hd_fill_2
XFILLER_3_151 vgnd vpwr scs8hd_decap_3
XFILLER_22_206 vgnd vpwr scs8hd_decap_8
XFILLER_0_187 vgnd vpwr scs8hd_decap_3
XFILLER_0_165 vpwr vgnd scs8hd_fill_2
XFILLER_12_272 vgnd vpwr scs8hd_decap_3
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_9.LATCH_0_.latch data_in _199_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _197_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_235 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _201_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.INVTX1_0_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_238 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_26_183 vgnd vpwr scs8hd_fill_1
XFILLER_25_62 vgnd vpwr scs8hd_decap_12
XFILLER_25_51 vgnd vpwr scs8hd_decap_8
X_195_ _195_/A _195_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__112__A _120_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_260 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _221_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_197 vpwr vgnd scs8hd_fill_2
XFILLER_23_175 vpwr vgnd scs8hd_fill_2
XFILLER_11_97 vpwr vgnd scs8hd_fill_2
XFILLER_11_86 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A _120_/A vgnd vpwr scs8hd_diode_2
X_178_ _178_/A _178_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_245 vgnd vpwr scs8hd_decap_8
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_145 vpwr vgnd scs8hd_fill_2
XFILLER_28_201 vgnd vpwr scs8hd_decap_12
X_101_ enable _102_/B vgnd vpwr scs8hd_inv_8
XFILLER_11_123 vgnd vpwr scs8hd_fill_1
XFILLER_11_101 vpwr vgnd scs8hd_fill_2
XFILLER_22_85 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _195_/A mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_19_256 vpwr vgnd scs8hd_fill_2
XFILLER_19_245 vpwr vgnd scs8hd_fill_2
XFILLER_19_212 vpwr vgnd scs8hd_fill_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_34_259 vgnd vpwr scs8hd_decap_12
XFILLER_19_267 vpwr vgnd scs8hd_fill_2
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _199_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_215 vgnd vpwr scs8hd_fill_1
XFILLER_4_108 vgnd vpwr scs8hd_decap_4
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_270 vgnd vpwr scs8hd_decap_4
XFILLER_17_74 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _203_/A vgnd
+ vpwr scs8hd_diode_2
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XANTENNA__104__B _110_/B vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _120_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_1_ mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _236_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_111 vpwr vgnd scs8hd_fill_2
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_199 vpwr vgnd scs8hd_fill_2
XFILLER_12_251 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _215_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__115__A _118_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _199_/Y mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_159 vgnd vpwr scs8hd_decap_12
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_77 vpwr vgnd scs8hd_fill_2
XFILLER_5_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _217_/HI vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_17.LATCH_0_.latch data_in _207_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XFILLER_2_206 vpwr vgnd scs8hd_fill_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XFILLER_25_74 vgnd vpwr scs8hd_decap_12
X_194_ _194_/A _194_/Y vgnd vpwr scs8hd_inv_8
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
XANTENNA__112__B _112_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_67 vgnd vpwr scs8hd_decap_4
XFILLER_2_23 vgnd vpwr scs8hd_decap_8
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_23_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.INVTX1_0_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_154 vgnd vpwr scs8hd_decap_3
XFILLER_14_143 vgnd vpwr scs8hd_decap_8
X_177_ _177_/A _177_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__107__B _104_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_176 vgnd vpwr scs8hd_decap_3
XANTENNA__123__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_20_157 vgnd vpwr scs8hd_decap_3
XFILLER_28_213 vgnd vpwr scs8hd_fill_1
X_100_ _100_/A _118_/C vgnd vpwr scs8hd_buf_1
XFILLER_11_146 vgnd vpwr scs8hd_decap_4
XFILLER_11_135 vpwr vgnd scs8hd_fill_2
XFILLER_19_235 vpwr vgnd scs8hd_fill_2
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
X_229_ _229_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_8_88 vpwr vgnd scs8hd_fill_2
XFILLER_8_77 vgnd vpwr scs8hd_decap_4
XFILLER_8_66 vgnd vpwr scs8hd_decap_4
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_205 vpwr vgnd scs8hd_fill_2
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XANTENNA__104__C _118_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__120__B _120_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_208 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _172_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
XFILLER_0_134 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_230 vpwr vgnd scs8hd_fill_2
XFILLER_8_234 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _201_/Y mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__115__B _118_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _211_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__131__A _135_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_193 vpwr vgnd scs8hd_fill_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XFILLER_39_51 vgnd vpwr scs8hd_decap_8
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_171 vgnd vpwr scs8hd_decap_12
XANTENNA__126__A _123_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_5.LATCH_0_.latch data_in _195_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_163 vgnd vpwr scs8hd_decap_12
XFILLER_26_141 vgnd vpwr scs8hd_decap_12
X_193_ _193_/A _193_/Y vgnd vpwr scs8hd_inv_8
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XFILLER_25_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_130 vpwr vgnd scs8hd_fill_2
XFILLER_2_46 vgnd vpwr scs8hd_fill_1
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_17_196 vpwr vgnd scs8hd_fill_2
XFILLER_17_174 vpwr vgnd scs8hd_fill_2
XFILLER_23_155 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _190_/A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_122 vgnd vpwr scs8hd_decap_6
X_176_ _176_/A _176_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_9_170 vpwr vgnd scs8hd_fill_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
XFILLER_11_169 vpwr vgnd scs8hd_fill_2
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XANTENNA__118__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_56 vgnd vpwr scs8hd_decap_3
X_159_ _169_/C _157_/X _159_/Y vgnd vpwr scs8hd_nor2_4
X_228_ _228_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__134__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_191 vgnd vpwr scs8hd_decap_6
XFILLER_6_184 vgnd vpwr scs8hd_decap_3
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
XFILLER_16_228 vgnd vpwr scs8hd_decap_4
XFILLER_16_206 vpwr vgnd scs8hd_fill_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XANTENNA__104__D _115_/D vgnd vpwr scs8hd_diode_2
XFILLER_3_176 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _214_/HI _194_/Y mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__129__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_220 vpwr vgnd scs8hd_fill_2
XFILLER_0_90 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_264 vgnd vpwr scs8hd_decap_8
XFILLER_8_246 vpwr vgnd scs8hd_fill_2
XANTENNA__115__C _118_/C vgnd vpwr scs8hd_diode_2
XANTENNA__131__B _131_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XFILLER_5_46 vgnd vpwr scs8hd_decap_4
XFILLER_38_161 vgnd vpwr scs8hd_decap_12
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_216 vpwr vgnd scs8hd_fill_2
XANTENNA__232__A _232_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XANTENNA__126__B _110_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _136_/A vgnd vpwr scs8hd_diode_2
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XFILLER_26_175 vgnd vpwr scs8hd_decap_8
XANTENNA__227__A _227_/A vgnd vpwr scs8hd_diode_2
X_192_ _192_/A _192_/Y vgnd vpwr scs8hd_inv_8
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
XFILLER_25_98 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_13.LATCH_0_.latch data_in _203_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_14.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_230 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_17_153 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__137__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _188_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_175_ _175_/A _175_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__C _118_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_193 vpwr vgnd scs8hd_fill_2
XFILLER_9_182 vgnd vpwr scs8hd_fill_1
XFILLER_28_215 vpwr vgnd scs8hd_fill_2
XFILLER_28_226 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_44 vgnd vpwr scs8hd_decap_12
XANTENNA__240__A _240_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_270 vgnd vpwr scs8hd_decap_6
X_227_ _227_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA__118__C _118_/C vgnd vpwr scs8hd_diode_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
X_158_ _152_/X _157_/X _158_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__B _118_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _196_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__150__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_262 vgnd vpwr scs8hd_decap_12
XFILLER_17_77 vgnd vpwr scs8hd_decap_12
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _200_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XANTENNA__235__A _235_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_199 vpwr vgnd scs8hd_fill_2
XFILLER_15_240 vpwr vgnd scs8hd_fill_2
XANTENNA__145__A _136_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _193_/A mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_265 vpwr vgnd scs8hd_fill_2
XFILLER_21_254 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_169 vgnd vpwr scs8hd_decap_3
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XANTENNA__115__D _115_/D vgnd vpwr scs8hd_diode_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_38_173 vgnd vpwr scs8hd_decap_12
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XANTENNA__126__C _118_/C vgnd vpwr scs8hd_diode_2
XANTENNA__142__B _141_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_261 vgnd vpwr scs8hd_decap_12
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _197_/Y mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XFILLER_26_198 vgnd vpwr scs8hd_decap_4
X_191_ _191_/A _191_/Y vgnd vpwr scs8hd_inv_8
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XANTENNA__243__A _243_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_15 vgnd vpwr scs8hd_decap_4
XFILLER_17_187 vpwr vgnd scs8hd_fill_2
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _198_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__153__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _202_/A vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_0_.latch data_in _191_/A _145_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XANTENNA__238__A _238_/A vgnd vpwr scs8hd_diode_2
X_243_ _243_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_14_168 vpwr vgnd scs8hd_fill_2
X_174_ _174_/A _174_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__D _115_/D vgnd vpwr scs8hd_diode_2
XANTENNA__148__A _136_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_105 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_80 vpwr vgnd scs8hd_fill_2
XFILLER_22_56 vpwr vgnd scs8hd_fill_2
XFILLER_19_216 vpwr vgnd scs8hd_fill_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
X_157_ _123_/A address[2] _139_/X _143_/D _157_/X vgnd vpwr scs8hd_or4_4
X_226_ _226_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA__134__C _100_/A vgnd vpwr scs8hd_diode_2
XANTENNA__118__D _118_/D vgnd vpwr scs8hd_diode_2
XFILLER_10_171 vgnd vpwr scs8hd_decap_8
XANTENNA__150__B _149_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_175 vgnd vpwr scs8hd_decap_6
XFILLER_6_164 vpwr vgnd scs8hd_fill_2
XFILLER_25_219 vpwr vgnd scs8hd_fill_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _173_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_274 vgnd vpwr scs8hd_decap_3
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_89 vgnd vpwr scs8hd_decap_12
Xmem_right_track_16.LATCH_0_.latch data_in _189_/A _142_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_274 vgnd vpwr scs8hd_fill_1
XFILLER_3_156 vgnd vpwr scs8hd_decap_3
XFILLER_3_134 vpwr vgnd scs8hd_fill_2
XFILLER_3_123 vpwr vgnd scs8hd_fill_2
XFILLER_3_101 vpwr vgnd scs8hd_fill_2
X_209_ _209_/HI _209_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__145__B _144_/B vgnd vpwr scs8hd_diode_2
XANTENNA__161__A _152_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_90 vpwr vgnd scs8hd_fill_2
XFILLER_0_115 vgnd vpwr scs8hd_decap_3
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_226 vpwr vgnd scs8hd_fill_2
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _216_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_10.tap_buf4_0_.scs8hd_inv_1 mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _229_/A vgnd vpwr scs8hd_inv_1
XANTENNA__156__A _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_7_270 vgnd vpwr scs8hd_decap_6
XFILLER_38_141 vgnd vpwr scs8hd_decap_12
XFILLER_38_185 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _222_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XANTENNA__126__D _118_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_273 vpwr vgnd scs8hd_fill_2
XPHY_12 vgnd vpwr scs8hd_decap_3
X_190_ _190_/A _190_/Y vgnd vpwr scs8hd_inv_8
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XFILLER_1_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_254 vgnd vpwr scs8hd_decap_4
XFILLER_17_166 vpwr vgnd scs8hd_fill_2
XANTENNA__153__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _175_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_136 vpwr vgnd scs8hd_fill_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
X_173_ _173_/A _173_/Y vgnd vpwr scs8hd_inv_8
X_242_ _242_/A chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__148__B _147_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_128 vgnd vpwr scs8hd_decap_8
XFILLER_20_117 vpwr vgnd scs8hd_fill_2
XANTENNA__164__A _152_/X vgnd vpwr scs8hd_diode_2
XFILLER_13_191 vpwr vgnd scs8hd_fill_2
XFILLER_9_184 vpwr vgnd scs8hd_fill_2
XFILLER_9_140 vpwr vgnd scs8hd_fill_2
XFILLER_11_139 vpwr vgnd scs8hd_fill_2
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XFILLER_19_239 vgnd vpwr scs8hd_decap_3
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
X_156_ _169_/C _153_/X _156_/Y vgnd vpwr scs8hd_nor2_4
X_225_ _225_/HI _225_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__134__D _118_/D vgnd vpwr scs8hd_diode_2
XFILLER_6_121 vpwr vgnd scs8hd_fill_2
XANTENNA__159__A _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XFILLER_25_209 vgnd vpwr scs8hd_decap_6
Xmux_right_track_10.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_168 vpwr vgnd scs8hd_fill_2
X_139_ _139_/A _139_/X vgnd vpwr scs8hd_buf_1
X_208_ _208_/HI _208_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__161__B _160_/X vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.tap_buf4_0_.scs8hd_inv_1 mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _232_/A vgnd vpwr scs8hd_inv_1
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_201 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XFILLER_12_234 vgnd vpwr scs8hd_decap_4
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _212_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__156__B _153_/X vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _172_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _213_/HI _192_/Y mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _242_/A vgnd vpwr scs8hd_inv_1
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XFILLER_5_208 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__167__A _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_17_101 vpwr vgnd scs8hd_fill_2
XFILLER_2_39 vgnd vpwr scs8hd_decap_4
XFILLER_1_266 vpwr vgnd scs8hd_fill_2
XFILLER_17_178 vpwr vgnd scs8hd_fill_2
XFILLER_17_156 vgnd vpwr scs8hd_fill_1
XFILLER_17_134 vpwr vgnd scs8hd_fill_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_4
XANTENNA__153__C _139_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_159 vgnd vpwr scs8hd_decap_4
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_9.LATCH_1_.latch data_in _198_/A _158_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _180_/A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
X_172_ _172_/A _172_/Y vgnd vpwr scs8hd_inv_8
X_241_ _241_/A chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__164__B _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_174 vpwr vgnd scs8hd_fill_2
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XFILLER_27_240 vpwr vgnd scs8hd_fill_2
X_224_ _224_/HI _224_/LO vgnd vpwr scs8hd_conb_1
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
X_155_ address[0] _169_/C vgnd vpwr scs8hd_buf_1
XFILLER_12_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_100 vgnd vpwr scs8hd_decap_3
XANTENNA__159__B _157_/X vgnd vpwr scs8hd_diode_2
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XFILLER_33_254 vpwr vgnd scs8hd_fill_2
XFILLER_18_251 vgnd vpwr scs8hd_decap_3
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_24_221 vgnd vpwr scs8hd_fill_1
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_232 vpwr vgnd scs8hd_fill_2
X_207_ _207_/A _207_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_202 vgnd vpwr scs8hd_decap_12
XFILLER_15_265 vgnd vpwr scs8hd_decap_12
XFILLER_15_254 vpwr vgnd scs8hd_fill_2
X_138_ address[4] _137_/Y _139_/A vgnd vpwr scs8hd_nand2_4
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_235 vpwr vgnd scs8hd_fill_2
XFILLER_0_94 vpwr vgnd scs8hd_fill_2
XFILLER_0_72 vpwr vgnd scs8hd_fill_2
XFILLER_0_139 vpwr vgnd scs8hd_fill_2
XFILLER_28_68 vgnd vpwr scs8hd_decap_12
XFILLER_8_206 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_12.LATCH_0_.latch data_in _185_/A _133_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_90 vpwr vgnd scs8hd_fill_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_4
XFILLER_38_198 vgnd vpwr scs8hd_decap_12
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _191_/A mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _199_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_80 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _188_/A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
XANTENNA__183__A _183_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _203_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XFILLER_1_234 vgnd vpwr scs8hd_decap_4
XFILLER_1_212 vgnd vpwr scs8hd_decap_3
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XANTENNA__153__D _140_/D vgnd vpwr scs8hd_diode_2
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_171 vgnd vpwr scs8hd_decap_12
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
X_240_ _240_/A chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
X_171_ _118_/D _170_/B _169_/C _171_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_22_193 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _195_/Y mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_17.LATCH_1_.latch data_in _206_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_153 vpwr vgnd scs8hd_fill_2
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
X_223_ _223_/HI _223_/LO vgnd vpwr scs8hd_conb_1
X_154_ _152_/X _153_/X _154_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_163 vpwr vgnd scs8hd_fill_2
XFILLER_6_189 vpwr vgnd scs8hd_fill_2
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
XFILLER_6_134 vpwr vgnd scs8hd_fill_2
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _238_/A vgnd vpwr scs8hd_inv_1
XANTENNA__191__A _191_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_233 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_0_.latch data_in _181_/A _125_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_137_ address[5] _137_/Y vgnd vpwr scs8hd_inv_8
X_206_ _206_/A _206_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_236 vgnd vpwr scs8hd_decap_8
XFILLER_30_247 vgnd vpwr scs8hd_decap_8
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_269 vgnd vpwr scs8hd_decap_8
XFILLER_21_258 vpwr vgnd scs8hd_fill_2
XANTENNA__186__A _186_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _205_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_107 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A _129_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _183_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_247 vpwr vgnd scs8hd_fill_2
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_243 vpwr vgnd scs8hd_fill_2
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
XFILLER_6_72 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_25_59 vpwr vgnd scs8hd_fill_2
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _191_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_19 vgnd vpwr scs8hd_fill_1
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_32_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_191 vgnd vpwr scs8hd_decap_3
XFILLER_15_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _172_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__194__A _194_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_39 vgnd vpwr scs8hd_decap_12
X_170_ _118_/D _170_/B _152_/X _170_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_14_139 vpwr vgnd scs8hd_fill_2
XFILLER_37_209 vgnd vpwr scs8hd_decap_12
XFILLER_26_80 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_7_ mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_84 vpwr vgnd scs8hd_fill_2
XFILLER_3_62 vpwr vgnd scs8hd_fill_2
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XANTENNA__099__A address[4] vgnd vpwr scs8hd_diode_2
X_153_ _123_/A address[2] _139_/X _140_/D _153_/X vgnd vpwr scs8hd_or4_4
X_222_ _222_/HI _222_/LO vgnd vpwr scs8hd_conb_1
Xmem_bottom_track_5.LATCH_1_.latch data_in _194_/A _150_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_93 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_33_245 vgnd vpwr scs8hd_decap_6
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_245 vgnd vpwr scs8hd_decap_4
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XFILLER_3_138 vpwr vgnd scs8hd_fill_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
X_136_ _136_/A _136_/B _136_/Y vgnd vpwr scs8hd_nor2_4
X_205_ _205_/A _205_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_259 vgnd vpwr scs8hd_decap_12
XFILLER_2_193 vpwr vgnd scs8hd_fill_2
XFILLER_0_85 vgnd vpwr scs8hd_decap_3
XFILLER_0_63 vpwr vgnd scs8hd_fill_2
XFILLER_0_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XFILLER_12_215 vpwr vgnd scs8hd_fill_2
XFILLER_20_270 vgnd vpwr scs8hd_decap_4
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd vpwr
+ scs8hd_diode_2
X_119_ _127_/A _120_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _223_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XFILLER_20_93 vgnd vpwr scs8hd_decap_12
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _208_/HI _190_/Y mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_32_129 vgnd vpwr scs8hd_decap_12
XFILLER_25_170 vgnd vpwr scs8hd_decap_8
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_107 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_162 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_195 vpwr vgnd scs8hd_fill_2
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XANTENNA__099__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_276 vgnd vpwr scs8hd_fill_1
XFILLER_27_254 vpwr vgnd scs8hd_fill_2
X_152_ _129_/A _152_/X vgnd vpwr scs8hd_buf_1
X_221_ _221_/HI _221_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_132 vpwr vgnd scs8hd_fill_2
XFILLER_6_158 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _178_/A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_210 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_13.LATCH_1_.latch data_in _202_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_191 vpwr vgnd scs8hd_fill_2
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_5_ mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_204_ _204_/A _204_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_227 vgnd vpwr scs8hd_decap_6
XFILLER_15_213 vpwr vgnd scs8hd_fill_2
X_135_ _135_/A _136_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_216 vpwr vgnd scs8hd_fill_2
XFILLER_9_62 vgnd vpwr scs8hd_decap_8
XFILLER_9_51 vgnd vpwr scs8hd_decap_8
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XFILLER_18_93 vgnd vpwr scs8hd_decap_12
X_118_ _118_/A _118_/B _118_/C _118_/D _120_/B vgnd vpwr scs8hd_or4_4
Xmem_right_track_4.LATCH_0_.latch data_in _177_/A _117_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A bottom_left_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_223 vgnd vpwr scs8hd_fill_1
XFILLER_4_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_52 vgnd vpwr scs8hd_fill_1
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_26_105 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_39 vgnd vpwr scs8hd_decap_12
XFILLER_1_226 vpwr vgnd scs8hd_fill_2
XFILLER_17_149 vgnd vpwr scs8hd_decap_4
XFILLER_17_127 vgnd vpwr scs8hd_fill_1
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XFILLER_16_193 vpwr vgnd scs8hd_fill_2
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _186_/A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_263 vgnd vpwr scs8hd_decap_12
XFILLER_22_174 vpwr vgnd scs8hd_fill_2
XFILLER_26_93 vgnd vpwr scs8hd_decap_12
XFILLER_13_152 vpwr vgnd scs8hd_fill_2
XFILLER_9_134 vgnd vpwr scs8hd_decap_4
XFILLER_9_123 vpwr vgnd scs8hd_fill_2
XFILLER_9_101 vpwr vgnd scs8hd_fill_2
XFILLER_9_189 vpwr vgnd scs8hd_fill_2
XFILLER_9_178 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_97 vpwr vgnd scs8hd_fill_2
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XFILLER_3_42 vpwr vgnd scs8hd_fill_2
XFILLER_3_31 vpwr vgnd scs8hd_fill_2
XFILLER_3_20 vpwr vgnd scs8hd_fill_2
X_220_ _220_/HI _220_/LO vgnd vpwr scs8hd_conb_1
XFILLER_27_266 vpwr vgnd scs8hd_fill_2
X_151_ _136_/A _149_/X _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_258 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _193_/Y mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
XFILLER_24_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _198_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
X_203_ _203_/A _203_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_258 vpwr vgnd scs8hd_fill_2
XFILLER_15_236 vpwr vgnd scs8hd_fill_2
X_134_ _123_/A _118_/B _100_/A _118_/D _136_/B vgnd vpwr scs8hd_or4_4
Xmem_bottom_track_1.LATCH_1_.latch data_in _190_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_10 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _202_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_54 vgnd vpwr scs8hd_decap_8
XFILLER_0_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_21 vgnd vpwr scs8hd_decap_8
XFILLER_21_239 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_206 vgnd vpwr scs8hd_decap_8
X_117_ _120_/A _116_/B _117_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_track_5.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_3_ mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XFILLER_7_254 vpwr vgnd scs8hd_fill_2
XFILLER_7_232 vgnd vpwr scs8hd_decap_4
XFILLER_7_276 vgnd vpwr scs8hd_fill_1
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _181_/A mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_27 vgnd vpwr scs8hd_decap_12
XFILLER_29_147 vgnd vpwr scs8hd_decap_12
XFILLER_37_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_257 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_1_.latch data_in _188_/A _141_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_26_117 vgnd vpwr scs8hd_decap_12
XFILLER_19_180 vgnd vpwr scs8hd_fill_1
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_15_62 vgnd vpwr scs8hd_decap_4
XFILLER_15_51 vgnd vpwr scs8hd_decap_8
XANTENNA__102__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_16_172 vpwr vgnd scs8hd_fill_2
XFILLER_39_275 vpwr vgnd scs8hd_fill_2
XFILLER_39_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_197 vgnd vpwr scs8hd_decap_6
XFILLER_13_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_131 vpwr vgnd scs8hd_fill_2
XFILLER_9_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _204_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_10 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_223 vpwr vgnd scs8hd_fill_2
XFILLER_27_201 vgnd vpwr scs8hd_decap_6
X_150_ _135_/A _149_/X _150_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_167 vpwr vgnd scs8hd_fill_2
XFILLER_10_145 vpwr vgnd scs8hd_fill_2
XFILLER_6_149 vpwr vgnd scs8hd_fill_2
XFILLER_6_138 vpwr vgnd scs8hd_fill_2
XFILLER_6_105 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_160 vpwr vgnd scs8hd_fill_2
XFILLER_24_215 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _175_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_204 vpwr vgnd scs8hd_fill_2
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
X_133_ _136_/A _131_/B _133_/Y vgnd vpwr scs8hd_nor2_4
X_202_ _202_/A _202_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_62 vgnd vpwr scs8hd_decap_12
XFILLER_23_51 vgnd vpwr scs8hd_decap_8
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ _189_/A mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_2_141 vpwr vgnd scs8hd_fill_2
XANTENNA__110__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_97 vpwr vgnd scs8hd_fill_2
XFILLER_9_86 vpwr vgnd scs8hd_fill_2
XFILLER_9_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd
+ vpwr scs8hd_diode_2
X_116_ _127_/A _116_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_240 vpwr vgnd scs8hd_fill_2
XFILLER_7_266 vpwr vgnd scs8hd_fill_2
XFILLER_29_159 vgnd vpwr scs8hd_decap_12
XFILLER_39_39 vgnd vpwr scs8hd_decap_12
XFILLER_37_192 vgnd vpwr scs8hd_decap_3
XFILLER_4_247 vgnd vpwr scs8hd_fill_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.INVTX1_1_.scs8hd_inv_1 bottom_left_grid_pin_1_ mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_26_129 vgnd vpwr scs8hd_decap_12
Xmem_right_track_0.LATCH_0_.latch data_in _173_/A _107_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_162 vpwr vgnd scs8hd_fill_2
XFILLER_15_74 vgnd vpwr scs8hd_decap_12
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XANTENNA__102__B _102_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_110 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_232 vgnd vpwr scs8hd_decap_12
XFILLER_22_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _177_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_13_187 vpwr vgnd scs8hd_fill_2
XFILLER_13_165 vpwr vgnd scs8hd_fill_2
XFILLER_9_114 vgnd vpwr scs8hd_decap_3
XANTENNA__113__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_66 vgnd vpwr scs8hd_decap_3
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_10_113 vpwr vgnd scs8hd_fill_2
XFILLER_6_117 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _234_/A vgnd vpwr scs8hd_inv_1
XFILLER_10_179 vgnd vpwr scs8hd_fill_1
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_246 vgnd vpwr scs8hd_decap_3
XANTENNA__108__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_32_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_132_ address[0] _136_/A vgnd vpwr scs8hd_buf_1
X_201_ _201_/A _201_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_74 vgnd vpwr scs8hd_decap_12
XFILLER_2_175 vgnd vpwr scs8hd_decap_3
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _226_/A vgnd vpwr scs8hd_inv_1
XANTENNA__110__B _110_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _176_/A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_274 vgnd vpwr scs8hd_fill_1
XFILLER_20_241 vpwr vgnd scs8hd_fill_2
XFILLER_18_74 vgnd vpwr scs8hd_fill_1
X_115_ _118_/A _118_/B _118_/C _115_/D _116_/B vgnd vpwr scs8hd_or4_4
XANTENNA__105__B _104_/X vgnd vpwr scs8hd_diode_2
XANTENNA__121__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XFILLER_37_160 vgnd vpwr scs8hd_decap_12
XFILLER_4_226 vgnd vpwr scs8hd_fill_1
XFILLER_4_204 vgnd vpwr scs8hd_decap_8
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _224_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_51 vgnd vpwr scs8hd_decap_8
XFILLER_29_62 vgnd vpwr scs8hd_decap_12
XANTENNA__116__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_88 vpwr vgnd scs8hd_fill_2
XFILLER_6_44 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _225_/HI _180_/Y mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_141 vgnd vpwr scs8hd_fill_1
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_86 vgnd vpwr scs8hd_decap_12
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XFILLER_0_262 vpwr vgnd scs8hd_fill_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

