magic
tech sky130A
magscale 1 2
timestamp 1606426090
<< locali >>
rect 8401 13175 8435 13481
rect 4445 12223 4479 12325
rect 7389 12087 7423 12393
rect 10793 12087 10827 12257
rect 10517 11543 10551 11645
rect 4077 11135 4111 11305
rect 7389 11067 7423 11169
rect 12173 10455 12207 10761
rect 13369 10455 13403 10557
rect 12173 9435 12207 9605
rect 7297 9027 7331 9129
rect 13185 8891 13219 9129
rect 3893 6851 3927 6953
rect 7205 6783 7239 6953
rect 13369 6783 13403 6953
rect 6561 6103 6595 6409
rect 10609 6171 10643 6273
rect 12173 6239 12207 6341
rect 6929 5763 6963 5865
rect 6561 4471 6595 4709
rect 5273 3519 5307 3621
rect 11529 3519 11563 3621
rect 12173 3383 12207 3485
rect 15393 3043 15427 3145
rect 5273 2499 5307 2601
<< viali >>
rect 15853 14501 15887 14535
rect 16773 14501 16807 14535
rect 4537 14433 4571 14467
rect 10149 14433 10183 14467
rect 14968 14433 15002 14467
rect 17417 14433 17451 14467
rect 4629 14365 4663 14399
rect 4721 14365 4755 14399
rect 10241 14365 10275 14399
rect 10333 14365 10367 14399
rect 15761 14365 15795 14399
rect 17509 14365 17543 14399
rect 17693 14365 17727 14399
rect 4169 14229 4203 14263
rect 9781 14229 9815 14263
rect 15071 14229 15105 14263
rect 17049 14229 17083 14263
rect 3893 14025 3927 14059
rect 9137 14025 9171 14059
rect 2881 13957 2915 13991
rect 10241 13957 10275 13991
rect 13553 13957 13587 13991
rect 18245 13957 18279 13991
rect 3433 13889 3467 13923
rect 4537 13889 4571 13923
rect 5365 13889 5399 13923
rect 5457 13889 5491 13923
rect 7481 13889 7515 13923
rect 9781 13889 9815 13923
rect 10701 13889 10735 13923
rect 10885 13889 10919 13923
rect 11621 13889 11655 13923
rect 13185 13889 13219 13923
rect 14197 13889 14231 13923
rect 15301 13889 15335 13923
rect 15485 13889 15519 13923
rect 15945 13889 15979 13923
rect 16957 13889 16991 13923
rect 3341 13821 3375 13855
rect 7205 13821 7239 13855
rect 7297 13821 7331 13855
rect 9505 13821 9539 13855
rect 11345 13821 11379 13855
rect 12449 13821 12483 13855
rect 12817 13821 12851 13855
rect 14013 13821 14047 13855
rect 15209 13821 15243 13855
rect 17233 13821 17267 13855
rect 18061 13821 18095 13855
rect 4261 13753 4295 13787
rect 16037 13753 16071 13787
rect 3249 13685 3283 13719
rect 4353 13685 4387 13719
rect 4905 13685 4939 13719
rect 5273 13685 5307 13719
rect 6837 13685 6871 13719
rect 9597 13685 9631 13719
rect 10609 13685 10643 13719
rect 13921 13685 13955 13719
rect 14841 13685 14875 13719
rect 17417 13685 17451 13719
rect 1961 13481 1995 13515
rect 2513 13481 2547 13515
rect 2881 13481 2915 13515
rect 4813 13481 4847 13515
rect 6377 13481 6411 13515
rect 8309 13481 8343 13515
rect 8401 13481 8435 13515
rect 10057 13481 10091 13515
rect 10701 13481 10735 13515
rect 11069 13481 11103 13515
rect 13277 13481 13311 13515
rect 13553 13481 13587 13515
rect 15301 13481 15335 13515
rect 17969 13481 18003 13515
rect 7196 13413 7230 13447
rect 1869 13345 1903 13379
rect 2973 13345 3007 13379
rect 5181 13345 5215 13379
rect 5273 13345 5307 13379
rect 6285 13345 6319 13379
rect 2145 13277 2179 13311
rect 3065 13277 3099 13311
rect 5457 13277 5491 13311
rect 6561 13277 6595 13311
rect 6929 13277 6963 13311
rect 8953 13345 8987 13379
rect 10149 13345 10183 13379
rect 12164 13345 12198 13379
rect 13921 13345 13955 13379
rect 15669 13345 15703 13379
rect 16681 13345 16715 13379
rect 17877 13345 17911 13379
rect 9045 13277 9079 13311
rect 9137 13277 9171 13311
rect 10241 13277 10275 13311
rect 11161 13277 11195 13311
rect 11345 13277 11379 13311
rect 11897 13277 11931 13311
rect 14013 13277 14047 13311
rect 14105 13277 14139 13311
rect 15761 13277 15795 13311
rect 15853 13277 15887 13311
rect 16773 13277 16807 13311
rect 16865 13277 16899 13311
rect 18061 13277 18095 13311
rect 8585 13209 8619 13243
rect 1501 13141 1535 13175
rect 5917 13141 5951 13175
rect 8401 13141 8435 13175
rect 9689 13141 9723 13175
rect 16313 13141 16347 13175
rect 17509 13141 17543 13175
rect 1777 12937 1811 12971
rect 4169 12937 4203 12971
rect 6193 12937 6227 12971
rect 8217 12937 8251 12971
rect 10241 12937 10275 12971
rect 11989 12937 12023 12971
rect 15945 12937 15979 12971
rect 16957 12937 16991 12971
rect 13829 12869 13863 12903
rect 2329 12801 2363 12835
rect 16497 12801 16531 12835
rect 17601 12801 17635 12835
rect 2789 12733 2823 12767
rect 4813 12733 4847 12767
rect 5080 12733 5114 12767
rect 6837 12733 6871 12767
rect 7104 12733 7138 12767
rect 8861 12733 8895 12767
rect 10609 12733 10643 12767
rect 12449 12733 12483 12767
rect 14289 12733 14323 12767
rect 17325 12733 17359 12767
rect 2237 12665 2271 12699
rect 3056 12665 3090 12699
rect 9128 12665 9162 12699
rect 10854 12665 10888 12699
rect 12716 12665 12750 12699
rect 14534 12665 14568 12699
rect 16313 12665 16347 12699
rect 2145 12597 2179 12631
rect 15669 12597 15703 12631
rect 16405 12597 16439 12631
rect 17417 12597 17451 12631
rect 2973 12393 3007 12427
rect 3341 12393 3375 12427
rect 4537 12393 4571 12427
rect 4997 12393 5031 12427
rect 5549 12393 5583 12427
rect 6929 12393 6963 12427
rect 7389 12393 7423 12427
rect 7573 12393 7607 12427
rect 8585 12393 8619 12427
rect 9965 12393 9999 12427
rect 11437 12393 11471 12427
rect 13921 12393 13955 12427
rect 15669 12393 15703 12427
rect 16129 12393 16163 12427
rect 3433 12325 3467 12359
rect 4445 12325 4479 12359
rect 2329 12257 2363 12291
rect 4905 12257 4939 12291
rect 5917 12257 5951 12291
rect 2421 12189 2455 12223
rect 2605 12189 2639 12223
rect 3617 12189 3651 12223
rect 4445 12189 4479 12223
rect 5089 12189 5123 12223
rect 6009 12189 6043 12223
rect 6193 12189 6227 12223
rect 7021 12189 7055 12223
rect 7205 12189 7239 12223
rect 1961 12121 1995 12155
rect 14289 12325 14323 12359
rect 16037 12325 16071 12359
rect 16948 12325 16982 12359
rect 7941 12257 7975 12291
rect 8953 12257 8987 12291
rect 10333 12257 10367 12291
rect 10793 12257 10827 12291
rect 11345 12257 11379 12291
rect 12357 12257 12391 12291
rect 16681 12257 16715 12291
rect 8033 12189 8067 12223
rect 8217 12189 8251 12223
rect 9045 12189 9079 12223
rect 9229 12189 9263 12223
rect 10425 12189 10459 12223
rect 10517 12189 10551 12223
rect 6561 12053 6595 12087
rect 7389 12053 7423 12087
rect 11529 12189 11563 12223
rect 12449 12189 12483 12223
rect 12633 12189 12667 12223
rect 13461 12189 13495 12223
rect 14381 12189 14415 12223
rect 14565 12189 14599 12223
rect 16221 12189 16255 12223
rect 10793 12053 10827 12087
rect 10977 12053 11011 12087
rect 11989 12053 12023 12087
rect 18061 12053 18095 12087
rect 2605 11849 2639 11883
rect 5733 11849 5767 11883
rect 8953 11849 8987 11883
rect 12541 11849 12575 11883
rect 13829 11849 13863 11883
rect 16957 11849 16991 11883
rect 1593 11781 1627 11815
rect 10701 11781 10735 11815
rect 16681 11781 16715 11815
rect 2237 11713 2271 11747
rect 3249 11713 3283 11747
rect 5273 11713 5307 11747
rect 6377 11713 6411 11747
rect 9229 11713 9263 11747
rect 10333 11713 10367 11747
rect 11161 11713 11195 11747
rect 11345 11713 11379 11747
rect 13093 11713 13127 11747
rect 14473 11713 14507 11747
rect 15301 11713 15335 11747
rect 17509 11713 17543 11747
rect 3617 11645 3651 11679
rect 3884 11645 3918 11679
rect 7573 11645 7607 11679
rect 7840 11645 7874 11679
rect 10517 11645 10551 11679
rect 14197 11645 14231 11679
rect 15568 11645 15602 11679
rect 1961 11577 1995 11611
rect 2973 11577 3007 11611
rect 6193 11577 6227 11611
rect 11069 11577 11103 11611
rect 12909 11577 12943 11611
rect 17325 11577 17359 11611
rect 2053 11509 2087 11543
rect 3065 11509 3099 11543
rect 4997 11509 5031 11543
rect 6101 11509 6135 11543
rect 9689 11509 9723 11543
rect 10057 11509 10091 11543
rect 10149 11509 10183 11543
rect 10517 11509 10551 11543
rect 13001 11509 13035 11543
rect 14289 11509 14323 11543
rect 17417 11509 17451 11543
rect 3709 11305 3743 11339
rect 4077 11305 4111 11339
rect 6837 11305 6871 11339
rect 11069 11305 11103 11339
rect 13645 11305 13679 11339
rect 13921 11305 13955 11339
rect 14381 11305 14415 11339
rect 16681 11305 16715 11339
rect 2596 11237 2630 11271
rect 1685 11169 1719 11203
rect 9934 11237 9968 11271
rect 12532 11237 12566 11271
rect 15568 11237 15602 11271
rect 4528 11169 4562 11203
rect 6101 11169 6135 11203
rect 7389 11169 7423 11203
rect 7665 11169 7699 11203
rect 8208 11169 8242 11203
rect 9689 11169 9723 11203
rect 11621 11169 11655 11203
rect 14289 11169 14323 11203
rect 15117 11169 15151 11203
rect 15301 11169 15335 11203
rect 17325 11169 17359 11203
rect 2329 11101 2363 11135
rect 4077 11101 4111 11135
rect 4261 11101 4295 11135
rect 6929 11101 6963 11135
rect 7113 11101 7147 11135
rect 7941 11101 7975 11135
rect 12265 11101 12299 11135
rect 14473 11101 14507 11135
rect 17417 11101 17451 11135
rect 17601 11101 17635 11135
rect 1869 11033 1903 11067
rect 5917 11033 5951 11067
rect 6469 11033 6503 11067
rect 7389 11033 7423 11067
rect 9321 11033 9355 11067
rect 14933 11033 14967 11067
rect 16957 11033 16991 11067
rect 5641 10965 5675 10999
rect 7481 10965 7515 10999
rect 11437 10965 11471 10999
rect 3709 10761 3743 10795
rect 9137 10761 9171 10795
rect 12173 10761 12207 10795
rect 4721 10693 4755 10727
rect 12081 10693 12115 10727
rect 4261 10625 4295 10659
rect 5365 10625 5399 10659
rect 6285 10625 6319 10659
rect 7757 10625 7791 10659
rect 9873 10625 9907 10659
rect 9965 10625 9999 10659
rect 10701 10625 10735 10659
rect 1409 10557 1443 10591
rect 1676 10557 1710 10591
rect 3065 10557 3099 10591
rect 6193 10557 6227 10591
rect 9781 10557 9815 10591
rect 6101 10489 6135 10523
rect 8024 10489 8058 10523
rect 10968 10489 11002 10523
rect 15301 10693 15335 10727
rect 13093 10625 13127 10659
rect 15945 10625 15979 10659
rect 18061 10625 18095 10659
rect 13369 10557 13403 10591
rect 13461 10557 13495 10591
rect 13728 10557 13762 10591
rect 15761 10557 15795 10591
rect 16313 10557 16347 10591
rect 16580 10557 16614 10591
rect 12909 10489 12943 10523
rect 15669 10489 15703 10523
rect 2789 10421 2823 10455
rect 3249 10421 3283 10455
rect 4077 10421 4111 10455
rect 4169 10421 4203 10455
rect 5089 10421 5123 10455
rect 5181 10421 5215 10455
rect 5733 10421 5767 10455
rect 9413 10421 9447 10455
rect 12173 10421 12207 10455
rect 12449 10421 12483 10455
rect 12817 10421 12851 10455
rect 13369 10421 13403 10455
rect 14841 10421 14875 10455
rect 17693 10421 17727 10455
rect 2237 10217 2271 10251
rect 2973 10217 3007 10251
rect 4629 10217 4663 10251
rect 4905 10217 4939 10251
rect 5273 10217 5307 10251
rect 11989 10217 12023 10251
rect 12265 10217 12299 10251
rect 13277 10217 13311 10251
rect 13737 10217 13771 10251
rect 14289 10217 14323 10251
rect 15761 10217 15795 10251
rect 18337 10217 18371 10251
rect 1409 10149 1443 10183
rect 9956 10149 9990 10183
rect 13645 10149 13679 10183
rect 15669 10149 15703 10183
rect 2329 10081 2363 10115
rect 3341 10081 3375 10115
rect 3433 10081 3467 10115
rect 4077 10081 4111 10115
rect 4813 10081 4847 10115
rect 5917 10081 5951 10115
rect 6184 10081 6218 10115
rect 8033 10081 8067 10115
rect 9689 10081 9723 10115
rect 12173 10081 12207 10115
rect 12633 10081 12667 10115
rect 16957 10081 16991 10115
rect 17224 10081 17258 10115
rect 2513 10013 2547 10047
rect 3525 10013 3559 10047
rect 5365 10013 5399 10047
rect 5457 10013 5491 10047
rect 8125 10013 8159 10047
rect 8217 10013 8251 10047
rect 8677 10013 8711 10047
rect 12725 10013 12759 10047
rect 12817 10013 12851 10047
rect 13921 10013 13955 10047
rect 15899 10013 15933 10047
rect 7297 9945 7331 9979
rect 1869 9877 1903 9911
rect 4261 9877 4295 9911
rect 7665 9877 7699 9911
rect 11069 9877 11103 9911
rect 15301 9877 15335 9911
rect 3709 9605 3743 9639
rect 5733 9605 5767 9639
rect 9321 9605 9355 9639
rect 10149 9605 10183 9639
rect 12173 9605 12207 9639
rect 13829 9605 13863 9639
rect 4353 9537 4387 9571
rect 5365 9537 5399 9571
rect 6377 9537 6411 9571
rect 7297 9537 7331 9571
rect 7481 9537 7515 9571
rect 8217 9537 8251 9571
rect 9045 9537 9079 9571
rect 9781 9537 9815 9571
rect 9873 9537 9907 9571
rect 10701 9537 10735 9571
rect 11897 9537 11931 9571
rect 1501 9469 1535 9503
rect 2053 9469 2087 9503
rect 4077 9469 4111 9503
rect 8033 9469 8067 9503
rect 8861 9469 8895 9503
rect 8953 9469 8987 9503
rect 10517 9469 10551 9503
rect 14197 9537 14231 9571
rect 17049 9537 17083 9571
rect 12449 9469 12483 9503
rect 14464 9469 14498 9503
rect 16773 9469 16807 9503
rect 2320 9401 2354 9435
rect 5181 9401 5215 9435
rect 6101 9401 6135 9435
rect 9689 9401 9723 9435
rect 11713 9401 11747 9435
rect 12173 9401 12207 9435
rect 12716 9401 12750 9435
rect 1685 9333 1719 9367
rect 3433 9333 3467 9367
rect 4169 9333 4203 9367
rect 4721 9333 4755 9367
rect 5089 9333 5123 9367
rect 6193 9333 6227 9367
rect 6837 9333 6871 9367
rect 7205 9333 7239 9367
rect 7665 9333 7699 9367
rect 8125 9333 8159 9367
rect 8493 9333 8527 9367
rect 10609 9333 10643 9367
rect 11345 9333 11379 9367
rect 11805 9333 11839 9367
rect 15577 9333 15611 9367
rect 16405 9333 16439 9367
rect 16865 9333 16899 9367
rect 7297 9129 7331 9163
rect 8769 9129 8803 9163
rect 10057 9129 10091 9163
rect 11805 9129 11839 9163
rect 12357 9129 12391 9163
rect 12725 9129 12759 9163
rect 13185 9129 13219 9163
rect 14657 9129 14691 9163
rect 17509 9129 17543 9163
rect 2421 9061 2455 9095
rect 5978 9061 6012 9095
rect 7634 9061 7668 9095
rect 10149 9061 10183 9095
rect 11713 9061 11747 9095
rect 12817 9061 12851 9095
rect 1409 8993 1443 9027
rect 2329 8993 2363 9027
rect 3341 8993 3375 9027
rect 4333 8993 4367 9027
rect 5733 8993 5767 9027
rect 7297 8993 7331 9027
rect 7389 8993 7423 9027
rect 10885 8993 10919 9027
rect 2513 8925 2547 8959
rect 3433 8925 3467 8959
rect 3525 8925 3559 8959
rect 4077 8925 4111 8959
rect 10333 8925 10367 8959
rect 10977 8925 11011 8959
rect 11161 8925 11195 8959
rect 11989 8925 12023 8959
rect 12909 8925 12943 8959
rect 14565 8993 14599 9027
rect 16129 8993 16163 9027
rect 16396 8993 16430 9027
rect 13369 8925 13403 8959
rect 14841 8925 14875 8959
rect 15301 8925 15335 8959
rect 1593 8857 1627 8891
rect 7113 8857 7147 8891
rect 9689 8857 9723 8891
rect 10517 8857 10551 8891
rect 11345 8857 11379 8891
rect 13185 8857 13219 8891
rect 1961 8789 1995 8823
rect 2973 8789 3007 8823
rect 5457 8789 5491 8823
rect 14197 8789 14231 8823
rect 6285 8585 6319 8619
rect 10517 8585 10551 8619
rect 12449 8585 12483 8619
rect 17233 8585 17267 8619
rect 2789 8517 2823 8551
rect 3065 8517 3099 8551
rect 4261 8517 4295 8551
rect 7021 8517 7055 8551
rect 11161 8517 11195 8551
rect 13553 8517 13587 8551
rect 18245 8517 18279 8551
rect 1409 8449 1443 8483
rect 3525 8449 3559 8483
rect 3709 8449 3743 8483
rect 11713 8449 11747 8483
rect 13001 8449 13035 8483
rect 14013 8449 14047 8483
rect 14197 8449 14231 8483
rect 15117 8449 15151 8483
rect 15853 8449 15887 8483
rect 1676 8381 1710 8415
rect 4077 8381 4111 8415
rect 4905 8381 4939 8415
rect 7181 8381 7215 8415
rect 7573 8381 7607 8415
rect 7840 8381 7874 8415
rect 11529 8381 11563 8415
rect 18061 8381 18095 8415
rect 5172 8313 5206 8347
rect 9229 8313 9263 8347
rect 11621 8313 11655 8347
rect 12909 8313 12943 8347
rect 13921 8313 13955 8347
rect 15025 8313 15059 8347
rect 16098 8313 16132 8347
rect 3433 8245 3467 8279
rect 8953 8245 8987 8279
rect 12817 8245 12851 8279
rect 14565 8245 14599 8279
rect 14933 8245 14967 8279
rect 2329 8041 2363 8075
rect 4077 8041 4111 8075
rect 4445 8041 4479 8075
rect 5089 8041 5123 8075
rect 6101 8041 6135 8075
rect 6469 8041 6503 8075
rect 7665 8041 7699 8075
rect 8677 8041 8711 8075
rect 12725 8041 12759 8075
rect 13369 8041 13403 8075
rect 14657 8041 14691 8075
rect 16681 8041 16715 8075
rect 16957 8041 16991 8075
rect 17325 8041 17359 8075
rect 3249 7973 3283 8007
rect 5457 7973 5491 8007
rect 8033 7973 8067 8007
rect 10057 7973 10091 8007
rect 11612 7973 11646 8007
rect 14565 7973 14599 8007
rect 2237 7905 2271 7939
rect 3341 7905 3375 7939
rect 7113 7905 7147 7939
rect 8125 7905 8159 7939
rect 10149 7905 10183 7939
rect 11345 7905 11379 7939
rect 15557 7905 15591 7939
rect 17969 7905 18003 7939
rect 2421 7837 2455 7871
rect 3525 7837 3559 7871
rect 4537 7837 4571 7871
rect 4721 7837 4755 7871
rect 5549 7837 5583 7871
rect 5733 7837 5767 7871
rect 6561 7837 6595 7871
rect 6745 7837 6779 7871
rect 8217 7837 8251 7871
rect 10241 7837 10275 7871
rect 10701 7837 10735 7871
rect 13461 7837 13495 7871
rect 13553 7837 13587 7871
rect 14841 7837 14875 7871
rect 15301 7837 15335 7871
rect 17417 7837 17451 7871
rect 17509 7837 17543 7871
rect 2881 7769 2915 7803
rect 18153 7769 18187 7803
rect 1869 7701 1903 7735
rect 7297 7701 7331 7735
rect 9689 7701 9723 7735
rect 13001 7701 13035 7735
rect 14197 7701 14231 7735
rect 3709 7497 3743 7531
rect 6377 7497 6411 7531
rect 7113 7497 7147 7531
rect 11713 7497 11747 7531
rect 11989 7497 12023 7531
rect 16589 7497 16623 7531
rect 13461 7429 13495 7463
rect 18245 7429 18279 7463
rect 4353 7361 4387 7395
rect 4997 7361 5031 7395
rect 7665 7361 7699 7395
rect 10333 7361 10367 7395
rect 12909 7361 12943 7395
rect 13093 7361 13127 7395
rect 13921 7361 13955 7395
rect 14013 7361 14047 7395
rect 15117 7361 15151 7395
rect 16037 7361 16071 7395
rect 16221 7361 16255 7395
rect 17049 7361 17083 7395
rect 17233 7361 17267 7395
rect 1593 7293 1627 7327
rect 1860 7293 1894 7327
rect 4905 7293 4939 7327
rect 7481 7293 7515 7327
rect 7573 7293 7607 7327
rect 8493 7293 8527 7327
rect 8760 7293 8794 7327
rect 12173 7293 12207 7327
rect 14933 7293 14967 7327
rect 16957 7293 16991 7327
rect 18061 7293 18095 7327
rect 3249 7225 3283 7259
rect 4077 7225 4111 7259
rect 4169 7225 4203 7259
rect 5264 7225 5298 7259
rect 10600 7225 10634 7259
rect 13829 7225 13863 7259
rect 15945 7225 15979 7259
rect 2973 7157 3007 7191
rect 4721 7157 4755 7191
rect 9873 7157 9907 7191
rect 12449 7157 12483 7191
rect 12817 7157 12851 7191
rect 14565 7157 14599 7191
rect 15025 7157 15059 7191
rect 15577 7157 15611 7191
rect 3893 6953 3927 6987
rect 6377 6953 6411 6987
rect 7205 6953 7239 6987
rect 8769 6953 8803 6987
rect 13369 6953 13403 6987
rect 14933 6953 14967 6987
rect 15669 6953 15703 6987
rect 6745 6885 6779 6919
rect 1685 6817 1719 6851
rect 2329 6817 2363 6851
rect 2596 6817 2630 6851
rect 3893 6817 3927 6851
rect 4084 6817 4118 6851
rect 4344 6817 4378 6851
rect 5733 6817 5767 6851
rect 7389 6817 7423 6851
rect 7656 6817 7690 6851
rect 9781 6817 9815 6851
rect 10048 6817 10082 6851
rect 11897 6817 11931 6851
rect 12909 6817 12943 6851
rect 16681 6885 16715 6919
rect 13553 6817 13587 6851
rect 13820 6817 13854 6851
rect 15761 6817 15795 6851
rect 17877 6817 17911 6851
rect 6837 6749 6871 6783
rect 7021 6749 7055 6783
rect 7205 6749 7239 6783
rect 9045 6749 9079 6783
rect 11989 6749 12023 6783
rect 12173 6749 12207 6783
rect 13001 6749 13035 6783
rect 13185 6749 13219 6783
rect 13369 6749 13403 6783
rect 15945 6749 15979 6783
rect 16773 6749 16807 6783
rect 16865 6749 16899 6783
rect 3709 6681 3743 6715
rect 5917 6681 5951 6715
rect 11529 6681 11563 6715
rect 12541 6681 12575 6715
rect 18061 6681 18095 6715
rect 1869 6613 1903 6647
rect 5457 6613 5491 6647
rect 11161 6613 11195 6647
rect 15301 6613 15335 6647
rect 16313 6613 16347 6647
rect 6561 6409 6595 6443
rect 8217 6409 8251 6443
rect 10793 6409 10827 6443
rect 11345 6409 11379 6443
rect 13553 6409 13587 6443
rect 18245 6409 18279 6443
rect 5733 6341 5767 6375
rect 2697 6273 2731 6307
rect 2881 6273 2915 6307
rect 4353 6273 4387 6307
rect 5273 6273 5307 6307
rect 6377 6273 6411 6307
rect 1685 6205 1719 6239
rect 2605 6205 2639 6239
rect 3249 6205 3283 6239
rect 4077 6137 4111 6171
rect 6193 6137 6227 6171
rect 10517 6341 10551 6375
rect 12173 6341 12207 6375
rect 15577 6341 15611 6375
rect 10609 6273 10643 6307
rect 11897 6273 11931 6307
rect 6837 6205 6871 6239
rect 9137 6205 9171 6239
rect 13185 6273 13219 6307
rect 14197 6273 14231 6307
rect 15117 6273 15151 6307
rect 16129 6273 16163 6307
rect 10977 6205 11011 6239
rect 12173 6205 12207 6239
rect 13921 6205 13955 6239
rect 17417 6205 17451 6239
rect 18061 6205 18095 6239
rect 7082 6137 7116 6171
rect 9404 6137 9438 6171
rect 10609 6137 10643 6171
rect 11713 6137 11747 6171
rect 1869 6069 1903 6103
rect 2237 6069 2271 6103
rect 3709 6069 3743 6103
rect 4169 6069 4203 6103
rect 4721 6069 4755 6103
rect 5089 6069 5123 6103
rect 5181 6069 5215 6103
rect 6101 6069 6135 6103
rect 6561 6069 6595 6103
rect 8493 6069 8527 6103
rect 11805 6069 11839 6103
rect 12541 6069 12575 6103
rect 12909 6069 12943 6103
rect 13001 6069 13035 6103
rect 14013 6069 14047 6103
rect 14565 6069 14599 6103
rect 14933 6069 14967 6103
rect 15025 6069 15059 6103
rect 15945 6069 15979 6103
rect 16037 6069 16071 6103
rect 17601 6069 17635 6103
rect 4077 5865 4111 5899
rect 6837 5865 6871 5899
rect 6929 5865 6963 5899
rect 9321 5865 9355 5899
rect 11897 5865 11931 5899
rect 14197 5865 14231 5899
rect 18061 5865 18095 5899
rect 1860 5797 1894 5831
rect 4537 5797 4571 5831
rect 14657 5797 14691 5831
rect 3249 5729 3283 5763
rect 4445 5729 4479 5763
rect 5273 5729 5307 5763
rect 5457 5729 5491 5763
rect 5724 5729 5758 5763
rect 6929 5729 6963 5763
rect 7113 5729 7147 5763
rect 7841 5729 7875 5763
rect 8208 5729 8242 5763
rect 9965 5729 9999 5763
rect 10232 5729 10266 5763
rect 12081 5729 12115 5763
rect 12440 5729 12474 5763
rect 14013 5729 14047 5763
rect 14565 5729 14599 5763
rect 15301 5729 15335 5763
rect 17325 5729 17359 5763
rect 17877 5729 17911 5763
rect 1593 5661 1627 5695
rect 4629 5661 4663 5695
rect 7941 5661 7975 5695
rect 12173 5661 12207 5695
rect 14841 5661 14875 5695
rect 13553 5593 13587 5627
rect 2973 5525 3007 5559
rect 3433 5525 3467 5559
rect 5089 5525 5123 5559
rect 7297 5525 7331 5559
rect 7665 5525 7699 5559
rect 11345 5525 11379 5559
rect 13829 5525 13863 5559
rect 17509 5525 17543 5559
rect 6193 5321 6227 5355
rect 8861 5321 8895 5355
rect 9873 5321 9907 5355
rect 10885 5321 10919 5355
rect 13829 5321 13863 5355
rect 15761 5321 15795 5355
rect 3985 5253 4019 5287
rect 4537 5185 4571 5219
rect 5549 5185 5583 5219
rect 7297 5185 7331 5219
rect 7389 5185 7423 5219
rect 8309 5185 8343 5219
rect 8493 5185 8527 5219
rect 9413 5185 9447 5219
rect 10425 5185 10459 5219
rect 11437 5185 11471 5219
rect 12449 5185 12483 5219
rect 14105 5185 14139 5219
rect 16313 5185 16347 5219
rect 1409 5117 1443 5151
rect 3065 5117 3099 5151
rect 5365 5117 5399 5151
rect 5457 5117 5491 5151
rect 6009 5117 6043 5151
rect 11253 5117 11287 5151
rect 17417 5117 17451 5151
rect 18061 5117 18095 5151
rect 1676 5049 1710 5083
rect 7205 5049 7239 5083
rect 9321 5049 9355 5083
rect 11345 5049 11379 5083
rect 12716 5049 12750 5083
rect 14372 5049 14406 5083
rect 16129 5049 16163 5083
rect 2789 4981 2823 5015
rect 3249 4981 3283 5015
rect 4353 4981 4387 5015
rect 4445 4981 4479 5015
rect 4997 4981 5031 5015
rect 6837 4981 6871 5015
rect 7849 4981 7883 5015
rect 8217 4981 8251 5015
rect 9229 4981 9263 5015
rect 10241 4981 10275 5015
rect 10333 4981 10367 5015
rect 11897 4981 11931 5015
rect 15485 4981 15519 5015
rect 16221 4981 16255 5015
rect 17601 4981 17635 5015
rect 18245 4981 18279 5015
rect 6101 4777 6135 4811
rect 9229 4777 9263 4811
rect 11805 4777 11839 4811
rect 11897 4777 11931 4811
rect 13185 4777 13219 4811
rect 13737 4777 13771 4811
rect 14105 4777 14139 4811
rect 15301 4777 15335 4811
rect 15669 4777 15703 4811
rect 2320 4709 2354 4743
rect 6561 4709 6595 4743
rect 13093 4709 13127 4743
rect 1501 4641 1535 4675
rect 4077 4641 4111 4675
rect 4344 4641 4378 4675
rect 6193 4641 6227 4675
rect 2053 4573 2087 4607
rect 6285 4573 6319 4607
rect 7113 4641 7147 4675
rect 7205 4641 7239 4675
rect 8116 4641 8150 4675
rect 9781 4641 9815 4675
rect 10048 4641 10082 4675
rect 17325 4641 17359 4675
rect 17877 4641 17911 4675
rect 7297 4573 7331 4607
rect 7849 4573 7883 4607
rect 11989 4573 12023 4607
rect 13369 4573 13403 4607
rect 14197 4573 14231 4607
rect 14381 4573 14415 4607
rect 15761 4573 15795 4607
rect 15945 4573 15979 4607
rect 1685 4437 1719 4471
rect 3433 4437 3467 4471
rect 5457 4437 5491 4471
rect 5733 4437 5767 4471
rect 6561 4437 6595 4471
rect 6745 4437 6779 4471
rect 11161 4437 11195 4471
rect 11437 4437 11471 4471
rect 12725 4437 12759 4471
rect 17509 4437 17543 4471
rect 18061 4437 18095 4471
rect 4077 4233 4111 4267
rect 15025 4233 15059 4267
rect 2329 4097 2363 4131
rect 2697 4097 2731 4131
rect 5549 4097 5583 4131
rect 8125 4097 8159 4131
rect 8309 4097 8343 4131
rect 9229 4097 9263 4131
rect 10241 4097 10275 4131
rect 10701 4097 10735 4131
rect 13001 4097 13035 4131
rect 13185 4097 13219 4131
rect 2053 4029 2087 4063
rect 4353 4029 4387 4063
rect 5365 4029 5399 4063
rect 6009 4029 6043 4063
rect 6837 4029 6871 4063
rect 8033 4029 8067 4063
rect 10149 4029 10183 4063
rect 13645 4029 13679 4063
rect 17417 4029 17451 4063
rect 18061 4029 18095 4063
rect 2964 3961 2998 3995
rect 6285 3961 6319 3995
rect 7113 3961 7147 3995
rect 9045 3961 9079 3995
rect 10057 3961 10091 3995
rect 10968 3961 11002 3995
rect 13912 3961 13946 3995
rect 1685 3893 1719 3927
rect 2145 3893 2179 3927
rect 4537 3893 4571 3927
rect 4997 3893 5031 3927
rect 5457 3893 5491 3927
rect 7665 3893 7699 3927
rect 8677 3893 8711 3927
rect 9137 3893 9171 3927
rect 9689 3893 9723 3927
rect 12081 3893 12115 3927
rect 12541 3893 12575 3927
rect 12909 3893 12943 3927
rect 17601 3893 17635 3927
rect 18245 3893 18279 3927
rect 2513 3689 2547 3723
rect 2973 3689 3007 3723
rect 4905 3689 4939 3723
rect 13921 3689 13955 3723
rect 14381 3689 14415 3723
rect 5273 3621 5307 3655
rect 5702 3621 5736 3655
rect 10057 3621 10091 3655
rect 11529 3621 11563 3655
rect 12510 3621 12544 3655
rect 1593 3553 1627 3587
rect 2329 3553 2363 3587
rect 3341 3553 3375 3587
rect 4813 3553 4847 3587
rect 7369 3553 7403 3587
rect 8769 3553 8803 3587
rect 10149 3553 10183 3587
rect 11069 3553 11103 3587
rect 11713 3553 11747 3587
rect 12265 3553 12299 3587
rect 14289 3553 14323 3587
rect 15301 3553 15335 3587
rect 17325 3553 17359 3587
rect 17877 3553 17911 3587
rect 1777 3485 1811 3519
rect 3433 3485 3467 3519
rect 3617 3485 3651 3519
rect 5089 3485 5123 3519
rect 5273 3485 5307 3519
rect 5457 3485 5491 3519
rect 7113 3485 7147 3519
rect 8953 3485 8987 3519
rect 10241 3485 10275 3519
rect 11161 3485 11195 3519
rect 11345 3485 11379 3519
rect 11529 3485 11563 3519
rect 12173 3485 12207 3519
rect 14473 3485 14507 3519
rect 15485 3485 15519 3519
rect 13645 3417 13679 3451
rect 4445 3349 4479 3383
rect 6837 3349 6871 3383
rect 8493 3349 8527 3383
rect 9689 3349 9723 3383
rect 10701 3349 10735 3383
rect 11897 3349 11931 3383
rect 12173 3349 12207 3383
rect 17509 3349 17543 3383
rect 18061 3349 18095 3383
rect 3157 3145 3191 3179
rect 5549 3145 5583 3179
rect 8125 3145 8159 3179
rect 9137 3145 9171 3179
rect 10149 3145 10183 3179
rect 15393 3145 15427 3179
rect 4537 3077 4571 3111
rect 12449 3077 12483 3111
rect 1869 3009 1903 3043
rect 3709 3009 3743 3043
rect 4997 3009 5031 3043
rect 5181 3009 5215 3043
rect 6101 3009 6135 3043
rect 8677 3009 8711 3043
rect 9597 3009 9631 3043
rect 9689 3009 9723 3043
rect 10609 3009 10643 3043
rect 10793 3009 10827 3043
rect 11621 3009 11655 3043
rect 11713 3009 11747 3043
rect 13001 3009 13035 3043
rect 14933 3009 14967 3043
rect 15393 3009 15427 3043
rect 15669 3009 15703 3043
rect 1593 2941 1627 2975
rect 2329 2941 2363 2975
rect 3525 2941 3559 2975
rect 3617 2941 3651 2975
rect 4905 2941 4939 2975
rect 6837 2941 6871 2975
rect 9505 2941 9539 2975
rect 10517 2941 10551 2975
rect 14013 2941 14047 2975
rect 14749 2941 14783 2975
rect 15516 2941 15550 2975
rect 16221 2941 16255 2975
rect 16865 2941 16899 2975
rect 17417 2941 17451 2975
rect 18061 2941 18095 2975
rect 2605 2873 2639 2907
rect 7665 2873 7699 2907
rect 11529 2873 11563 2907
rect 12817 2873 12851 2907
rect 14289 2873 14323 2907
rect 5917 2805 5951 2839
rect 6009 2805 6043 2839
rect 8493 2805 8527 2839
rect 8585 2805 8619 2839
rect 11161 2805 11195 2839
rect 12909 2805 12943 2839
rect 16405 2805 16439 2839
rect 17049 2805 17083 2839
rect 17601 2805 17635 2839
rect 18245 2805 18279 2839
rect 1869 2601 1903 2635
rect 3341 2601 3375 2635
rect 3433 2601 3467 2635
rect 4905 2601 4939 2635
rect 5273 2601 5307 2635
rect 6377 2601 6411 2635
rect 9045 2601 9079 2635
rect 10241 2601 10275 2635
rect 10701 2601 10735 2635
rect 11713 2601 11747 2635
rect 4813 2533 4847 2567
rect 11621 2533 11655 2567
rect 12909 2533 12943 2567
rect 1685 2465 1719 2499
rect 2237 2465 2271 2499
rect 5273 2465 5307 2499
rect 5457 2465 5491 2499
rect 6193 2465 6227 2499
rect 6929 2465 6963 2499
rect 7757 2465 7791 2499
rect 10609 2465 10643 2499
rect 12633 2465 12667 2499
rect 13369 2465 13403 2499
rect 14105 2465 14139 2499
rect 17417 2465 17451 2499
rect 2513 2397 2547 2431
rect 3617 2397 3651 2431
rect 4997 2397 5031 2431
rect 5641 2397 5675 2431
rect 7113 2397 7147 2431
rect 7941 2397 7975 2431
rect 9137 2397 9171 2431
rect 9321 2397 9355 2431
rect 10885 2397 10919 2431
rect 11805 2397 11839 2431
rect 13553 2397 13587 2431
rect 14289 2397 14323 2431
rect 2973 2329 3007 2363
rect 11253 2329 11287 2363
rect 4445 2261 4479 2295
rect 8677 2261 8711 2295
rect 17601 2261 17635 2295
<< metal1 >>
rect 4062 15172 4068 15224
rect 4120 15212 4126 15224
rect 9490 15212 9496 15224
rect 4120 15184 9496 15212
rect 4120 15172 4126 15184
rect 9490 15172 9496 15184
rect 9548 15172 9554 15224
rect 1104 14714 18860 14736
rect 1104 14662 6912 14714
rect 6964 14662 6976 14714
rect 7028 14662 7040 14714
rect 7092 14662 7104 14714
rect 7156 14662 12843 14714
rect 12895 14662 12907 14714
rect 12959 14662 12971 14714
rect 13023 14662 13035 14714
rect 13087 14662 18860 14714
rect 1104 14640 18860 14662
rect 3418 14560 3424 14612
rect 3476 14600 3482 14612
rect 11146 14600 11152 14612
rect 3476 14572 11152 14600
rect 3476 14560 3482 14572
rect 11146 14560 11152 14572
rect 11204 14560 11210 14612
rect 5350 14492 5356 14544
rect 5408 14532 5414 14544
rect 14274 14532 14280 14544
rect 5408 14504 14280 14532
rect 5408 14492 5414 14504
rect 14274 14492 14280 14504
rect 14332 14492 14338 14544
rect 15841 14535 15899 14541
rect 15841 14532 15853 14535
rect 15212 14504 15853 14532
rect 4522 14464 4528 14476
rect 4483 14436 4528 14464
rect 4522 14424 4528 14436
rect 4580 14424 4586 14476
rect 10042 14424 10048 14476
rect 10100 14424 10106 14476
rect 10137 14467 10195 14473
rect 10137 14433 10149 14467
rect 10183 14464 10195 14467
rect 10410 14464 10416 14476
rect 10183 14436 10416 14464
rect 10183 14433 10195 14436
rect 10137 14427 10195 14433
rect 10410 14424 10416 14436
rect 10468 14424 10474 14476
rect 13906 14424 13912 14476
rect 13964 14464 13970 14476
rect 14366 14464 14372 14476
rect 13964 14436 14372 14464
rect 13964 14424 13970 14436
rect 14366 14424 14372 14436
rect 14424 14464 14430 14476
rect 14956 14467 15014 14473
rect 14956 14464 14968 14467
rect 14424 14436 14968 14464
rect 14424 14424 14430 14436
rect 14956 14433 14968 14436
rect 15002 14464 15014 14467
rect 15212 14464 15240 14504
rect 15841 14501 15853 14504
rect 15887 14501 15899 14535
rect 15841 14495 15899 14501
rect 16761 14535 16819 14541
rect 16761 14501 16773 14535
rect 16807 14532 16819 14535
rect 18782 14532 18788 14544
rect 16807 14504 18788 14532
rect 16807 14501 16819 14504
rect 16761 14495 16819 14501
rect 18782 14492 18788 14504
rect 18840 14492 18846 14544
rect 17402 14464 17408 14476
rect 15002 14436 15240 14464
rect 17363 14436 17408 14464
rect 15002 14433 15014 14436
rect 14956 14427 15014 14433
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 3050 14356 3056 14408
rect 3108 14396 3114 14408
rect 4617 14399 4675 14405
rect 4617 14396 4629 14399
rect 3108 14368 4629 14396
rect 3108 14356 3114 14368
rect 4617 14365 4629 14368
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 4706 14356 4712 14408
rect 4764 14396 4770 14408
rect 10060 14396 10088 14424
rect 10229 14399 10287 14405
rect 10229 14396 10241 14399
rect 4764 14368 4809 14396
rect 10060 14368 10241 14396
rect 4764 14356 4770 14368
rect 10229 14365 10241 14368
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14396 10379 14399
rect 10502 14396 10508 14408
rect 10367 14368 10508 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 10502 14356 10508 14368
rect 10560 14396 10566 14408
rect 11054 14396 11060 14408
rect 10560 14368 11060 14396
rect 10560 14356 10566 14368
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 15378 14356 15384 14408
rect 15436 14396 15442 14408
rect 15749 14399 15807 14405
rect 15749 14396 15761 14399
rect 15436 14368 15761 14396
rect 15436 14356 15442 14368
rect 15749 14365 15761 14368
rect 15795 14365 15807 14399
rect 17494 14396 17500 14408
rect 17455 14368 17500 14396
rect 15749 14359 15807 14365
rect 17494 14356 17500 14368
rect 17552 14356 17558 14408
rect 17678 14396 17684 14408
rect 17639 14368 17684 14396
rect 17678 14356 17684 14368
rect 17736 14356 17742 14408
rect 3326 14288 3332 14340
rect 3384 14328 3390 14340
rect 18046 14328 18052 14340
rect 3384 14300 18052 14328
rect 3384 14288 3390 14300
rect 18046 14288 18052 14300
rect 18104 14288 18110 14340
rect 4157 14263 4215 14269
rect 4157 14229 4169 14263
rect 4203 14260 4215 14263
rect 9674 14260 9680 14272
rect 4203 14232 9680 14260
rect 4203 14229 4215 14232
rect 4157 14223 4215 14229
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 9769 14263 9827 14269
rect 9769 14229 9781 14263
rect 9815 14260 9827 14263
rect 10778 14260 10784 14272
rect 9815 14232 10784 14260
rect 9815 14229 9827 14232
rect 9769 14223 9827 14229
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 15059 14263 15117 14269
rect 15059 14229 15071 14263
rect 15105 14260 15117 14263
rect 15654 14260 15660 14272
rect 15105 14232 15660 14260
rect 15105 14229 15117 14232
rect 15059 14223 15117 14229
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 17034 14260 17040 14272
rect 16995 14232 17040 14260
rect 17034 14220 17040 14232
rect 17092 14220 17098 14272
rect 1104 14170 18860 14192
rect 1104 14118 3947 14170
rect 3999 14118 4011 14170
rect 4063 14118 4075 14170
rect 4127 14118 4139 14170
rect 4191 14118 9878 14170
rect 9930 14118 9942 14170
rect 9994 14118 10006 14170
rect 10058 14118 10070 14170
rect 10122 14118 15808 14170
rect 15860 14118 15872 14170
rect 15924 14118 15936 14170
rect 15988 14118 16000 14170
rect 16052 14118 18860 14170
rect 1104 14096 18860 14118
rect 3881 14059 3939 14065
rect 3881 14025 3893 14059
rect 3927 14056 3939 14059
rect 4522 14056 4528 14068
rect 3927 14028 4528 14056
rect 3927 14025 3939 14028
rect 3881 14019 3939 14025
rect 4522 14016 4528 14028
rect 4580 14016 4586 14068
rect 9125 14059 9183 14065
rect 9125 14025 9137 14059
rect 9171 14056 9183 14059
rect 10686 14056 10692 14068
rect 9171 14028 10692 14056
rect 9171 14025 9183 14028
rect 9125 14019 9183 14025
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 13446 14056 13452 14068
rect 10796 14028 13452 14056
rect 2869 13991 2927 13997
rect 2869 13957 2881 13991
rect 2915 13988 2927 13991
rect 2958 13988 2964 14000
rect 2915 13960 2964 13988
rect 2915 13957 2927 13960
rect 2869 13951 2927 13957
rect 2958 13948 2964 13960
rect 3016 13948 3022 14000
rect 3602 13948 3608 14000
rect 3660 13988 3666 14000
rect 10229 13991 10287 13997
rect 3660 13960 9536 13988
rect 3660 13948 3666 13960
rect 2682 13880 2688 13932
rect 2740 13920 2746 13932
rect 3421 13923 3479 13929
rect 3421 13920 3433 13923
rect 2740 13892 3433 13920
rect 2740 13880 2746 13892
rect 3421 13889 3433 13892
rect 3467 13889 3479 13923
rect 3421 13883 3479 13889
rect 4525 13923 4583 13929
rect 4525 13889 4537 13923
rect 4571 13920 4583 13923
rect 4798 13920 4804 13932
rect 4571 13892 4804 13920
rect 4571 13889 4583 13892
rect 4525 13883 4583 13889
rect 4798 13880 4804 13892
rect 4856 13880 4862 13932
rect 5350 13920 5356 13932
rect 5311 13892 5356 13920
rect 5350 13880 5356 13892
rect 5408 13880 5414 13932
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 7466 13920 7472 13932
rect 5500 13892 5545 13920
rect 7427 13892 7472 13920
rect 5500 13880 5506 13892
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 2774 13812 2780 13864
rect 2832 13852 2838 13864
rect 3329 13855 3387 13861
rect 3329 13852 3341 13855
rect 2832 13824 3341 13852
rect 2832 13812 2838 13824
rect 3329 13821 3341 13824
rect 3375 13821 3387 13855
rect 3329 13815 3387 13821
rect 6638 13812 6644 13864
rect 6696 13852 6702 13864
rect 7193 13855 7251 13861
rect 7193 13852 7205 13855
rect 6696 13824 7205 13852
rect 6696 13812 6702 13824
rect 7193 13821 7205 13824
rect 7239 13821 7251 13855
rect 7193 13815 7251 13821
rect 7285 13855 7343 13861
rect 7285 13821 7297 13855
rect 7331 13852 7343 13855
rect 8110 13852 8116 13864
rect 7331 13824 8116 13852
rect 7331 13821 7343 13824
rect 7285 13815 7343 13821
rect 8110 13812 8116 13824
rect 8168 13812 8174 13864
rect 9508 13861 9536 13960
rect 10229 13957 10241 13991
rect 10275 13988 10287 13991
rect 10594 13988 10600 14000
rect 10275 13960 10600 13988
rect 10275 13957 10287 13960
rect 10229 13951 10287 13957
rect 10594 13948 10600 13960
rect 10652 13948 10658 14000
rect 9769 13923 9827 13929
rect 9769 13889 9781 13923
rect 9815 13920 9827 13923
rect 10502 13920 10508 13932
rect 9815 13892 10508 13920
rect 9815 13889 9827 13892
rect 9769 13883 9827 13889
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13920 10747 13923
rect 10796 13920 10824 14028
rect 13446 14016 13452 14028
rect 13504 14056 13510 14068
rect 16206 14056 16212 14068
rect 13504 14028 16212 14056
rect 13504 14016 13510 14028
rect 16206 14016 16212 14028
rect 16264 14016 16270 14068
rect 13541 13991 13599 13997
rect 13541 13957 13553 13991
rect 13587 13988 13599 13991
rect 14734 13988 14740 14000
rect 13587 13960 14740 13988
rect 13587 13957 13599 13960
rect 13541 13951 13599 13957
rect 14734 13948 14740 13960
rect 14792 13948 14798 14000
rect 14918 13948 14924 14000
rect 14976 13988 14982 14000
rect 17126 13988 17132 14000
rect 14976 13960 15332 13988
rect 14976 13948 14982 13960
rect 10735 13892 10824 13920
rect 10873 13923 10931 13929
rect 10735 13889 10747 13892
rect 10689 13883 10747 13889
rect 10873 13889 10885 13923
rect 10919 13920 10931 13923
rect 11054 13920 11060 13932
rect 10919 13892 11060 13920
rect 10919 13889 10931 13892
rect 10873 13883 10931 13889
rect 11054 13880 11060 13892
rect 11112 13880 11118 13932
rect 11609 13923 11667 13929
rect 11609 13889 11621 13923
rect 11655 13920 11667 13923
rect 12158 13920 12164 13932
rect 11655 13892 12164 13920
rect 11655 13889 11667 13892
rect 11609 13883 11667 13889
rect 12158 13880 12164 13892
rect 12216 13880 12222 13932
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13920 13231 13923
rect 13906 13920 13912 13932
rect 13219 13892 13912 13920
rect 13219 13889 13231 13892
rect 13173 13883 13231 13889
rect 13906 13880 13912 13892
rect 13964 13880 13970 13932
rect 14182 13920 14188 13932
rect 14143 13892 14188 13920
rect 14182 13880 14188 13892
rect 14240 13880 14246 13932
rect 15304 13929 15332 13960
rect 15488 13960 17132 13988
rect 15488 13929 15516 13960
rect 17126 13948 17132 13960
rect 17184 13988 17190 14000
rect 17678 13988 17684 14000
rect 17184 13960 17684 13988
rect 17184 13948 17190 13960
rect 17678 13948 17684 13960
rect 17736 13948 17742 14000
rect 18233 13991 18291 13997
rect 18233 13957 18245 13991
rect 18279 13988 18291 13991
rect 18506 13988 18512 14000
rect 18279 13960 18512 13988
rect 18279 13957 18291 13960
rect 18233 13951 18291 13957
rect 18506 13948 18512 13960
rect 18564 13948 18570 14000
rect 15289 13923 15347 13929
rect 15289 13889 15301 13923
rect 15335 13889 15347 13923
rect 15289 13883 15347 13889
rect 15473 13923 15531 13929
rect 15473 13889 15485 13923
rect 15519 13889 15531 13923
rect 15473 13883 15531 13889
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13920 15991 13923
rect 16574 13920 16580 13932
rect 15979 13892 16580 13920
rect 15979 13889 15991 13892
rect 15933 13883 15991 13889
rect 16574 13880 16580 13892
rect 16632 13880 16638 13932
rect 16945 13923 17003 13929
rect 16945 13889 16957 13923
rect 16991 13920 17003 13923
rect 17586 13920 17592 13932
rect 16991 13892 17592 13920
rect 16991 13889 17003 13892
rect 16945 13883 17003 13889
rect 17586 13880 17592 13892
rect 17644 13880 17650 13932
rect 9493 13855 9551 13861
rect 9493 13821 9505 13855
rect 9539 13852 9551 13855
rect 9582 13852 9588 13864
rect 9539 13824 9588 13852
rect 9539 13821 9551 13824
rect 9493 13815 9551 13821
rect 9582 13812 9588 13824
rect 9640 13812 9646 13864
rect 9674 13812 9680 13864
rect 9732 13852 9738 13864
rect 11333 13855 11391 13861
rect 11333 13852 11345 13855
rect 9732 13824 11345 13852
rect 9732 13812 9738 13824
rect 11333 13821 11345 13824
rect 11379 13821 11391 13855
rect 11333 13815 11391 13821
rect 12434 13812 12440 13864
rect 12492 13852 12498 13864
rect 12805 13855 12863 13861
rect 12492 13824 12537 13852
rect 12492 13812 12498 13824
rect 12805 13821 12817 13855
rect 12851 13852 12863 13855
rect 13262 13852 13268 13864
rect 12851 13824 13268 13852
rect 12851 13821 12863 13824
rect 12805 13815 12863 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 14001 13855 14059 13861
rect 14001 13821 14013 13855
rect 14047 13852 14059 13855
rect 14047 13824 15148 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 4249 13787 4307 13793
rect 4249 13753 4261 13787
rect 4295 13784 4307 13787
rect 4295 13756 4936 13784
rect 4295 13753 4307 13756
rect 4249 13747 4307 13753
rect 1946 13676 1952 13728
rect 2004 13716 2010 13728
rect 3237 13719 3295 13725
rect 3237 13716 3249 13719
rect 2004 13688 3249 13716
rect 2004 13676 2010 13688
rect 3237 13685 3249 13688
rect 3283 13685 3295 13719
rect 3237 13679 3295 13685
rect 4338 13676 4344 13728
rect 4396 13716 4402 13728
rect 4908 13725 4936 13756
rect 5534 13744 5540 13796
rect 5592 13784 5598 13796
rect 10134 13784 10140 13796
rect 5592 13756 7144 13784
rect 5592 13744 5598 13756
rect 4893 13719 4951 13725
rect 4396 13688 4441 13716
rect 4396 13676 4402 13688
rect 4893 13685 4905 13719
rect 4939 13685 4951 13719
rect 5258 13716 5264 13728
rect 5219 13688 5264 13716
rect 4893 13679 4951 13685
rect 5258 13676 5264 13688
rect 5316 13676 5322 13728
rect 6362 13676 6368 13728
rect 6420 13716 6426 13728
rect 6825 13719 6883 13725
rect 6825 13716 6837 13719
rect 6420 13688 6837 13716
rect 6420 13676 6426 13688
rect 6825 13685 6837 13688
rect 6871 13685 6883 13719
rect 7116 13716 7144 13756
rect 9048 13756 10140 13784
rect 9048 13716 9076 13756
rect 10134 13744 10140 13756
rect 10192 13744 10198 13796
rect 10318 13744 10324 13796
rect 10376 13784 10382 13796
rect 10376 13756 11192 13784
rect 10376 13744 10382 13756
rect 7116 13688 9076 13716
rect 9585 13719 9643 13725
rect 6825 13679 6883 13685
rect 9585 13685 9597 13719
rect 9631 13716 9643 13719
rect 10502 13716 10508 13728
rect 9631 13688 10508 13716
rect 9631 13685 9643 13688
rect 9585 13679 9643 13685
rect 10502 13676 10508 13688
rect 10560 13676 10566 13728
rect 10597 13719 10655 13725
rect 10597 13685 10609 13719
rect 10643 13716 10655 13719
rect 10686 13716 10692 13728
rect 10643 13688 10692 13716
rect 10643 13685 10655 13688
rect 10597 13679 10655 13685
rect 10686 13676 10692 13688
rect 10744 13676 10750 13728
rect 11164 13716 11192 13756
rect 11238 13744 11244 13796
rect 11296 13784 11302 13796
rect 15120 13784 15148 13824
rect 15194 13812 15200 13864
rect 15252 13852 15258 13864
rect 15252 13824 15297 13852
rect 15252 13812 15258 13824
rect 15654 13812 15660 13864
rect 15712 13852 15718 13864
rect 17218 13852 17224 13864
rect 15712 13824 15792 13852
rect 17179 13824 17224 13852
rect 15712 13812 15718 13824
rect 15286 13784 15292 13796
rect 11296 13756 14964 13784
rect 15120 13756 15292 13784
rect 11296 13744 11302 13756
rect 13262 13716 13268 13728
rect 11164 13688 13268 13716
rect 13262 13676 13268 13688
rect 13320 13676 13326 13728
rect 13906 13716 13912 13728
rect 13867 13688 13912 13716
rect 13906 13676 13912 13688
rect 13964 13676 13970 13728
rect 14826 13716 14832 13728
rect 14787 13688 14832 13716
rect 14826 13676 14832 13688
rect 14884 13676 14890 13728
rect 14936 13716 14964 13756
rect 15286 13744 15292 13756
rect 15344 13744 15350 13796
rect 15764 13784 15792 13824
rect 17218 13812 17224 13824
rect 17276 13812 17282 13864
rect 18046 13852 18052 13864
rect 18007 13824 18052 13852
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 16025 13787 16083 13793
rect 16025 13784 16037 13787
rect 15764 13756 16037 13784
rect 16025 13753 16037 13756
rect 16071 13753 16083 13787
rect 16025 13747 16083 13753
rect 17405 13719 17463 13725
rect 17405 13716 17417 13719
rect 14936 13688 17417 13716
rect 17405 13685 17417 13688
rect 17451 13685 17463 13719
rect 17405 13679 17463 13685
rect 1104 13626 18860 13648
rect 1104 13574 6912 13626
rect 6964 13574 6976 13626
rect 7028 13574 7040 13626
rect 7092 13574 7104 13626
rect 7156 13574 12843 13626
rect 12895 13574 12907 13626
rect 12959 13574 12971 13626
rect 13023 13574 13035 13626
rect 13087 13574 18860 13626
rect 1104 13552 18860 13574
rect 1949 13515 2007 13521
rect 1949 13481 1961 13515
rect 1995 13512 2007 13515
rect 2501 13515 2559 13521
rect 2501 13512 2513 13515
rect 1995 13484 2513 13512
rect 1995 13481 2007 13484
rect 1949 13475 2007 13481
rect 2501 13481 2513 13484
rect 2547 13481 2559 13515
rect 2866 13512 2872 13524
rect 2779 13484 2872 13512
rect 2501 13475 2559 13481
rect 2866 13472 2872 13484
rect 2924 13512 2930 13524
rect 4062 13512 4068 13524
rect 2924 13484 4068 13512
rect 2924 13472 2930 13484
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 4338 13472 4344 13524
rect 4396 13512 4402 13524
rect 4801 13515 4859 13521
rect 4801 13512 4813 13515
rect 4396 13484 4813 13512
rect 4396 13472 4402 13484
rect 4801 13481 4813 13484
rect 4847 13481 4859 13515
rect 6362 13512 6368 13524
rect 6323 13484 6368 13512
rect 4801 13475 4859 13481
rect 6362 13472 6368 13484
rect 6420 13472 6426 13524
rect 7466 13472 7472 13524
rect 7524 13512 7530 13524
rect 8297 13515 8355 13521
rect 8297 13512 8309 13515
rect 7524 13484 8309 13512
rect 7524 13472 7530 13484
rect 8297 13481 8309 13484
rect 8343 13481 8355 13515
rect 8297 13475 8355 13481
rect 8389 13515 8447 13521
rect 8389 13481 8401 13515
rect 8435 13512 8447 13515
rect 9950 13512 9956 13524
rect 8435 13484 9956 13512
rect 8435 13481 8447 13484
rect 8389 13475 8447 13481
rect 9950 13472 9956 13484
rect 10008 13472 10014 13524
rect 10045 13515 10103 13521
rect 10045 13481 10057 13515
rect 10091 13512 10103 13515
rect 10689 13515 10747 13521
rect 10689 13512 10701 13515
rect 10091 13484 10701 13512
rect 10091 13481 10103 13484
rect 10045 13475 10103 13481
rect 10689 13481 10701 13484
rect 10735 13481 10747 13515
rect 10689 13475 10747 13481
rect 11057 13515 11115 13521
rect 11057 13481 11069 13515
rect 11103 13512 11115 13515
rect 11146 13512 11152 13524
rect 11103 13484 11152 13512
rect 11103 13481 11115 13484
rect 11057 13475 11115 13481
rect 11146 13472 11152 13484
rect 11204 13512 11210 13524
rect 11514 13512 11520 13524
rect 11204 13484 11520 13512
rect 11204 13472 11210 13484
rect 11514 13472 11520 13484
rect 11572 13472 11578 13524
rect 13262 13512 13268 13524
rect 13223 13484 13268 13512
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 13541 13515 13599 13521
rect 13541 13481 13553 13515
rect 13587 13512 13599 13515
rect 13906 13512 13912 13524
rect 13587 13484 13912 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 13906 13472 13912 13484
rect 13964 13472 13970 13524
rect 15286 13512 15292 13524
rect 15247 13484 15292 13512
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 17954 13512 17960 13524
rect 17915 13484 17960 13512
rect 17954 13472 17960 13484
rect 18012 13472 18018 13524
rect 7184 13447 7242 13453
rect 2884 13416 6408 13444
rect 1762 13336 1768 13388
rect 1820 13376 1826 13388
rect 1857 13379 1915 13385
rect 1857 13376 1869 13379
rect 1820 13348 1869 13376
rect 1820 13336 1826 13348
rect 1857 13345 1869 13348
rect 1903 13345 1915 13379
rect 2884 13376 2912 13416
rect 1857 13339 1915 13345
rect 2056 13348 2912 13376
rect 2961 13379 3019 13385
rect 1118 13268 1124 13320
rect 1176 13308 1182 13320
rect 2056 13308 2084 13348
rect 2961 13345 2973 13379
rect 3007 13376 3019 13379
rect 3142 13376 3148 13388
rect 3007 13348 3148 13376
rect 3007 13345 3019 13348
rect 2961 13339 3019 13345
rect 3142 13336 3148 13348
rect 3200 13336 3206 13388
rect 3786 13336 3792 13388
rect 3844 13376 3850 13388
rect 5169 13379 5227 13385
rect 5169 13376 5181 13379
rect 3844 13348 5181 13376
rect 3844 13336 3850 13348
rect 5169 13345 5181 13348
rect 5215 13345 5227 13379
rect 5169 13339 5227 13345
rect 5261 13379 5319 13385
rect 5261 13345 5273 13379
rect 5307 13376 5319 13379
rect 5350 13376 5356 13388
rect 5307 13348 5356 13376
rect 5307 13345 5319 13348
rect 5261 13339 5319 13345
rect 1176 13280 2084 13308
rect 2133 13311 2191 13317
rect 1176 13268 1182 13280
rect 2133 13277 2145 13311
rect 2179 13308 2191 13311
rect 2682 13308 2688 13320
rect 2179 13280 2688 13308
rect 2179 13277 2191 13280
rect 2133 13271 2191 13277
rect 2682 13268 2688 13280
rect 2740 13268 2746 13320
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13277 3111 13311
rect 3053 13271 3111 13277
rect 2038 13200 2044 13252
rect 2096 13240 2102 13252
rect 3068 13240 3096 13271
rect 2096 13212 3096 13240
rect 5184 13240 5212 13339
rect 5350 13336 5356 13348
rect 5408 13336 5414 13388
rect 6270 13376 6276 13388
rect 6231 13348 6276 13376
rect 6270 13336 6276 13348
rect 6328 13336 6334 13388
rect 6380 13376 6408 13416
rect 7184 13413 7196 13447
rect 7230 13444 7242 13447
rect 7742 13444 7748 13456
rect 7230 13416 7748 13444
rect 7230 13413 7242 13416
rect 7184 13407 7242 13413
rect 7742 13404 7748 13416
rect 7800 13404 7806 13456
rect 12434 13444 12440 13456
rect 7852 13416 12440 13444
rect 7852 13376 7880 13416
rect 12434 13404 12440 13416
rect 12492 13404 12498 13456
rect 14108 13416 15884 13444
rect 6380 13348 7880 13376
rect 8294 13336 8300 13388
rect 8352 13376 8358 13388
rect 8941 13379 8999 13385
rect 8941 13376 8953 13379
rect 8352 13348 8953 13376
rect 8352 13336 8358 13348
rect 8941 13345 8953 13348
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13376 10195 13379
rect 10686 13376 10692 13388
rect 10183 13348 10692 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 10686 13336 10692 13348
rect 10744 13336 10750 13388
rect 12152 13379 12210 13385
rect 12152 13345 12164 13379
rect 12198 13376 12210 13379
rect 13906 13376 13912 13388
rect 12198 13348 13492 13376
rect 13867 13348 13912 13376
rect 12198 13345 12210 13348
rect 12152 13339 12210 13345
rect 5442 13308 5448 13320
rect 5355 13280 5448 13308
rect 5442 13268 5448 13280
rect 5500 13308 5506 13320
rect 6546 13308 6552 13320
rect 5500 13280 6552 13308
rect 5500 13268 5506 13280
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 6914 13308 6920 13320
rect 6875 13280 6920 13308
rect 6914 13268 6920 13280
rect 6972 13268 6978 13320
rect 9030 13308 9036 13320
rect 8991 13280 9036 13308
rect 9030 13268 9036 13280
rect 9088 13268 9094 13320
rect 9122 13268 9128 13320
rect 9180 13308 9186 13320
rect 10229 13311 10287 13317
rect 10229 13308 10241 13311
rect 9180 13280 10241 13308
rect 9180 13268 9186 13280
rect 10229 13277 10241 13280
rect 10275 13277 10287 13311
rect 11146 13308 11152 13320
rect 11107 13280 11152 13308
rect 10229 13271 10287 13277
rect 11146 13268 11152 13280
rect 11204 13268 11210 13320
rect 11330 13308 11336 13320
rect 11291 13280 11336 13308
rect 11330 13268 11336 13280
rect 11388 13268 11394 13320
rect 11882 13308 11888 13320
rect 11843 13280 11888 13308
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 8573 13243 8631 13249
rect 5184 13212 6040 13240
rect 2096 13200 2102 13212
rect 1489 13175 1547 13181
rect 1489 13141 1501 13175
rect 1535 13172 1547 13175
rect 2222 13172 2228 13184
rect 1535 13144 2228 13172
rect 1535 13141 1547 13144
rect 1489 13135 1547 13141
rect 2222 13132 2228 13144
rect 2280 13132 2286 13184
rect 4338 13132 4344 13184
rect 4396 13172 4402 13184
rect 5905 13175 5963 13181
rect 5905 13172 5917 13175
rect 4396 13144 5917 13172
rect 4396 13132 4402 13144
rect 5905 13141 5917 13144
rect 5951 13141 5963 13175
rect 6012 13172 6040 13212
rect 8573 13209 8585 13243
rect 8619 13240 8631 13243
rect 9766 13240 9772 13252
rect 8619 13212 9772 13240
rect 8619 13209 8631 13212
rect 8573 13203 8631 13209
rect 9766 13200 9772 13212
rect 9824 13200 9830 13252
rect 9858 13200 9864 13252
rect 9916 13200 9922 13252
rect 9950 13200 9956 13252
rect 10008 13240 10014 13252
rect 11698 13240 11704 13252
rect 10008 13212 11704 13240
rect 10008 13200 10014 13212
rect 11698 13200 11704 13212
rect 11756 13200 11762 13252
rect 13464 13240 13492 13348
rect 13906 13336 13912 13348
rect 13964 13336 13970 13388
rect 14108 13320 14136 13416
rect 15562 13336 15568 13388
rect 15620 13376 15626 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15620 13348 15669 13376
rect 15620 13336 15626 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 13998 13308 14004 13320
rect 13959 13280 14004 13308
rect 13998 13268 14004 13280
rect 14056 13268 14062 13320
rect 14090 13268 14096 13320
rect 14148 13308 14154 13320
rect 15856 13317 15884 13416
rect 16669 13379 16727 13385
rect 16669 13345 16681 13379
rect 16715 13376 16727 13379
rect 16942 13376 16948 13388
rect 16715 13348 16948 13376
rect 16715 13345 16727 13348
rect 16669 13339 16727 13345
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 17862 13376 17868 13388
rect 17823 13348 17868 13376
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 15749 13311 15807 13317
rect 15749 13308 15761 13311
rect 14148 13280 14193 13308
rect 15672 13280 15761 13308
rect 14148 13268 14154 13280
rect 15672 13252 15700 13280
rect 15749 13277 15761 13280
rect 15795 13277 15807 13311
rect 15749 13271 15807 13277
rect 15841 13311 15899 13317
rect 15841 13277 15853 13311
rect 15887 13277 15899 13311
rect 16758 13308 16764 13320
rect 16719 13280 16764 13308
rect 15841 13271 15899 13277
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 16850 13268 16856 13320
rect 16908 13308 16914 13320
rect 18049 13311 18107 13317
rect 16908 13280 16953 13308
rect 16908 13268 16914 13280
rect 18049 13277 18061 13311
rect 18095 13277 18107 13311
rect 18049 13271 18107 13277
rect 14182 13240 14188 13252
rect 13464 13212 14188 13240
rect 14182 13200 14188 13212
rect 14240 13200 14246 13252
rect 15654 13200 15660 13252
rect 15712 13200 15718 13252
rect 17678 13200 17684 13252
rect 17736 13240 17742 13252
rect 18064 13240 18092 13271
rect 17736 13212 18092 13240
rect 17736 13200 17742 13212
rect 8389 13175 8447 13181
rect 8389 13172 8401 13175
rect 6012 13144 8401 13172
rect 5905 13135 5963 13141
rect 8389 13141 8401 13144
rect 8435 13141 8447 13175
rect 9674 13172 9680 13184
rect 9635 13144 9680 13172
rect 8389 13135 8447 13141
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 9876 13172 9904 13200
rect 12618 13172 12624 13184
rect 9876 13144 12624 13172
rect 12618 13132 12624 13144
rect 12676 13132 12682 13184
rect 15470 13132 15476 13184
rect 15528 13172 15534 13184
rect 16301 13175 16359 13181
rect 16301 13172 16313 13175
rect 15528 13144 16313 13172
rect 15528 13132 15534 13144
rect 16301 13141 16313 13144
rect 16347 13141 16359 13175
rect 16301 13135 16359 13141
rect 17310 13132 17316 13184
rect 17368 13172 17374 13184
rect 17497 13175 17555 13181
rect 17497 13172 17509 13175
rect 17368 13144 17509 13172
rect 17368 13132 17374 13144
rect 17497 13141 17509 13144
rect 17543 13141 17555 13175
rect 17497 13135 17555 13141
rect 1104 13082 18860 13104
rect 1104 13030 3947 13082
rect 3999 13030 4011 13082
rect 4063 13030 4075 13082
rect 4127 13030 4139 13082
rect 4191 13030 9878 13082
rect 9930 13030 9942 13082
rect 9994 13030 10006 13082
rect 10058 13030 10070 13082
rect 10122 13030 15808 13082
rect 15860 13030 15872 13082
rect 15924 13030 15936 13082
rect 15988 13030 16000 13082
rect 16052 13030 18860 13082
rect 1104 13008 18860 13030
rect 1762 12968 1768 12980
rect 1723 12940 1768 12968
rect 1762 12928 1768 12940
rect 1820 12928 1826 12980
rect 4157 12971 4215 12977
rect 4157 12937 4169 12971
rect 4203 12968 4215 12971
rect 4246 12968 4252 12980
rect 4203 12940 4252 12968
rect 4203 12937 4215 12940
rect 4157 12931 4215 12937
rect 4246 12928 4252 12940
rect 4304 12968 4310 12980
rect 4706 12968 4712 12980
rect 4304 12940 4712 12968
rect 4304 12928 4310 12940
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 4798 12928 4804 12980
rect 4856 12968 4862 12980
rect 6181 12971 6239 12977
rect 6181 12968 6193 12971
rect 4856 12940 6193 12968
rect 4856 12928 4862 12940
rect 6181 12937 6193 12940
rect 6227 12937 6239 12971
rect 6181 12931 6239 12937
rect 6546 12928 6552 12980
rect 6604 12968 6610 12980
rect 8205 12971 8263 12977
rect 8205 12968 8217 12971
rect 6604 12940 8217 12968
rect 6604 12928 6610 12940
rect 8205 12937 8217 12940
rect 8251 12937 8263 12971
rect 8205 12931 8263 12937
rect 9122 12928 9128 12980
rect 9180 12968 9186 12980
rect 10229 12971 10287 12977
rect 10229 12968 10241 12971
rect 9180 12940 10241 12968
rect 9180 12928 9186 12940
rect 10229 12937 10241 12940
rect 10275 12937 10287 12971
rect 11238 12968 11244 12980
rect 10229 12931 10287 12937
rect 10336 12940 11244 12968
rect 2038 12792 2044 12844
rect 2096 12832 2102 12844
rect 2317 12835 2375 12841
rect 2317 12832 2329 12835
rect 2096 12804 2329 12832
rect 2096 12792 2102 12804
rect 2317 12801 2329 12804
rect 2363 12801 2375 12835
rect 2317 12795 2375 12801
rect 7926 12792 7932 12844
rect 7984 12832 7990 12844
rect 7984 12804 8984 12832
rect 7984 12792 7990 12804
rect 2777 12767 2835 12773
rect 2777 12733 2789 12767
rect 2823 12764 2835 12767
rect 4430 12764 4436 12776
rect 2823 12736 4436 12764
rect 2823 12733 2835 12736
rect 2777 12727 2835 12733
rect 4430 12724 4436 12736
rect 4488 12764 4494 12776
rect 5074 12773 5080 12776
rect 4801 12767 4859 12773
rect 4801 12764 4813 12767
rect 4488 12736 4813 12764
rect 4488 12724 4494 12736
rect 4801 12733 4813 12736
rect 4847 12733 4859 12767
rect 5068 12764 5080 12773
rect 4987 12736 5080 12764
rect 4801 12727 4859 12733
rect 5068 12727 5080 12736
rect 5132 12764 5138 12776
rect 5442 12764 5448 12776
rect 5132 12736 5448 12764
rect 5074 12724 5080 12727
rect 5132 12724 5138 12736
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12733 6883 12767
rect 6825 12727 6883 12733
rect 7092 12767 7150 12773
rect 7092 12733 7104 12767
rect 7138 12764 7150 12767
rect 7466 12764 7472 12776
rect 7138 12736 7472 12764
rect 7138 12733 7150 12736
rect 7092 12727 7150 12733
rect 2225 12699 2283 12705
rect 2225 12665 2237 12699
rect 2271 12696 2283 12699
rect 2314 12696 2320 12708
rect 2271 12668 2320 12696
rect 2271 12665 2283 12668
rect 2225 12659 2283 12665
rect 2314 12656 2320 12668
rect 2372 12656 2378 12708
rect 3044 12699 3102 12705
rect 3044 12665 3056 12699
rect 3090 12696 3102 12699
rect 3602 12696 3608 12708
rect 3090 12668 3608 12696
rect 3090 12665 3102 12668
rect 3044 12659 3102 12665
rect 3602 12656 3608 12668
rect 3660 12696 3666 12708
rect 4706 12696 4712 12708
rect 3660 12668 4712 12696
rect 3660 12656 3666 12668
rect 4706 12656 4712 12668
rect 4764 12656 4770 12708
rect 6730 12696 6736 12708
rect 5184 12668 6736 12696
rect 2130 12628 2136 12640
rect 2091 12600 2136 12628
rect 2130 12588 2136 12600
rect 2188 12588 2194 12640
rect 3970 12588 3976 12640
rect 4028 12628 4034 12640
rect 5184 12628 5212 12668
rect 6730 12656 6736 12668
rect 6788 12656 6794 12708
rect 6840 12696 6868 12727
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 7650 12764 7656 12776
rect 7563 12736 7656 12764
rect 6914 12696 6920 12708
rect 6827 12668 6920 12696
rect 6914 12656 6920 12668
rect 6972 12696 6978 12708
rect 7576 12696 7604 12736
rect 7650 12724 7656 12736
rect 7708 12764 7714 12776
rect 8849 12767 8907 12773
rect 8849 12764 8861 12767
rect 7708 12736 8861 12764
rect 7708 12724 7714 12736
rect 8849 12733 8861 12736
rect 8895 12733 8907 12767
rect 8956 12764 8984 12804
rect 10336 12764 10364 12940
rect 11238 12928 11244 12940
rect 11296 12928 11302 12980
rect 11330 12928 11336 12980
rect 11388 12968 11394 12980
rect 11977 12971 12035 12977
rect 11977 12968 11989 12971
rect 11388 12940 11989 12968
rect 11388 12928 11394 12940
rect 11977 12937 11989 12940
rect 12023 12937 12035 12971
rect 11977 12931 12035 12937
rect 15562 12928 15568 12980
rect 15620 12968 15626 12980
rect 15933 12971 15991 12977
rect 15933 12968 15945 12971
rect 15620 12940 15945 12968
rect 15620 12928 15626 12940
rect 15933 12937 15945 12940
rect 15979 12937 15991 12971
rect 16942 12968 16948 12980
rect 16903 12940 16948 12968
rect 15933 12931 15991 12937
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 13817 12903 13875 12909
rect 13817 12869 13829 12903
rect 13863 12900 13875 12903
rect 14182 12900 14188 12912
rect 13863 12872 14188 12900
rect 13863 12869 13875 12872
rect 13817 12863 13875 12869
rect 14182 12860 14188 12872
rect 14240 12860 14246 12912
rect 16482 12832 16488 12844
rect 16443 12804 16488 12832
rect 16482 12792 16488 12804
rect 16540 12792 16546 12844
rect 17589 12835 17647 12841
rect 17589 12801 17601 12835
rect 17635 12832 17647 12835
rect 17770 12832 17776 12844
rect 17635 12804 17776 12832
rect 17635 12801 17647 12804
rect 17589 12795 17647 12801
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 8956 12736 10364 12764
rect 10597 12767 10655 12773
rect 8849 12727 8907 12733
rect 10597 12733 10609 12767
rect 10643 12764 10655 12767
rect 11422 12764 11428 12776
rect 10643 12736 11428 12764
rect 10643 12733 10655 12736
rect 10597 12727 10655 12733
rect 11422 12724 11428 12736
rect 11480 12764 11486 12776
rect 11882 12764 11888 12776
rect 11480 12736 11888 12764
rect 11480 12724 11486 12736
rect 11882 12724 11888 12736
rect 11940 12764 11946 12776
rect 12437 12767 12495 12773
rect 12437 12764 12449 12767
rect 11940 12736 12449 12764
rect 11940 12724 11946 12736
rect 12437 12733 12449 12736
rect 12483 12733 12495 12767
rect 13814 12764 13820 12776
rect 12437 12727 12495 12733
rect 12636 12736 13820 12764
rect 6972 12668 7604 12696
rect 9116 12699 9174 12705
rect 6972 12656 6978 12668
rect 9116 12665 9128 12699
rect 9162 12696 9174 12699
rect 9214 12696 9220 12708
rect 9162 12668 9220 12696
rect 9162 12665 9174 12668
rect 9116 12659 9174 12665
rect 9214 12656 9220 12668
rect 9272 12656 9278 12708
rect 10318 12656 10324 12708
rect 10376 12696 10382 12708
rect 10842 12699 10900 12705
rect 10842 12696 10854 12699
rect 10376 12668 10854 12696
rect 10376 12656 10382 12668
rect 10842 12665 10854 12668
rect 10888 12665 10900 12699
rect 10842 12659 10900 12665
rect 11238 12656 11244 12708
rect 11296 12696 11302 12708
rect 12636 12696 12664 12736
rect 13814 12724 13820 12736
rect 13872 12724 13878 12776
rect 14277 12767 14335 12773
rect 14277 12733 14289 12767
rect 14323 12764 14335 12767
rect 15286 12764 15292 12776
rect 14323 12736 15292 12764
rect 14323 12733 14335 12736
rect 14277 12727 14335 12733
rect 15286 12724 15292 12736
rect 15344 12724 15350 12776
rect 17310 12764 17316 12776
rect 17271 12736 17316 12764
rect 17310 12724 17316 12736
rect 17368 12724 17374 12776
rect 11296 12668 12664 12696
rect 12704 12699 12762 12705
rect 11296 12656 11302 12668
rect 12704 12665 12716 12699
rect 12750 12696 12762 12699
rect 14090 12696 14096 12708
rect 12750 12668 14096 12696
rect 12750 12665 12762 12668
rect 12704 12659 12762 12665
rect 14090 12656 14096 12668
rect 14148 12656 14154 12708
rect 14458 12656 14464 12708
rect 14516 12705 14522 12708
rect 14516 12699 14580 12705
rect 14516 12665 14534 12699
rect 14568 12665 14580 12699
rect 16298 12696 16304 12708
rect 16259 12668 16304 12696
rect 14516 12659 14580 12665
rect 14516 12656 14522 12659
rect 16298 12656 16304 12668
rect 16356 12656 16362 12708
rect 4028 12600 5212 12628
rect 4028 12588 4034 12600
rect 5350 12588 5356 12640
rect 5408 12628 5414 12640
rect 7926 12628 7932 12640
rect 5408 12600 7932 12628
rect 5408 12588 5414 12600
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 8110 12588 8116 12640
rect 8168 12628 8174 12640
rect 11606 12628 11612 12640
rect 8168 12600 11612 12628
rect 8168 12588 8174 12600
rect 11606 12588 11612 12600
rect 11664 12588 11670 12640
rect 14108 12628 14136 12656
rect 15657 12631 15715 12637
rect 15657 12628 15669 12631
rect 14108 12600 15669 12628
rect 15657 12597 15669 12600
rect 15703 12597 15715 12631
rect 16390 12628 16396 12640
rect 16351 12600 16396 12628
rect 15657 12591 15715 12597
rect 16390 12588 16396 12600
rect 16448 12588 16454 12640
rect 16574 12588 16580 12640
rect 16632 12628 16638 12640
rect 17405 12631 17463 12637
rect 17405 12628 17417 12631
rect 16632 12600 17417 12628
rect 16632 12588 16638 12600
rect 17405 12597 17417 12600
rect 17451 12597 17463 12631
rect 17405 12591 17463 12597
rect 1104 12538 18860 12560
rect 1104 12486 6912 12538
rect 6964 12486 6976 12538
rect 7028 12486 7040 12538
rect 7092 12486 7104 12538
rect 7156 12486 12843 12538
rect 12895 12486 12907 12538
rect 12959 12486 12971 12538
rect 13023 12486 13035 12538
rect 13087 12486 18860 12538
rect 1104 12464 18860 12486
rect 2961 12427 3019 12433
rect 2961 12393 2973 12427
rect 3007 12424 3019 12427
rect 3050 12424 3056 12436
rect 3007 12396 3056 12424
rect 3007 12393 3019 12396
rect 2961 12387 3019 12393
rect 3050 12384 3056 12396
rect 3108 12384 3114 12436
rect 3329 12427 3387 12433
rect 3329 12393 3341 12427
rect 3375 12424 3387 12427
rect 4525 12427 4583 12433
rect 4525 12424 4537 12427
rect 3375 12396 4537 12424
rect 3375 12393 3387 12396
rect 3329 12387 3387 12393
rect 4525 12393 4537 12396
rect 4571 12393 4583 12427
rect 4525 12387 4583 12393
rect 4985 12427 5043 12433
rect 4985 12393 4997 12427
rect 5031 12424 5043 12427
rect 5537 12427 5595 12433
rect 5537 12424 5549 12427
rect 5031 12396 5549 12424
rect 5031 12393 5043 12396
rect 4985 12387 5043 12393
rect 5537 12393 5549 12396
rect 5583 12393 5595 12427
rect 6917 12427 6975 12433
rect 6917 12424 6929 12427
rect 5537 12387 5595 12393
rect 5644 12396 6929 12424
rect 3421 12359 3479 12365
rect 3421 12325 3433 12359
rect 3467 12356 3479 12359
rect 4338 12356 4344 12368
rect 3467 12328 4344 12356
rect 3467 12325 3479 12328
rect 3421 12319 3479 12325
rect 4338 12316 4344 12328
rect 4396 12316 4402 12368
rect 4433 12359 4491 12365
rect 4433 12325 4445 12359
rect 4479 12356 4491 12359
rect 4479 12328 4936 12356
rect 4479 12325 4491 12328
rect 4433 12319 4491 12325
rect 4908 12300 4936 12328
rect 5166 12316 5172 12368
rect 5224 12356 5230 12368
rect 5644 12356 5672 12396
rect 6917 12393 6929 12396
rect 6963 12424 6975 12427
rect 7377 12427 7435 12433
rect 7377 12424 7389 12427
rect 6963 12396 7389 12424
rect 6963 12393 6975 12396
rect 6917 12387 6975 12393
rect 7377 12393 7389 12396
rect 7423 12393 7435 12427
rect 7377 12387 7435 12393
rect 7561 12427 7619 12433
rect 7561 12393 7573 12427
rect 7607 12424 7619 12427
rect 8294 12424 8300 12436
rect 7607 12396 8300 12424
rect 7607 12393 7619 12396
rect 7561 12387 7619 12393
rect 8294 12384 8300 12396
rect 8352 12384 8358 12436
rect 8573 12427 8631 12433
rect 8573 12393 8585 12427
rect 8619 12424 8631 12427
rect 9030 12424 9036 12436
rect 8619 12396 9036 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 9953 12427 10011 12433
rect 9953 12393 9965 12427
rect 9999 12424 10011 12427
rect 11146 12424 11152 12436
rect 9999 12396 11152 12424
rect 9999 12393 10011 12396
rect 9953 12387 10011 12393
rect 11146 12384 11152 12396
rect 11204 12384 11210 12436
rect 11330 12384 11336 12436
rect 11388 12384 11394 12436
rect 11425 12427 11483 12433
rect 11425 12393 11437 12427
rect 11471 12424 11483 12427
rect 11606 12424 11612 12436
rect 11471 12396 11612 12424
rect 11471 12393 11483 12396
rect 11425 12387 11483 12393
rect 11606 12384 11612 12396
rect 11664 12424 11670 12436
rect 13262 12424 13268 12436
rect 11664 12396 13268 12424
rect 11664 12384 11670 12396
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 13909 12427 13967 12433
rect 13909 12393 13921 12427
rect 13955 12424 13967 12427
rect 13998 12424 14004 12436
rect 13955 12396 14004 12424
rect 13955 12393 13967 12396
rect 13909 12387 13967 12393
rect 13998 12384 14004 12396
rect 14056 12384 14062 12436
rect 15654 12424 15660 12436
rect 15615 12396 15660 12424
rect 15654 12384 15660 12396
rect 15712 12384 15718 12436
rect 16117 12427 16175 12433
rect 16117 12393 16129 12427
rect 16163 12424 16175 12427
rect 17034 12424 17040 12436
rect 16163 12396 17040 12424
rect 16163 12393 16175 12396
rect 16117 12387 16175 12393
rect 17034 12384 17040 12396
rect 17092 12384 17098 12436
rect 5224 12328 5672 12356
rect 5224 12316 5230 12328
rect 6730 12316 6736 12368
rect 6788 12356 6794 12368
rect 8478 12356 8484 12368
rect 6788 12328 8484 12356
rect 6788 12316 6794 12328
rect 8478 12316 8484 12328
rect 8536 12316 8542 12368
rect 11348 12356 11376 12384
rect 9784 12328 11376 12356
rect 2317 12291 2375 12297
rect 2317 12288 2329 12291
rect 2240 12260 2329 12288
rect 1946 12152 1952 12164
rect 1907 12124 1952 12152
rect 1946 12112 1952 12124
rect 2004 12112 2010 12164
rect 2240 12084 2268 12260
rect 2317 12257 2329 12260
rect 2363 12257 2375 12291
rect 2317 12251 2375 12257
rect 4890 12248 4896 12300
rect 4948 12288 4954 12300
rect 5905 12291 5963 12297
rect 4948 12260 4993 12288
rect 4948 12248 4954 12260
rect 5905 12257 5917 12291
rect 5951 12288 5963 12291
rect 6362 12288 6368 12300
rect 5951 12260 6368 12288
rect 5951 12257 5963 12260
rect 5905 12251 5963 12257
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12288 7987 12291
rect 8846 12288 8852 12300
rect 7975 12260 8852 12288
rect 7975 12257 7987 12260
rect 7929 12251 7987 12257
rect 8846 12248 8852 12260
rect 8904 12248 8910 12300
rect 8941 12291 8999 12297
rect 8941 12257 8953 12291
rect 8987 12288 8999 12291
rect 9398 12288 9404 12300
rect 8987 12260 9404 12288
rect 8987 12257 8999 12260
rect 8941 12251 8999 12257
rect 9398 12248 9404 12260
rect 9456 12248 9462 12300
rect 2406 12220 2412 12232
rect 2367 12192 2412 12220
rect 2406 12180 2412 12192
rect 2464 12180 2470 12232
rect 2590 12180 2596 12232
rect 2648 12220 2654 12232
rect 3602 12220 3608 12232
rect 2648 12192 2693 12220
rect 3563 12192 3608 12220
rect 2648 12180 2654 12192
rect 3602 12180 3608 12192
rect 3660 12180 3666 12232
rect 4154 12180 4160 12232
rect 4212 12220 4218 12232
rect 4433 12223 4491 12229
rect 4433 12220 4445 12223
rect 4212 12192 4445 12220
rect 4212 12180 4218 12192
rect 4433 12189 4445 12192
rect 4479 12189 4491 12223
rect 4433 12183 4491 12189
rect 5074 12180 5080 12232
rect 5132 12220 5138 12232
rect 5132 12192 5177 12220
rect 5132 12180 5138 12192
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 5997 12223 6055 12229
rect 5997 12220 6009 12223
rect 5592 12192 6009 12220
rect 5592 12180 5598 12192
rect 5997 12189 6009 12192
rect 6043 12189 6055 12223
rect 5997 12183 6055 12189
rect 6181 12223 6239 12229
rect 6181 12189 6193 12223
rect 6227 12189 6239 12223
rect 7006 12220 7012 12232
rect 6967 12192 7012 12220
rect 6181 12183 6239 12189
rect 3510 12112 3516 12164
rect 3568 12152 3574 12164
rect 4614 12152 4620 12164
rect 3568 12124 4620 12152
rect 3568 12112 3574 12124
rect 4614 12112 4620 12124
rect 4672 12112 4678 12164
rect 6196 12152 6224 12183
rect 7006 12180 7012 12192
rect 7064 12180 7070 12232
rect 7193 12223 7251 12229
rect 7193 12189 7205 12223
rect 7239 12220 7251 12223
rect 7374 12220 7380 12232
rect 7239 12192 7380 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 7374 12180 7380 12192
rect 7432 12180 7438 12232
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 8021 12223 8079 12229
rect 8021 12220 8033 12223
rect 7616 12192 8033 12220
rect 7616 12180 7622 12192
rect 8021 12189 8033 12192
rect 8067 12220 8079 12223
rect 8110 12220 8116 12232
rect 8067 12192 8116 12220
rect 8067 12189 8079 12192
rect 8021 12183 8079 12189
rect 8110 12180 8116 12192
rect 8168 12180 8174 12232
rect 8205 12223 8263 12229
rect 8205 12189 8217 12223
rect 8251 12189 8263 12223
rect 9030 12220 9036 12232
rect 8991 12192 9036 12220
rect 8205 12183 8263 12189
rect 6914 12152 6920 12164
rect 6196 12124 6920 12152
rect 6914 12112 6920 12124
rect 6972 12152 6978 12164
rect 7466 12152 7472 12164
rect 6972 12124 7472 12152
rect 6972 12112 6978 12124
rect 7466 12112 7472 12124
rect 7524 12112 7530 12164
rect 8220 12152 8248 12183
rect 9030 12180 9036 12192
rect 9088 12180 9094 12232
rect 9214 12220 9220 12232
rect 9127 12192 9220 12220
rect 9214 12180 9220 12192
rect 9272 12220 9278 12232
rect 9784 12220 9812 12328
rect 11698 12316 11704 12368
rect 11756 12356 11762 12368
rect 14090 12356 14096 12368
rect 11756 12328 14096 12356
rect 11756 12316 11762 12328
rect 14090 12316 14096 12328
rect 14148 12356 14154 12368
rect 14277 12359 14335 12365
rect 14277 12356 14289 12359
rect 14148 12328 14289 12356
rect 14148 12316 14154 12328
rect 14277 12325 14289 12328
rect 14323 12325 14335 12359
rect 14277 12319 14335 12325
rect 14826 12316 14832 12368
rect 14884 12356 14890 12368
rect 16025 12359 16083 12365
rect 16025 12356 16037 12359
rect 14884 12328 16037 12356
rect 14884 12316 14890 12328
rect 16025 12325 16037 12328
rect 16071 12325 16083 12359
rect 16025 12319 16083 12325
rect 16936 12359 16994 12365
rect 16936 12325 16948 12359
rect 16982 12356 16994 12359
rect 17126 12356 17132 12368
rect 16982 12328 17132 12356
rect 16982 12325 16994 12328
rect 16936 12319 16994 12325
rect 17126 12316 17132 12328
rect 17184 12316 17190 12368
rect 10321 12291 10379 12297
rect 10321 12257 10333 12291
rect 10367 12288 10379 12291
rect 10781 12291 10839 12297
rect 10367 12260 10732 12288
rect 10367 12257 10379 12260
rect 10321 12251 10379 12257
rect 10413 12223 10471 12229
rect 10413 12220 10425 12223
rect 9272 12192 9812 12220
rect 9876 12192 10425 12220
rect 9272 12180 9278 12192
rect 9232 12152 9260 12180
rect 8220 12124 9260 12152
rect 9306 12112 9312 12164
rect 9364 12152 9370 12164
rect 9876 12152 9904 12192
rect 10413 12189 10425 12192
rect 10459 12189 10471 12223
rect 10413 12183 10471 12189
rect 10505 12223 10563 12229
rect 10505 12189 10517 12223
rect 10551 12189 10563 12223
rect 10505 12183 10563 12189
rect 9364 12124 9904 12152
rect 9364 12112 9370 12124
rect 10318 12112 10324 12164
rect 10376 12152 10382 12164
rect 10520 12152 10548 12183
rect 10376 12124 10548 12152
rect 10704 12152 10732 12260
rect 10781 12257 10793 12291
rect 10827 12288 10839 12291
rect 11333 12291 11391 12297
rect 11333 12288 11345 12291
rect 10827 12260 11345 12288
rect 10827 12257 10839 12260
rect 10781 12251 10839 12257
rect 11333 12257 11345 12260
rect 11379 12288 11391 12291
rect 11974 12288 11980 12300
rect 11379 12260 11980 12288
rect 11379 12257 11391 12260
rect 11333 12251 11391 12257
rect 11974 12248 11980 12260
rect 12032 12248 12038 12300
rect 12342 12288 12348 12300
rect 12303 12260 12348 12288
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 15102 12288 15108 12300
rect 14384 12260 15108 12288
rect 14384 12232 14412 12260
rect 15102 12248 15108 12260
rect 15160 12248 15166 12300
rect 15286 12248 15292 12300
rect 15344 12288 15350 12300
rect 16669 12291 16727 12297
rect 16669 12288 16681 12291
rect 15344 12260 16681 12288
rect 15344 12248 15350 12260
rect 16669 12257 16681 12260
rect 16715 12257 16727 12291
rect 16669 12251 16727 12257
rect 11238 12180 11244 12232
rect 11296 12220 11302 12232
rect 11517 12223 11575 12229
rect 11517 12220 11529 12223
rect 11296 12192 11529 12220
rect 11296 12180 11302 12192
rect 11517 12189 11529 12192
rect 11563 12189 11575 12223
rect 11517 12183 11575 12189
rect 11606 12180 11612 12232
rect 11664 12220 11670 12232
rect 12437 12223 12495 12229
rect 12437 12220 12449 12223
rect 11664 12192 12449 12220
rect 11664 12180 11670 12192
rect 12437 12189 12449 12192
rect 12483 12189 12495 12223
rect 12618 12220 12624 12232
rect 12579 12192 12624 12220
rect 12437 12183 12495 12189
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12220 13507 12223
rect 13722 12220 13728 12232
rect 13495 12192 13728 12220
rect 13495 12189 13507 12192
rect 13449 12183 13507 12189
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 14366 12220 14372 12232
rect 13872 12192 14372 12220
rect 13872 12180 13878 12192
rect 14366 12180 14372 12192
rect 14424 12180 14430 12232
rect 14458 12180 14464 12232
rect 14516 12220 14522 12232
rect 14553 12223 14611 12229
rect 14553 12220 14565 12223
rect 14516 12192 14565 12220
rect 14516 12180 14522 12192
rect 14553 12189 14565 12192
rect 14599 12220 14611 12223
rect 16209 12223 16267 12229
rect 16209 12220 16221 12223
rect 14599 12192 16221 12220
rect 14599 12189 14611 12192
rect 14553 12183 14611 12189
rect 16209 12189 16221 12192
rect 16255 12220 16267 12223
rect 16482 12220 16488 12232
rect 16255 12192 16488 12220
rect 16255 12189 16267 12192
rect 16209 12183 16267 12189
rect 16298 12152 16304 12164
rect 10704 12124 16304 12152
rect 10376 12112 10382 12124
rect 10888 12096 10916 12124
rect 16298 12112 16304 12124
rect 16356 12112 16362 12164
rect 2866 12084 2872 12096
rect 2240 12056 2872 12084
rect 2866 12044 2872 12056
rect 2924 12084 2930 12096
rect 3786 12084 3792 12096
rect 2924 12056 3792 12084
rect 2924 12044 2930 12056
rect 3786 12044 3792 12056
rect 3844 12044 3850 12096
rect 6549 12087 6607 12093
rect 6549 12053 6561 12087
rect 6595 12084 6607 12087
rect 7282 12084 7288 12096
rect 6595 12056 7288 12084
rect 6595 12053 6607 12056
rect 6549 12047 6607 12053
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 7377 12087 7435 12093
rect 7377 12053 7389 12087
rect 7423 12084 7435 12087
rect 8202 12084 8208 12096
rect 7423 12056 8208 12084
rect 7423 12053 7435 12056
rect 7377 12047 7435 12053
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 8294 12044 8300 12096
rect 8352 12084 8358 12096
rect 10781 12087 10839 12093
rect 10781 12084 10793 12087
rect 8352 12056 10793 12084
rect 8352 12044 8358 12056
rect 10781 12053 10793 12056
rect 10827 12053 10839 12087
rect 10781 12047 10839 12053
rect 10870 12044 10876 12096
rect 10928 12044 10934 12096
rect 10965 12087 11023 12093
rect 10965 12053 10977 12087
rect 11011 12084 11023 12087
rect 11146 12084 11152 12096
rect 11011 12056 11152 12084
rect 11011 12053 11023 12056
rect 10965 12047 11023 12053
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 11977 12087 12035 12093
rect 11977 12053 11989 12087
rect 12023 12084 12035 12087
rect 14182 12084 14188 12096
rect 12023 12056 14188 12084
rect 12023 12053 12035 12056
rect 11977 12047 12035 12053
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 16408 12084 16436 12192
rect 16482 12180 16488 12192
rect 16540 12180 16546 12232
rect 18049 12087 18107 12093
rect 18049 12084 18061 12087
rect 16408 12056 18061 12084
rect 18049 12053 18061 12056
rect 18095 12053 18107 12087
rect 18049 12047 18107 12053
rect 1104 11994 18860 12016
rect 1104 11942 3947 11994
rect 3999 11942 4011 11994
rect 4063 11942 4075 11994
rect 4127 11942 4139 11994
rect 4191 11942 9878 11994
rect 9930 11942 9942 11994
rect 9994 11942 10006 11994
rect 10058 11942 10070 11994
rect 10122 11942 15808 11994
rect 15860 11942 15872 11994
rect 15924 11942 15936 11994
rect 15988 11942 16000 11994
rect 16052 11942 18860 11994
rect 1104 11920 18860 11942
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 2593 11883 2651 11889
rect 2593 11880 2605 11883
rect 2464 11852 2605 11880
rect 2464 11840 2470 11852
rect 2593 11849 2605 11852
rect 2639 11849 2651 11883
rect 2593 11843 2651 11849
rect 3786 11840 3792 11892
rect 3844 11880 3850 11892
rect 5721 11883 5779 11889
rect 3844 11852 4568 11880
rect 3844 11840 3850 11852
rect 1581 11815 1639 11821
rect 1581 11781 1593 11815
rect 1627 11812 1639 11815
rect 2774 11812 2780 11824
rect 1627 11784 2780 11812
rect 1627 11781 1639 11784
rect 1581 11775 1639 11781
rect 2774 11772 2780 11784
rect 2832 11772 2838 11824
rect 4540 11812 4568 11852
rect 5721 11849 5733 11883
rect 5767 11880 5779 11883
rect 6270 11880 6276 11892
rect 5767 11852 6276 11880
rect 5767 11849 5779 11852
rect 5721 11843 5779 11849
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 8938 11880 8944 11892
rect 8899 11852 8944 11880
rect 8938 11840 8944 11852
rect 8996 11840 9002 11892
rect 9030 11840 9036 11892
rect 9088 11880 9094 11892
rect 11790 11880 11796 11892
rect 9088 11852 11796 11880
rect 9088 11840 9094 11852
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 12342 11840 12348 11892
rect 12400 11880 12406 11892
rect 12529 11883 12587 11889
rect 12529 11880 12541 11883
rect 12400 11852 12541 11880
rect 12400 11840 12406 11852
rect 12529 11849 12541 11852
rect 12575 11849 12587 11883
rect 12529 11843 12587 11849
rect 13817 11883 13875 11889
rect 13817 11849 13829 11883
rect 13863 11880 13875 11883
rect 13906 11880 13912 11892
rect 13863 11852 13912 11880
rect 13863 11849 13875 11852
rect 13817 11843 13875 11849
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 13998 11840 14004 11892
rect 14056 11880 14062 11892
rect 14918 11880 14924 11892
rect 14056 11852 14924 11880
rect 14056 11840 14062 11852
rect 14918 11840 14924 11852
rect 14976 11840 14982 11892
rect 16390 11840 16396 11892
rect 16448 11880 16454 11892
rect 16945 11883 17003 11889
rect 16945 11880 16957 11883
rect 16448 11852 16957 11880
rect 16448 11840 16454 11852
rect 16945 11849 16957 11852
rect 16991 11849 17003 11883
rect 16945 11843 17003 11849
rect 7466 11812 7472 11824
rect 4540 11784 7472 11812
rect 7466 11772 7472 11784
rect 7524 11772 7530 11824
rect 8570 11772 8576 11824
rect 8628 11812 8634 11824
rect 10686 11812 10692 11824
rect 8628 11784 10548 11812
rect 10647 11784 10692 11812
rect 8628 11772 8634 11784
rect 2038 11704 2044 11756
rect 2096 11744 2102 11756
rect 2225 11747 2283 11753
rect 2225 11744 2237 11747
rect 2096 11716 2237 11744
rect 2096 11704 2102 11716
rect 2225 11713 2237 11716
rect 2271 11744 2283 11747
rect 2590 11744 2596 11756
rect 2271 11716 2596 11744
rect 2271 11713 2283 11716
rect 2225 11707 2283 11713
rect 2590 11704 2596 11716
rect 2648 11704 2654 11756
rect 3237 11747 3295 11753
rect 3237 11713 3249 11747
rect 3283 11744 3295 11747
rect 5258 11744 5264 11756
rect 3283 11716 3740 11744
rect 5219 11716 5264 11744
rect 3283 11713 3295 11716
rect 3237 11707 3295 11713
rect 3605 11679 3663 11685
rect 3605 11645 3617 11679
rect 3651 11645 3663 11679
rect 3605 11639 3663 11645
rect 1949 11611 2007 11617
rect 1949 11577 1961 11611
rect 1995 11608 2007 11611
rect 2866 11608 2872 11620
rect 1995 11580 2872 11608
rect 1995 11577 2007 11580
rect 1949 11571 2007 11577
rect 2866 11568 2872 11580
rect 2924 11568 2930 11620
rect 2961 11611 3019 11617
rect 2961 11577 2973 11611
rect 3007 11608 3019 11611
rect 3510 11608 3516 11620
rect 3007 11580 3516 11608
rect 3007 11577 3019 11580
rect 2961 11571 3019 11577
rect 3510 11568 3516 11580
rect 3568 11568 3574 11620
rect 2041 11543 2099 11549
rect 2041 11509 2053 11543
rect 2087 11540 2099 11543
rect 2774 11540 2780 11552
rect 2087 11512 2780 11540
rect 2087 11509 2099 11512
rect 2041 11503 2099 11509
rect 2774 11500 2780 11512
rect 2832 11500 2838 11552
rect 3053 11543 3111 11549
rect 3053 11509 3065 11543
rect 3099 11540 3111 11543
rect 3418 11540 3424 11552
rect 3099 11512 3424 11540
rect 3099 11509 3111 11512
rect 3053 11503 3111 11509
rect 3418 11500 3424 11512
rect 3476 11500 3482 11552
rect 3620 11540 3648 11639
rect 3712 11608 3740 11716
rect 5258 11704 5264 11716
rect 5316 11704 5322 11756
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11744 6423 11747
rect 6914 11744 6920 11756
rect 6411 11716 6920 11744
rect 6411 11713 6423 11716
rect 6365 11707 6423 11713
rect 6914 11704 6920 11716
rect 6972 11704 6978 11756
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 9217 11747 9275 11753
rect 9217 11744 9229 11747
rect 8904 11716 9229 11744
rect 8904 11704 8910 11716
rect 9217 11713 9229 11716
rect 9263 11713 9275 11747
rect 10318 11744 10324 11756
rect 10279 11716 10324 11744
rect 9217 11707 9275 11713
rect 10318 11704 10324 11716
rect 10376 11704 10382 11756
rect 10520 11744 10548 11784
rect 10686 11772 10692 11784
rect 10744 11772 10750 11824
rect 15010 11812 15016 11824
rect 10796 11784 15016 11812
rect 10796 11744 10824 11784
rect 15010 11772 15016 11784
rect 15068 11772 15074 11824
rect 16669 11815 16727 11821
rect 16669 11781 16681 11815
rect 16715 11812 16727 11815
rect 17126 11812 17132 11824
rect 16715 11784 17132 11812
rect 16715 11781 16727 11784
rect 16669 11775 16727 11781
rect 17126 11772 17132 11784
rect 17184 11812 17190 11824
rect 17184 11784 17540 11812
rect 17184 11772 17190 11784
rect 11146 11744 11152 11756
rect 10520 11716 10824 11744
rect 11107 11716 11152 11744
rect 11146 11704 11152 11716
rect 11204 11704 11210 11756
rect 11330 11744 11336 11756
rect 11291 11716 11336 11744
rect 11330 11704 11336 11716
rect 11388 11704 11394 11756
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 13081 11747 13139 11753
rect 13081 11744 13093 11747
rect 12124 11716 13093 11744
rect 12124 11704 12130 11716
rect 13081 11713 13093 11716
rect 13127 11713 13139 11747
rect 14458 11744 14464 11756
rect 13081 11707 13139 11713
rect 13648 11716 14320 11744
rect 14419 11716 14464 11744
rect 3872 11679 3930 11685
rect 3872 11645 3884 11679
rect 3918 11676 3930 11679
rect 4246 11676 4252 11688
rect 3918 11648 4252 11676
rect 3918 11645 3930 11648
rect 3872 11639 3930 11645
rect 4246 11636 4252 11648
rect 4304 11636 4310 11688
rect 4706 11636 4712 11688
rect 4764 11676 4770 11688
rect 7006 11676 7012 11688
rect 4764 11648 7012 11676
rect 4764 11636 4770 11648
rect 7006 11636 7012 11648
rect 7064 11636 7070 11688
rect 7561 11679 7619 11685
rect 7561 11645 7573 11679
rect 7607 11676 7619 11679
rect 7650 11676 7656 11688
rect 7607 11648 7656 11676
rect 7607 11645 7619 11648
rect 7561 11639 7619 11645
rect 7650 11636 7656 11648
rect 7708 11636 7714 11688
rect 7828 11679 7886 11685
rect 7828 11645 7840 11679
rect 7874 11676 7886 11679
rect 9122 11676 9128 11688
rect 7874 11648 9128 11676
rect 7874 11645 7886 11648
rect 7828 11639 7886 11645
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 10505 11679 10563 11685
rect 10505 11676 10517 11679
rect 9232 11648 10517 11676
rect 3786 11608 3792 11620
rect 3712 11580 3792 11608
rect 3786 11568 3792 11580
rect 3844 11568 3850 11620
rect 3970 11568 3976 11620
rect 4028 11608 4034 11620
rect 6181 11611 6239 11617
rect 6181 11608 6193 11611
rect 4028 11580 6193 11608
rect 4028 11568 4034 11580
rect 6181 11577 6193 11580
rect 6227 11608 6239 11611
rect 9232 11608 9260 11648
rect 10505 11645 10517 11648
rect 10551 11645 10563 11679
rect 10505 11639 10563 11645
rect 10686 11636 10692 11688
rect 10744 11676 10750 11688
rect 13648 11676 13676 11716
rect 10744 11648 13676 11676
rect 10744 11636 10750 11648
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 14185 11679 14243 11685
rect 14185 11676 14197 11679
rect 13780 11648 14197 11676
rect 13780 11636 13786 11648
rect 14185 11645 14197 11648
rect 14231 11645 14243 11679
rect 14185 11639 14243 11645
rect 11057 11611 11115 11617
rect 11057 11608 11069 11611
rect 6227 11580 9260 11608
rect 9692 11580 11069 11608
rect 6227 11577 6239 11580
rect 6181 11571 6239 11577
rect 4430 11540 4436 11552
rect 3620 11512 4436 11540
rect 4430 11500 4436 11512
rect 4488 11500 4494 11552
rect 4982 11540 4988 11552
rect 4943 11512 4988 11540
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 6086 11540 6092 11552
rect 6047 11512 6092 11540
rect 6086 11500 6092 11512
rect 6144 11500 6150 11552
rect 6362 11500 6368 11552
rect 6420 11540 6426 11552
rect 9582 11540 9588 11552
rect 6420 11512 9588 11540
rect 6420 11500 6426 11512
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 9692 11549 9720 11580
rect 11057 11577 11069 11580
rect 11103 11577 11115 11611
rect 11057 11571 11115 11577
rect 12897 11611 12955 11617
rect 12897 11577 12909 11611
rect 12943 11608 12955 11611
rect 13906 11608 13912 11620
rect 12943 11580 13912 11608
rect 12943 11577 12955 11580
rect 12897 11571 12955 11577
rect 13906 11568 13912 11580
rect 13964 11568 13970 11620
rect 14292 11608 14320 11716
rect 14458 11704 14464 11716
rect 14516 11704 14522 11756
rect 15286 11744 15292 11756
rect 15247 11716 15292 11744
rect 15286 11704 15292 11716
rect 15344 11704 15350 11756
rect 16482 11704 16488 11756
rect 16540 11744 16546 11756
rect 17402 11744 17408 11756
rect 16540 11716 17408 11744
rect 16540 11704 16546 11716
rect 17402 11704 17408 11716
rect 17460 11704 17466 11756
rect 17512 11753 17540 11784
rect 17497 11747 17555 11753
rect 17497 11713 17509 11747
rect 17543 11713 17555 11747
rect 17497 11707 17555 11713
rect 15556 11679 15614 11685
rect 15556 11645 15568 11679
rect 15602 11676 15614 11679
rect 16850 11676 16856 11688
rect 15602 11648 16856 11676
rect 15602 11645 15614 11648
rect 15556 11639 15614 11645
rect 16850 11636 16856 11648
rect 16908 11636 16914 11688
rect 17313 11611 17371 11617
rect 17313 11608 17325 11611
rect 14292 11580 17325 11608
rect 17313 11577 17325 11580
rect 17359 11608 17371 11611
rect 18138 11608 18144 11620
rect 17359 11580 18144 11608
rect 17359 11577 17371 11580
rect 17313 11571 17371 11577
rect 18138 11568 18144 11580
rect 18196 11568 18202 11620
rect 9677 11543 9735 11549
rect 9677 11509 9689 11543
rect 9723 11509 9735 11543
rect 10042 11540 10048 11552
rect 10003 11512 10048 11540
rect 9677 11503 9735 11509
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 10137 11543 10195 11549
rect 10137 11509 10149 11543
rect 10183 11540 10195 11543
rect 10505 11543 10563 11549
rect 10505 11540 10517 11543
rect 10183 11512 10517 11540
rect 10183 11509 10195 11512
rect 10137 11503 10195 11509
rect 10505 11509 10517 11512
rect 10551 11540 10563 11543
rect 11698 11540 11704 11552
rect 10551 11512 11704 11540
rect 10551 11509 10563 11512
rect 10505 11503 10563 11509
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 12989 11543 13047 11549
rect 12989 11509 13001 11543
rect 13035 11540 13047 11543
rect 13262 11540 13268 11552
rect 13035 11512 13268 11540
rect 13035 11509 13047 11512
rect 12989 11503 13047 11509
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 13630 11500 13636 11552
rect 13688 11540 13694 11552
rect 14274 11540 14280 11552
rect 13688 11512 14280 11540
rect 13688 11500 13694 11512
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 17402 11500 17408 11552
rect 17460 11540 17466 11552
rect 17460 11512 17505 11540
rect 17460 11500 17466 11512
rect 1104 11450 18860 11472
rect 1104 11398 6912 11450
rect 6964 11398 6976 11450
rect 7028 11398 7040 11450
rect 7092 11398 7104 11450
rect 7156 11398 12843 11450
rect 12895 11398 12907 11450
rect 12959 11398 12971 11450
rect 13023 11398 13035 11450
rect 13087 11398 18860 11450
rect 1104 11376 18860 11398
rect 2406 11296 2412 11348
rect 2464 11336 2470 11348
rect 2682 11336 2688 11348
rect 2464 11308 2688 11336
rect 2464 11296 2470 11308
rect 2682 11296 2688 11308
rect 2740 11336 2746 11348
rect 3697 11339 3755 11345
rect 3697 11336 3709 11339
rect 2740 11308 3709 11336
rect 2740 11296 2746 11308
rect 3697 11305 3709 11308
rect 3743 11305 3755 11339
rect 3697 11299 3755 11305
rect 4065 11339 4123 11345
rect 4065 11305 4077 11339
rect 4111 11336 4123 11339
rect 6825 11339 6883 11345
rect 4111 11308 6776 11336
rect 4111 11305 4123 11308
rect 4065 11299 4123 11305
rect 2314 11228 2320 11280
rect 2372 11228 2378 11280
rect 2590 11277 2596 11280
rect 2584 11268 2596 11277
rect 2551 11240 2596 11268
rect 2584 11231 2596 11240
rect 2590 11228 2596 11231
rect 2648 11228 2654 11280
rect 6748 11268 6776 11308
rect 6825 11305 6837 11339
rect 6871 11336 6883 11339
rect 9306 11336 9312 11348
rect 6871 11308 9312 11336
rect 6871 11305 6883 11308
rect 6825 11299 6883 11305
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 9582 11296 9588 11348
rect 9640 11336 9646 11348
rect 9640 11308 10272 11336
rect 9640 11296 9646 11308
rect 7006 11268 7012 11280
rect 6748 11240 7012 11268
rect 7006 11228 7012 11240
rect 7064 11228 7070 11280
rect 9122 11268 9128 11280
rect 7116 11240 9128 11268
rect 1673 11203 1731 11209
rect 1673 11169 1685 11203
rect 1719 11200 1731 11203
rect 2332 11200 2360 11228
rect 1719 11172 2360 11200
rect 1719 11169 1731 11172
rect 1673 11163 1731 11169
rect 3786 11160 3792 11212
rect 3844 11200 3850 11212
rect 4516 11203 4574 11209
rect 4516 11200 4528 11203
rect 3844 11172 4528 11200
rect 3844 11160 3850 11172
rect 4516 11169 4528 11172
rect 4562 11200 4574 11203
rect 4982 11200 4988 11212
rect 4562 11172 4988 11200
rect 4562 11169 4574 11172
rect 4516 11163 4574 11169
rect 4982 11160 4988 11172
rect 5040 11160 5046 11212
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11200 6147 11203
rect 6638 11200 6644 11212
rect 6135 11172 6644 11200
rect 6135 11169 6147 11172
rect 6089 11163 6147 11169
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 2038 11092 2044 11144
rect 2096 11132 2102 11144
rect 2317 11135 2375 11141
rect 2317 11132 2329 11135
rect 2096 11104 2329 11132
rect 2096 11092 2102 11104
rect 2317 11101 2329 11104
rect 2363 11101 2375 11135
rect 2317 11095 2375 11101
rect 3510 11092 3516 11144
rect 3568 11132 3574 11144
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 3568 11104 4077 11132
rect 3568 11092 3574 11104
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 4246 11132 4252 11144
rect 4207 11104 4252 11132
rect 4065 11095 4123 11101
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 5718 11092 5724 11144
rect 5776 11132 5782 11144
rect 7116 11141 7144 11240
rect 9122 11228 9128 11240
rect 9180 11268 9186 11280
rect 9922 11271 9980 11277
rect 9922 11268 9934 11271
rect 9180 11240 9934 11268
rect 9180 11228 9186 11240
rect 9922 11237 9934 11240
rect 9968 11237 9980 11271
rect 10244 11268 10272 11308
rect 10318 11296 10324 11348
rect 10376 11336 10382 11348
rect 11057 11339 11115 11345
rect 11057 11336 11069 11339
rect 10376 11308 11069 11336
rect 10376 11296 10382 11308
rect 11057 11305 11069 11308
rect 11103 11336 11115 11339
rect 11238 11336 11244 11348
rect 11103 11308 11244 11336
rect 11103 11305 11115 11308
rect 11057 11299 11115 11305
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 12066 11296 12072 11348
rect 12124 11336 12130 11348
rect 12124 11308 12563 11336
rect 12124 11296 12130 11308
rect 10686 11268 10692 11280
rect 10244 11240 10692 11268
rect 9922 11231 9980 11237
rect 10686 11228 10692 11240
rect 10744 11228 10750 11280
rect 11974 11268 11980 11280
rect 11624 11240 11980 11268
rect 7377 11203 7435 11209
rect 7377 11169 7389 11203
rect 7423 11200 7435 11203
rect 7653 11203 7711 11209
rect 7653 11200 7665 11203
rect 7423 11172 7665 11200
rect 7423 11169 7435 11172
rect 7377 11163 7435 11169
rect 7653 11169 7665 11172
rect 7699 11169 7711 11203
rect 7653 11163 7711 11169
rect 8196 11203 8254 11209
rect 8196 11169 8208 11203
rect 8242 11200 8254 11203
rect 8938 11200 8944 11212
rect 8242 11172 8944 11200
rect 8242 11169 8254 11172
rect 8196 11163 8254 11169
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 9582 11160 9588 11212
rect 9640 11200 9646 11212
rect 11624 11209 11652 11240
rect 11974 11228 11980 11240
rect 12032 11228 12038 11280
rect 12535 11277 12563 11308
rect 12618 11296 12624 11348
rect 12676 11336 12682 11348
rect 13633 11339 13691 11345
rect 13633 11336 13645 11339
rect 12676 11308 13645 11336
rect 12676 11296 12682 11308
rect 13633 11305 13645 11308
rect 13679 11336 13691 11339
rect 13722 11336 13728 11348
rect 13679 11308 13728 11336
rect 13679 11305 13691 11308
rect 13633 11299 13691 11305
rect 13722 11296 13728 11308
rect 13780 11296 13786 11348
rect 13906 11336 13912 11348
rect 13867 11308 13912 11336
rect 13906 11296 13912 11308
rect 13964 11296 13970 11348
rect 14369 11339 14427 11345
rect 14369 11305 14381 11339
rect 14415 11336 14427 11339
rect 15010 11336 15016 11348
rect 14415 11308 15016 11336
rect 14415 11305 14427 11308
rect 14369 11299 14427 11305
rect 15010 11296 15016 11308
rect 15068 11296 15074 11348
rect 16669 11339 16727 11345
rect 16669 11305 16681 11339
rect 16715 11336 16727 11339
rect 16850 11336 16856 11348
rect 16715 11308 16856 11336
rect 16715 11305 16727 11308
rect 16669 11299 16727 11305
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 12520 11271 12578 11277
rect 12520 11237 12532 11271
rect 12566 11237 12578 11271
rect 12520 11231 12578 11237
rect 13814 11228 13820 11280
rect 13872 11268 13878 11280
rect 15556 11271 15614 11277
rect 13872 11240 15332 11268
rect 13872 11228 13878 11240
rect 15304 11212 15332 11240
rect 15556 11237 15568 11271
rect 15602 11268 15614 11271
rect 17770 11268 17776 11280
rect 15602 11240 17776 11268
rect 15602 11237 15614 11240
rect 15556 11231 15614 11237
rect 17770 11228 17776 11240
rect 17828 11228 17834 11280
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 9640 11172 9689 11200
rect 9640 11160 9646 11172
rect 9677 11169 9689 11172
rect 9723 11200 9735 11203
rect 11609 11203 11667 11209
rect 9723 11172 10732 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 6917 11135 6975 11141
rect 6917 11132 6929 11135
rect 5776 11104 6929 11132
rect 5776 11092 5782 11104
rect 6917 11101 6929 11104
rect 6963 11101 6975 11135
rect 6917 11095 6975 11101
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11101 7159 11135
rect 7101 11095 7159 11101
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 1394 11024 1400 11076
rect 1452 11064 1458 11076
rect 1857 11067 1915 11073
rect 1857 11064 1869 11067
rect 1452 11036 1869 11064
rect 1452 11024 1458 11036
rect 1857 11033 1869 11036
rect 1903 11033 1915 11067
rect 1857 11027 1915 11033
rect 3326 11024 3332 11076
rect 3384 11064 3390 11076
rect 3970 11064 3976 11076
rect 3384 11036 3976 11064
rect 3384 11024 3390 11036
rect 3970 11024 3976 11036
rect 4028 11024 4034 11076
rect 5810 11024 5816 11076
rect 5868 11064 5874 11076
rect 5905 11067 5963 11073
rect 5905 11064 5917 11067
rect 5868 11036 5917 11064
rect 5868 11024 5874 11036
rect 5905 11033 5917 11036
rect 5951 11033 5963 11067
rect 6454 11064 6460 11076
rect 6415 11036 6460 11064
rect 5905 11027 5963 11033
rect 2590 10956 2596 11008
rect 2648 10996 2654 11008
rect 5629 10999 5687 11005
rect 5629 10996 5641 10999
rect 2648 10968 5641 10996
rect 2648 10956 2654 10968
rect 5629 10965 5641 10968
rect 5675 10965 5687 10999
rect 5920 10996 5948 11027
rect 6454 11024 6460 11036
rect 6512 11024 6518 11076
rect 7377 11067 7435 11073
rect 7377 11064 7389 11067
rect 6840 11036 7389 11064
rect 6840 10996 6868 11036
rect 7377 11033 7389 11036
rect 7423 11033 7435 11067
rect 7377 11027 7435 11033
rect 5920 10968 6868 10996
rect 7469 10999 7527 11005
rect 5629 10959 5687 10965
rect 7469 10965 7481 10999
rect 7515 10996 7527 10999
rect 7650 10996 7656 11008
rect 7515 10968 7656 10996
rect 7515 10965 7527 10968
rect 7469 10959 7527 10965
rect 7650 10956 7656 10968
rect 7708 10996 7714 11008
rect 7944 10996 7972 11095
rect 9309 11067 9367 11073
rect 9309 11033 9321 11067
rect 9355 11064 9367 11067
rect 9355 11036 9720 11064
rect 9355 11033 9367 11036
rect 9309 11027 9367 11033
rect 7708 10968 7972 10996
rect 9692 10996 9720 11036
rect 10704 11008 10732 11172
rect 11609 11169 11621 11203
rect 11655 11169 11667 11203
rect 11609 11163 11667 11169
rect 11698 11160 11704 11212
rect 11756 11200 11762 11212
rect 13998 11200 14004 11212
rect 11756 11172 14004 11200
rect 11756 11160 11762 11172
rect 13998 11160 14004 11172
rect 14056 11160 14062 11212
rect 14274 11200 14280 11212
rect 14235 11172 14280 11200
rect 14274 11160 14280 11172
rect 14332 11160 14338 11212
rect 14826 11160 14832 11212
rect 14884 11200 14890 11212
rect 15105 11203 15163 11209
rect 15105 11200 15117 11203
rect 14884 11172 15117 11200
rect 14884 11160 14890 11172
rect 15105 11169 15117 11172
rect 15151 11169 15163 11203
rect 15286 11200 15292 11212
rect 15247 11172 15292 11200
rect 15105 11163 15163 11169
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 16390 11160 16396 11212
rect 16448 11200 16454 11212
rect 16666 11200 16672 11212
rect 16448 11172 16672 11200
rect 16448 11160 16454 11172
rect 16666 11160 16672 11172
rect 16724 11160 16730 11212
rect 17126 11160 17132 11212
rect 17184 11200 17190 11212
rect 17313 11203 17371 11209
rect 17313 11200 17325 11203
rect 17184 11172 17325 11200
rect 17184 11160 17190 11172
rect 17313 11169 17325 11172
rect 17359 11169 17371 11203
rect 17313 11163 17371 11169
rect 12250 11132 12256 11144
rect 12211 11104 12256 11132
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 13906 11092 13912 11144
rect 13964 11132 13970 11144
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 13964 11104 14473 11132
rect 13964 11092 13970 11104
rect 14461 11101 14473 11104
rect 14507 11101 14519 11135
rect 15194 11132 15200 11144
rect 14461 11095 14519 11101
rect 14660 11104 15200 11132
rect 10318 10996 10324 11008
rect 9692 10968 10324 10996
rect 7708 10956 7714 10968
rect 10318 10956 10324 10968
rect 10376 10956 10382 11008
rect 10686 10956 10692 11008
rect 10744 10996 10750 11008
rect 11422 10996 11428 11008
rect 10744 10968 11428 10996
rect 10744 10956 10750 10968
rect 11422 10956 11428 10968
rect 11480 10996 11486 11008
rect 12268 10996 12296 11092
rect 13354 11024 13360 11076
rect 13412 11064 13418 11076
rect 14660 11064 14688 11104
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 13412 11036 14688 11064
rect 14921 11067 14979 11073
rect 13412 11024 13418 11036
rect 14921 11033 14933 11067
rect 14967 11064 14979 11067
rect 15304 11064 15332 11160
rect 17405 11135 17463 11141
rect 17405 11101 17417 11135
rect 17451 11101 17463 11135
rect 17405 11095 17463 11101
rect 17589 11135 17647 11141
rect 17589 11101 17601 11135
rect 17635 11132 17647 11135
rect 17678 11132 17684 11144
rect 17635 11104 17684 11132
rect 17635 11101 17647 11104
rect 17589 11095 17647 11101
rect 16942 11064 16948 11076
rect 14967 11036 15332 11064
rect 16903 11036 16948 11064
rect 14967 11033 14979 11036
rect 14921 11027 14979 11033
rect 16942 11024 16948 11036
rect 17000 11024 17006 11076
rect 17310 11024 17316 11076
rect 17368 11064 17374 11076
rect 17420 11064 17448 11095
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 17368 11036 17448 11064
rect 17368 11024 17374 11036
rect 11480 10968 12296 10996
rect 11480 10956 11486 10968
rect 13170 10956 13176 11008
rect 13228 10996 13234 11008
rect 17034 10996 17040 11008
rect 13228 10968 17040 10996
rect 13228 10956 13234 10968
rect 17034 10956 17040 10968
rect 17092 10956 17098 11008
rect 1104 10906 18860 10928
rect 1104 10854 3947 10906
rect 3999 10854 4011 10906
rect 4063 10854 4075 10906
rect 4127 10854 4139 10906
rect 4191 10854 9878 10906
rect 9930 10854 9942 10906
rect 9994 10854 10006 10906
rect 10058 10854 10070 10906
rect 10122 10854 15808 10906
rect 15860 10854 15872 10906
rect 15924 10854 15936 10906
rect 15988 10854 16000 10906
rect 16052 10854 18860 10906
rect 1104 10832 18860 10854
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 3697 10795 3755 10801
rect 3697 10792 3709 10795
rect 2832 10764 3709 10792
rect 2832 10752 2838 10764
rect 3697 10761 3709 10764
rect 3743 10761 3755 10795
rect 5166 10792 5172 10804
rect 3697 10755 3755 10761
rect 4172 10764 5172 10792
rect 4172 10736 4200 10764
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 8018 10792 8024 10804
rect 7064 10764 8024 10792
rect 7064 10752 7070 10764
rect 8018 10752 8024 10764
rect 8076 10792 8082 10804
rect 9122 10792 9128 10804
rect 8076 10764 8892 10792
rect 9083 10764 9128 10792
rect 8076 10752 8082 10764
rect 4154 10684 4160 10736
rect 4212 10684 4218 10736
rect 4709 10727 4767 10733
rect 4709 10693 4721 10727
rect 4755 10724 4767 10727
rect 5994 10724 6000 10736
rect 4755 10696 6000 10724
rect 4755 10693 4767 10696
rect 4709 10687 4767 10693
rect 5994 10684 6000 10696
rect 6052 10684 6058 10736
rect 3510 10616 3516 10668
rect 3568 10656 3574 10668
rect 3786 10656 3792 10668
rect 3568 10628 3792 10656
rect 3568 10616 3574 10628
rect 3786 10616 3792 10628
rect 3844 10656 3850 10668
rect 4249 10659 4307 10665
rect 4249 10656 4261 10659
rect 3844 10628 4261 10656
rect 3844 10616 3850 10628
rect 4249 10625 4261 10628
rect 4295 10625 4307 10659
rect 4249 10619 4307 10625
rect 5353 10659 5411 10665
rect 5353 10625 5365 10659
rect 5399 10656 5411 10659
rect 5902 10656 5908 10668
rect 5399 10628 5908 10656
rect 5399 10625 5411 10628
rect 5353 10619 5411 10625
rect 5902 10616 5908 10628
rect 5960 10616 5966 10668
rect 6270 10656 6276 10668
rect 6231 10628 6276 10656
rect 6270 10616 6276 10628
rect 6328 10616 6334 10668
rect 7650 10616 7656 10668
rect 7708 10656 7714 10668
rect 7745 10659 7803 10665
rect 7745 10656 7757 10659
rect 7708 10628 7757 10656
rect 7708 10616 7714 10628
rect 7745 10625 7757 10628
rect 7791 10625 7803 10659
rect 8864 10656 8892 10764
rect 9122 10752 9128 10764
rect 9180 10752 9186 10804
rect 9490 10752 9496 10804
rect 9548 10792 9554 10804
rect 12161 10795 12219 10801
rect 9548 10764 11744 10792
rect 9548 10752 9554 10764
rect 8938 10684 8944 10736
rect 8996 10724 9002 10736
rect 8996 10696 9996 10724
rect 8996 10684 9002 10696
rect 8864 10628 9628 10656
rect 7745 10619 7803 10625
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10557 1455 10591
rect 1397 10551 1455 10557
rect 1664 10591 1722 10597
rect 1664 10557 1676 10591
rect 1710 10588 1722 10591
rect 2406 10588 2412 10600
rect 1710 10560 2412 10588
rect 1710 10557 1722 10560
rect 1664 10551 1722 10557
rect 1412 10520 1440 10551
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 3053 10591 3111 10597
rect 3053 10557 3065 10591
rect 3099 10588 3111 10591
rect 6181 10591 6239 10597
rect 6181 10588 6193 10591
rect 3099 10560 6193 10588
rect 3099 10557 3111 10560
rect 3053 10551 3111 10557
rect 6181 10557 6193 10560
rect 6227 10588 6239 10591
rect 7558 10588 7564 10600
rect 6227 10560 7564 10588
rect 6227 10557 6239 10560
rect 6181 10551 6239 10557
rect 7558 10548 7564 10560
rect 7616 10548 7622 10600
rect 7834 10548 7840 10600
rect 7892 10588 7898 10600
rect 7892 10560 9444 10588
rect 7892 10548 7898 10560
rect 2038 10520 2044 10532
rect 1412 10492 2044 10520
rect 2038 10480 2044 10492
rect 2096 10480 2102 10532
rect 3418 10480 3424 10532
rect 3476 10520 3482 10532
rect 8018 10529 8024 10532
rect 6089 10523 6147 10529
rect 3476 10492 5856 10520
rect 3476 10480 3482 10492
rect 2498 10412 2504 10464
rect 2556 10452 2562 10464
rect 2777 10455 2835 10461
rect 2777 10452 2789 10455
rect 2556 10424 2789 10452
rect 2556 10412 2562 10424
rect 2777 10421 2789 10424
rect 2823 10421 2835 10455
rect 3234 10452 3240 10464
rect 3195 10424 3240 10452
rect 2777 10415 2835 10421
rect 3234 10412 3240 10424
rect 3292 10412 3298 10464
rect 4062 10452 4068 10464
rect 4023 10424 4068 10452
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 4157 10455 4215 10461
rect 4157 10421 4169 10455
rect 4203 10452 4215 10455
rect 4706 10452 4712 10464
rect 4203 10424 4712 10452
rect 4203 10421 4215 10424
rect 4157 10415 4215 10421
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 5074 10452 5080 10464
rect 5035 10424 5080 10452
rect 5074 10412 5080 10424
rect 5132 10412 5138 10464
rect 5166 10412 5172 10464
rect 5224 10452 5230 10464
rect 5224 10424 5269 10452
rect 5224 10412 5230 10424
rect 5442 10412 5448 10464
rect 5500 10452 5506 10464
rect 5721 10455 5779 10461
rect 5721 10452 5733 10455
rect 5500 10424 5733 10452
rect 5500 10412 5506 10424
rect 5721 10421 5733 10424
rect 5767 10421 5779 10455
rect 5828 10452 5856 10492
rect 6089 10489 6101 10523
rect 6135 10520 6147 10523
rect 8012 10520 8024 10529
rect 6135 10492 7880 10520
rect 7979 10492 8024 10520
rect 6135 10489 6147 10492
rect 6089 10483 6147 10489
rect 6730 10452 6736 10464
rect 5828 10424 6736 10452
rect 5721 10415 5779 10421
rect 6730 10412 6736 10424
rect 6788 10412 6794 10464
rect 7852 10452 7880 10492
rect 8012 10483 8024 10492
rect 8018 10480 8024 10483
rect 8076 10480 8082 10532
rect 8570 10452 8576 10464
rect 7852 10424 8576 10452
rect 8570 10412 8576 10424
rect 8628 10412 8634 10464
rect 9416 10461 9444 10560
rect 9401 10455 9459 10461
rect 9401 10421 9413 10455
rect 9447 10421 9459 10455
rect 9600 10452 9628 10628
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 9968 10665 9996 10696
rect 9861 10659 9919 10665
rect 9861 10656 9873 10659
rect 9732 10628 9873 10656
rect 9732 10616 9738 10628
rect 9861 10625 9873 10628
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10625 10011 10659
rect 10686 10656 10692 10668
rect 10647 10628 10692 10656
rect 9953 10619 10011 10625
rect 10686 10616 10692 10628
rect 10744 10616 10750 10668
rect 9766 10588 9772 10600
rect 9727 10560 9772 10588
rect 9766 10548 9772 10560
rect 9824 10548 9830 10600
rect 11716 10588 11744 10764
rect 12161 10761 12173 10795
rect 12207 10792 12219 10795
rect 16206 10792 16212 10804
rect 12207 10764 16212 10792
rect 12207 10761 12219 10764
rect 12161 10755 12219 10761
rect 16206 10752 16212 10764
rect 16264 10752 16270 10804
rect 16574 10792 16580 10804
rect 16316 10764 16580 10792
rect 12066 10724 12072 10736
rect 12027 10696 12072 10724
rect 12066 10684 12072 10696
rect 12124 10684 12130 10736
rect 15289 10727 15347 10733
rect 15289 10693 15301 10727
rect 15335 10724 15347 10727
rect 16316 10724 16344 10764
rect 16574 10752 16580 10764
rect 16632 10752 16638 10804
rect 16666 10752 16672 10804
rect 16724 10792 16730 10804
rect 17494 10792 17500 10804
rect 16724 10764 17500 10792
rect 16724 10752 16730 10764
rect 17494 10752 17500 10764
rect 17552 10752 17558 10804
rect 15335 10696 16344 10724
rect 15335 10693 15347 10696
rect 15289 10687 15347 10693
rect 13078 10656 13084 10668
rect 13039 10628 13084 10656
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 14458 10616 14464 10668
rect 14516 10656 14522 10668
rect 14642 10656 14648 10668
rect 14516 10628 14648 10656
rect 14516 10616 14522 10628
rect 14642 10616 14648 10628
rect 14700 10616 14706 10668
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10656 15991 10659
rect 15979 10628 16436 10656
rect 15979 10625 15991 10628
rect 15933 10619 15991 10625
rect 13722 10597 13728 10600
rect 13357 10591 13415 10597
rect 13357 10588 13369 10591
rect 11716 10560 13369 10588
rect 13357 10557 13369 10560
rect 13403 10557 13415 10591
rect 13357 10551 13415 10557
rect 13449 10591 13507 10597
rect 13449 10557 13461 10591
rect 13495 10557 13507 10591
rect 13449 10551 13507 10557
rect 13716 10551 13728 10597
rect 13780 10588 13786 10600
rect 13780 10560 13816 10588
rect 10956 10523 11014 10529
rect 10956 10489 10968 10523
rect 11002 10520 11014 10523
rect 11698 10520 11704 10532
rect 11002 10492 11704 10520
rect 11002 10489 11014 10492
rect 10956 10483 11014 10489
rect 11698 10480 11704 10492
rect 11756 10480 11762 10532
rect 12250 10480 12256 10532
rect 12308 10520 12314 10532
rect 12897 10523 12955 10529
rect 12897 10520 12909 10523
rect 12308 10492 12909 10520
rect 12308 10480 12314 10492
rect 12897 10489 12909 10492
rect 12943 10489 12955 10523
rect 13464 10520 13492 10551
rect 13722 10548 13728 10551
rect 13780 10548 13786 10560
rect 14918 10548 14924 10600
rect 14976 10588 14982 10600
rect 15749 10591 15807 10597
rect 15749 10588 15761 10591
rect 14976 10560 15761 10588
rect 14976 10548 14982 10560
rect 15749 10557 15761 10560
rect 15795 10588 15807 10591
rect 16114 10588 16120 10600
rect 15795 10560 16120 10588
rect 15795 10557 15807 10560
rect 15749 10551 15807 10557
rect 16114 10548 16120 10560
rect 16172 10548 16178 10600
rect 16298 10588 16304 10600
rect 16259 10560 16304 10588
rect 16298 10548 16304 10560
rect 16356 10548 16362 10600
rect 16408 10588 16436 10628
rect 17862 10616 17868 10668
rect 17920 10656 17926 10668
rect 18049 10659 18107 10665
rect 18049 10656 18061 10659
rect 17920 10628 18061 10656
rect 17920 10616 17926 10628
rect 18049 10625 18061 10628
rect 18095 10625 18107 10659
rect 18049 10619 18107 10625
rect 16568 10591 16626 10597
rect 16568 10588 16580 10591
rect 16408 10560 16580 10588
rect 16568 10557 16580 10560
rect 16614 10588 16626 10591
rect 17678 10588 17684 10600
rect 16614 10560 17684 10588
rect 16614 10557 16626 10560
rect 16568 10551 16626 10557
rect 17678 10548 17684 10560
rect 17736 10548 17742 10600
rect 13814 10520 13820 10532
rect 13464 10492 13820 10520
rect 12897 10483 12955 10489
rect 13814 10480 13820 10492
rect 13872 10480 13878 10532
rect 15657 10523 15715 10529
rect 15657 10520 15669 10523
rect 13924 10492 15669 10520
rect 12161 10455 12219 10461
rect 12161 10452 12173 10455
rect 9600 10424 12173 10452
rect 9401 10415 9459 10421
rect 12161 10421 12173 10424
rect 12207 10421 12219 10455
rect 12161 10415 12219 10421
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12526 10452 12532 10464
rect 12483 10424 12532 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 12805 10455 12863 10461
rect 12805 10452 12817 10455
rect 12768 10424 12817 10452
rect 12768 10412 12774 10424
rect 12805 10421 12817 10424
rect 12851 10452 12863 10455
rect 13170 10452 13176 10464
rect 12851 10424 13176 10452
rect 12851 10421 12863 10424
rect 12805 10415 12863 10421
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 13357 10455 13415 10461
rect 13357 10421 13369 10455
rect 13403 10452 13415 10455
rect 13924 10452 13952 10492
rect 15657 10489 15669 10492
rect 15703 10520 15715 10523
rect 18046 10520 18052 10532
rect 15703 10492 18052 10520
rect 15703 10489 15715 10492
rect 15657 10483 15715 10489
rect 18046 10480 18052 10492
rect 18104 10480 18110 10532
rect 14826 10452 14832 10464
rect 13403 10424 13952 10452
rect 14787 10424 14832 10452
rect 13403 10421 13415 10424
rect 13357 10415 13415 10421
rect 14826 10412 14832 10424
rect 14884 10412 14890 10464
rect 17586 10412 17592 10464
rect 17644 10452 17650 10464
rect 17681 10455 17739 10461
rect 17681 10452 17693 10455
rect 17644 10424 17693 10452
rect 17644 10412 17650 10424
rect 17681 10421 17693 10424
rect 17727 10452 17739 10455
rect 17770 10452 17776 10464
rect 17727 10424 17776 10452
rect 17727 10421 17739 10424
rect 17681 10415 17739 10421
rect 17770 10412 17776 10424
rect 17828 10412 17834 10464
rect 1104 10362 18860 10384
rect 1104 10310 6912 10362
rect 6964 10310 6976 10362
rect 7028 10310 7040 10362
rect 7092 10310 7104 10362
rect 7156 10310 12843 10362
rect 12895 10310 12907 10362
rect 12959 10310 12971 10362
rect 13023 10310 13035 10362
rect 13087 10310 18860 10362
rect 1104 10288 18860 10310
rect 2222 10248 2228 10260
rect 2183 10220 2228 10248
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 2866 10208 2872 10260
rect 2924 10248 2930 10260
rect 2961 10251 3019 10257
rect 2961 10248 2973 10251
rect 2924 10220 2973 10248
rect 2924 10208 2930 10220
rect 2961 10217 2973 10220
rect 3007 10217 3019 10251
rect 2961 10211 3019 10217
rect 4430 10208 4436 10260
rect 4488 10248 4494 10260
rect 4617 10251 4675 10257
rect 4617 10248 4629 10251
rect 4488 10220 4629 10248
rect 4488 10208 4494 10220
rect 4617 10217 4629 10220
rect 4663 10217 4675 10251
rect 4617 10211 4675 10217
rect 4893 10251 4951 10257
rect 4893 10217 4905 10251
rect 4939 10248 4951 10251
rect 5166 10248 5172 10260
rect 4939 10220 5172 10248
rect 4939 10217 4951 10220
rect 4893 10211 4951 10217
rect 5166 10208 5172 10220
rect 5224 10208 5230 10260
rect 5261 10251 5319 10257
rect 5261 10217 5273 10251
rect 5307 10248 5319 10251
rect 8110 10248 8116 10260
rect 5307 10220 8116 10248
rect 5307 10217 5319 10220
rect 5261 10211 5319 10217
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 8202 10208 8208 10260
rect 8260 10248 8266 10260
rect 9122 10248 9128 10260
rect 8260 10220 9128 10248
rect 8260 10208 8266 10220
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 11974 10248 11980 10260
rect 9640 10220 9720 10248
rect 11935 10220 11980 10248
rect 9640 10208 9646 10220
rect 1397 10183 1455 10189
rect 1397 10149 1409 10183
rect 1443 10180 1455 10183
rect 2130 10180 2136 10192
rect 1443 10152 2136 10180
rect 1443 10149 1455 10152
rect 1397 10143 1455 10149
rect 2130 10140 2136 10152
rect 2188 10140 2194 10192
rect 3970 10140 3976 10192
rect 4028 10180 4034 10192
rect 5534 10180 5540 10192
rect 4028 10152 5540 10180
rect 4028 10140 4034 10152
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 7650 10180 7656 10192
rect 5920 10152 7656 10180
rect 2317 10115 2375 10121
rect 2317 10081 2329 10115
rect 2363 10112 2375 10115
rect 2958 10112 2964 10124
rect 2363 10084 2964 10112
rect 2363 10081 2375 10084
rect 2317 10075 2375 10081
rect 2958 10072 2964 10084
rect 3016 10072 3022 10124
rect 3142 10072 3148 10124
rect 3200 10112 3206 10124
rect 3329 10115 3387 10121
rect 3329 10112 3341 10115
rect 3200 10084 3341 10112
rect 3200 10072 3206 10084
rect 3329 10081 3341 10084
rect 3375 10081 3387 10115
rect 3329 10075 3387 10081
rect 3418 10072 3424 10124
rect 3476 10112 3482 10124
rect 4065 10115 4123 10121
rect 3476 10084 3521 10112
rect 3476 10072 3482 10084
rect 4065 10081 4077 10115
rect 4111 10081 4123 10115
rect 4065 10075 4123 10081
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10112 4859 10115
rect 5810 10112 5816 10124
rect 4847 10084 5816 10112
rect 4847 10081 4859 10084
rect 4801 10075 4859 10081
rect 2498 10044 2504 10056
rect 2459 10016 2504 10044
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 3510 10044 3516 10056
rect 3471 10016 3516 10044
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 4080 10044 4108 10075
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 5920 10121 5948 10152
rect 7650 10140 7656 10152
rect 7708 10140 7714 10192
rect 8938 10180 8944 10192
rect 7944 10152 8944 10180
rect 5905 10115 5963 10121
rect 5905 10081 5917 10115
rect 5951 10081 5963 10115
rect 5905 10075 5963 10081
rect 6172 10115 6230 10121
rect 6172 10081 6184 10115
rect 6218 10112 6230 10115
rect 7466 10112 7472 10124
rect 6218 10084 7472 10112
rect 6218 10081 6230 10084
rect 6172 10075 6230 10081
rect 7466 10072 7472 10084
rect 7524 10072 7530 10124
rect 5350 10044 5356 10056
rect 4080 10016 5120 10044
rect 5311 10016 5356 10044
rect 4154 9936 4160 9988
rect 4212 9976 4218 9988
rect 4890 9976 4896 9988
rect 4212 9948 4896 9976
rect 4212 9936 4218 9948
rect 4890 9936 4896 9948
rect 4948 9936 4954 9988
rect 1578 9868 1584 9920
rect 1636 9908 1642 9920
rect 1857 9911 1915 9917
rect 1857 9908 1869 9911
rect 1636 9880 1869 9908
rect 1636 9868 1642 9880
rect 1857 9877 1869 9880
rect 1903 9877 1915 9911
rect 4246 9908 4252 9920
rect 4207 9880 4252 9908
rect 1857 9871 1915 9877
rect 4246 9868 4252 9880
rect 4304 9868 4310 9920
rect 5092 9908 5120 10016
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10013 5503 10047
rect 7944 10044 7972 10152
rect 8938 10140 8944 10152
rect 8996 10140 9002 10192
rect 9692 10121 9720 10220
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 12250 10248 12256 10260
rect 12211 10220 12256 10248
rect 12250 10208 12256 10220
rect 12308 10208 12314 10260
rect 13262 10248 13268 10260
rect 13223 10220 13268 10248
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 13446 10208 13452 10260
rect 13504 10248 13510 10260
rect 13725 10251 13783 10257
rect 13725 10248 13737 10251
rect 13504 10220 13737 10248
rect 13504 10208 13510 10220
rect 13725 10217 13737 10220
rect 13771 10217 13783 10251
rect 14274 10248 14280 10260
rect 14235 10220 14280 10248
rect 13725 10211 13783 10217
rect 14274 10208 14280 10220
rect 14332 10208 14338 10260
rect 15749 10251 15807 10257
rect 15749 10217 15761 10251
rect 15795 10248 15807 10251
rect 16206 10248 16212 10260
rect 15795 10220 16212 10248
rect 15795 10217 15807 10220
rect 15749 10211 15807 10217
rect 16206 10208 16212 10220
rect 16264 10248 16270 10260
rect 16666 10248 16672 10260
rect 16264 10220 16672 10248
rect 16264 10208 16270 10220
rect 16666 10208 16672 10220
rect 16724 10208 16730 10260
rect 17678 10208 17684 10260
rect 17736 10248 17742 10260
rect 18325 10251 18383 10257
rect 18325 10248 18337 10251
rect 17736 10220 18337 10248
rect 17736 10208 17742 10220
rect 18325 10217 18337 10220
rect 18371 10217 18383 10251
rect 18325 10211 18383 10217
rect 9944 10183 10002 10189
rect 9944 10149 9956 10183
rect 9990 10180 10002 10183
rect 10318 10180 10324 10192
rect 9990 10152 10324 10180
rect 9990 10149 10002 10152
rect 9944 10143 10002 10149
rect 10318 10140 10324 10152
rect 10376 10180 10382 10192
rect 10686 10180 10692 10192
rect 10376 10152 10692 10180
rect 10376 10140 10382 10152
rect 10686 10140 10692 10152
rect 10744 10140 10750 10192
rect 11146 10140 11152 10192
rect 11204 10180 11210 10192
rect 13464 10180 13492 10208
rect 11204 10152 13492 10180
rect 11204 10140 11210 10152
rect 13538 10140 13544 10192
rect 13596 10180 13602 10192
rect 13633 10183 13691 10189
rect 13633 10180 13645 10183
rect 13596 10152 13645 10180
rect 13596 10140 13602 10152
rect 13633 10149 13645 10152
rect 13679 10149 13691 10183
rect 13633 10143 13691 10149
rect 15657 10183 15715 10189
rect 15657 10149 15669 10183
rect 15703 10180 15715 10183
rect 16114 10180 16120 10192
rect 15703 10152 16120 10180
rect 15703 10149 15715 10152
rect 15657 10143 15715 10149
rect 8021 10115 8079 10121
rect 8021 10081 8033 10115
rect 8067 10112 8079 10115
rect 9677 10115 9735 10121
rect 8067 10084 8892 10112
rect 8067 10081 8079 10084
rect 8021 10075 8079 10081
rect 5445 10007 5503 10013
rect 7208 10016 7972 10044
rect 8113 10047 8171 10053
rect 5166 9936 5172 9988
rect 5224 9976 5230 9988
rect 5460 9976 5488 10007
rect 5224 9948 5488 9976
rect 5224 9936 5230 9948
rect 7208 9908 7236 10016
rect 8113 10013 8125 10047
rect 8159 10013 8171 10047
rect 8113 10007 8171 10013
rect 7285 9979 7343 9985
rect 7285 9945 7297 9979
rect 7331 9976 7343 9979
rect 8018 9976 8024 9988
rect 7331 9948 8024 9976
rect 7331 9945 7343 9948
rect 7285 9939 7343 9945
rect 8018 9936 8024 9948
rect 8076 9936 8082 9988
rect 8128 9976 8156 10007
rect 8202 10004 8208 10056
rect 8260 10044 8266 10056
rect 8662 10044 8668 10056
rect 8260 10016 8305 10044
rect 8404 10016 8524 10044
rect 8623 10016 8668 10044
rect 8260 10004 8266 10016
rect 8404 9976 8432 10016
rect 8128 9948 8432 9976
rect 8496 9976 8524 10016
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 8864 10044 8892 10084
rect 9677 10081 9689 10115
rect 9723 10081 9735 10115
rect 12158 10112 12164 10124
rect 12119 10084 12164 10112
rect 9677 10075 9735 10081
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 12618 10072 12624 10124
rect 12676 10112 12682 10124
rect 13648 10112 13676 10143
rect 16114 10140 16120 10152
rect 16172 10180 16178 10192
rect 16482 10180 16488 10192
rect 16172 10152 16488 10180
rect 16172 10140 16178 10152
rect 16482 10140 16488 10152
rect 16540 10140 16546 10192
rect 16574 10140 16580 10192
rect 16632 10180 16638 10192
rect 17954 10180 17960 10192
rect 16632 10152 17960 10180
rect 16632 10140 16638 10152
rect 17954 10140 17960 10152
rect 18012 10140 18018 10192
rect 12676 10084 12721 10112
rect 13648 10084 16252 10112
rect 12676 10072 12682 10084
rect 9490 10044 9496 10056
rect 8864 10016 9496 10044
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 12713 10047 12771 10053
rect 12713 10013 12725 10047
rect 12759 10013 12771 10047
rect 12713 10007 12771 10013
rect 8754 9976 8760 9988
rect 8496 9948 8760 9976
rect 8754 9936 8760 9948
rect 8812 9936 8818 9988
rect 12618 9936 12624 9988
rect 12676 9976 12682 9988
rect 12728 9976 12756 10007
rect 12802 10004 12808 10056
rect 12860 10044 12866 10056
rect 13906 10044 13912 10056
rect 12860 10016 12905 10044
rect 13867 10016 13912 10044
rect 12860 10004 12866 10016
rect 13906 10004 13912 10016
rect 13964 10004 13970 10056
rect 14826 10004 14832 10056
rect 14884 10044 14890 10056
rect 15887 10047 15945 10053
rect 15887 10044 15899 10047
rect 14884 10016 15899 10044
rect 14884 10004 14890 10016
rect 15887 10013 15899 10016
rect 15933 10013 15945 10047
rect 16224 10044 16252 10084
rect 16298 10072 16304 10124
rect 16356 10112 16362 10124
rect 16945 10115 17003 10121
rect 16945 10112 16957 10115
rect 16356 10084 16957 10112
rect 16356 10072 16362 10084
rect 16945 10081 16957 10084
rect 16991 10081 17003 10115
rect 16945 10075 17003 10081
rect 17212 10115 17270 10121
rect 17212 10081 17224 10115
rect 17258 10112 17270 10115
rect 17494 10112 17500 10124
rect 17258 10084 17500 10112
rect 17258 10081 17270 10084
rect 17212 10075 17270 10081
rect 17494 10072 17500 10084
rect 17552 10072 17558 10124
rect 16224 10016 16988 10044
rect 15887 10007 15945 10013
rect 12676 9948 12756 9976
rect 12676 9936 12682 9948
rect 13814 9936 13820 9988
rect 13872 9976 13878 9988
rect 14182 9976 14188 9988
rect 13872 9948 14188 9976
rect 13872 9936 13878 9948
rect 14182 9936 14188 9948
rect 14240 9936 14246 9988
rect 5092 9880 7236 9908
rect 7653 9911 7711 9917
rect 7653 9877 7665 9911
rect 7699 9908 7711 9911
rect 8294 9908 8300 9920
rect 7699 9880 8300 9908
rect 7699 9877 7711 9880
rect 7653 9871 7711 9877
rect 8294 9868 8300 9880
rect 8352 9868 8358 9920
rect 11054 9908 11060 9920
rect 10967 9880 11060 9908
rect 11054 9868 11060 9880
rect 11112 9908 11118 9920
rect 11974 9908 11980 9920
rect 11112 9880 11980 9908
rect 11112 9868 11118 9880
rect 11974 9868 11980 9880
rect 12032 9868 12038 9920
rect 15286 9908 15292 9920
rect 15247 9880 15292 9908
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 16960 9908 16988 10016
rect 17954 9908 17960 9920
rect 16960 9880 17960 9908
rect 17954 9868 17960 9880
rect 18012 9868 18018 9920
rect 1104 9818 18860 9840
rect 1104 9766 3947 9818
rect 3999 9766 4011 9818
rect 4063 9766 4075 9818
rect 4127 9766 4139 9818
rect 4191 9766 9878 9818
rect 9930 9766 9942 9818
rect 9994 9766 10006 9818
rect 10058 9766 10070 9818
rect 10122 9766 15808 9818
rect 15860 9766 15872 9818
rect 15924 9766 15936 9818
rect 15988 9766 16000 9818
rect 16052 9766 18860 9818
rect 1104 9744 18860 9766
rect 8294 9704 8300 9716
rect 3620 9676 8300 9704
rect 1504 9540 2176 9568
rect 1504 9509 1532 9540
rect 1489 9503 1547 9509
rect 1489 9469 1501 9503
rect 1535 9469 1547 9503
rect 2038 9500 2044 9512
rect 1999 9472 2044 9500
rect 1489 9463 1547 9469
rect 2038 9460 2044 9472
rect 2096 9460 2102 9512
rect 2148 9500 2176 9540
rect 3050 9500 3056 9512
rect 2148 9472 3056 9500
rect 3050 9460 3056 9472
rect 3108 9500 3114 9512
rect 3620 9500 3648 9676
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 8386 9664 8392 9716
rect 8444 9704 8450 9716
rect 11422 9704 11428 9716
rect 8444 9676 11428 9704
rect 8444 9664 8450 9676
rect 11422 9664 11428 9676
rect 11480 9664 11486 9716
rect 11698 9664 11704 9716
rect 11756 9704 11762 9716
rect 11756 9676 13860 9704
rect 11756 9664 11762 9676
rect 3697 9639 3755 9645
rect 3697 9605 3709 9639
rect 3743 9636 3755 9639
rect 5074 9636 5080 9648
rect 3743 9608 5080 9636
rect 3743 9605 3755 9608
rect 3697 9599 3755 9605
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 5718 9636 5724 9648
rect 5679 9608 5724 9636
rect 5718 9596 5724 9608
rect 5776 9596 5782 9648
rect 8018 9636 8024 9648
rect 6380 9608 8024 9636
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9568 4399 9571
rect 5166 9568 5172 9580
rect 4387 9540 5172 9568
rect 4387 9537 4399 9540
rect 4341 9531 4399 9537
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 5353 9571 5411 9577
rect 5353 9537 5365 9571
rect 5399 9568 5411 9571
rect 6270 9568 6276 9580
rect 5399 9540 6276 9568
rect 5399 9537 5411 9540
rect 5353 9531 5411 9537
rect 5736 9512 5764 9540
rect 6270 9528 6276 9540
rect 6328 9528 6334 9580
rect 6380 9577 6408 9608
rect 8018 9596 8024 9608
rect 8076 9636 8082 9648
rect 9306 9636 9312 9648
rect 8076 9608 9159 9636
rect 9267 9608 9312 9636
rect 8076 9596 8082 9608
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9537 6423 9571
rect 7282 9568 7288 9580
rect 7243 9540 7288 9568
rect 6365 9531 6423 9537
rect 7282 9528 7288 9540
rect 7340 9528 7346 9580
rect 7466 9568 7472 9580
rect 7427 9540 7472 9568
rect 7466 9528 7472 9540
rect 7524 9568 7530 9580
rect 8202 9568 8208 9580
rect 7524 9540 8208 9568
rect 7524 9528 7530 9540
rect 8202 9528 8208 9540
rect 8260 9568 8266 9580
rect 9033 9571 9091 9577
rect 9033 9568 9045 9571
rect 8260 9540 9045 9568
rect 8260 9528 8266 9540
rect 9033 9537 9045 9540
rect 9079 9537 9091 9571
rect 9131 9568 9159 9608
rect 9306 9596 9312 9608
rect 9364 9596 9370 9648
rect 10137 9639 10195 9645
rect 9416 9608 9904 9636
rect 9416 9568 9444 9608
rect 9131 9540 9444 9568
rect 9033 9531 9091 9537
rect 9490 9528 9496 9580
rect 9548 9568 9554 9580
rect 9876 9577 9904 9608
rect 10137 9605 10149 9639
rect 10183 9636 10195 9639
rect 10226 9636 10232 9648
rect 10183 9608 10232 9636
rect 10183 9605 10195 9608
rect 10137 9599 10195 9605
rect 10226 9596 10232 9608
rect 10284 9596 10290 9648
rect 13832 9645 13860 9676
rect 14182 9664 14188 9716
rect 14240 9704 14246 9716
rect 16298 9704 16304 9716
rect 14240 9676 16304 9704
rect 14240 9664 14246 9676
rect 16298 9664 16304 9676
rect 16356 9664 16362 9716
rect 12161 9639 12219 9645
rect 12161 9636 12173 9639
rect 10520 9608 12173 9636
rect 9769 9571 9827 9577
rect 9769 9568 9781 9571
rect 9548 9540 9781 9568
rect 9548 9528 9554 9540
rect 9769 9537 9781 9540
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9537 9919 9571
rect 9861 9531 9919 9537
rect 3108 9472 3648 9500
rect 4065 9503 4123 9509
rect 3108 9460 3114 9472
rect 4065 9469 4077 9503
rect 4111 9500 4123 9503
rect 5442 9500 5448 9512
rect 4111 9472 5448 9500
rect 4111 9469 4123 9472
rect 4065 9463 4123 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 5718 9460 5724 9512
rect 5776 9460 5782 9512
rect 7558 9460 7564 9512
rect 7616 9500 7622 9512
rect 8021 9503 8079 9509
rect 8021 9500 8033 9503
rect 7616 9472 8033 9500
rect 7616 9460 7622 9472
rect 8021 9469 8033 9472
rect 8067 9500 8079 9503
rect 8386 9500 8392 9512
rect 8067 9472 8392 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 8662 9460 8668 9512
rect 8720 9500 8726 9512
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 8720 9472 8861 9500
rect 8720 9460 8726 9472
rect 8849 9469 8861 9472
rect 8895 9469 8907 9503
rect 8849 9463 8907 9469
rect 8938 9460 8944 9512
rect 8996 9500 9002 9512
rect 8996 9472 9041 9500
rect 8996 9460 9002 9472
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 10520 9509 10548 9608
rect 12161 9605 12173 9608
rect 12207 9605 12219 9639
rect 12161 9599 12219 9605
rect 13817 9639 13875 9645
rect 13817 9605 13829 9639
rect 13863 9636 13875 9639
rect 13906 9636 13912 9648
rect 13863 9608 13912 9636
rect 13863 9605 13875 9608
rect 13817 9599 13875 9605
rect 13906 9596 13912 9608
rect 13964 9596 13970 9648
rect 10686 9568 10692 9580
rect 10647 9540 10692 9568
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 11698 9528 11704 9580
rect 11756 9568 11762 9580
rect 14200 9577 14228 9664
rect 11885 9571 11943 9577
rect 11885 9568 11897 9571
rect 11756 9540 11897 9568
rect 11756 9528 11762 9540
rect 11885 9537 11897 9540
rect 11931 9537 11943 9571
rect 14185 9571 14243 9577
rect 11885 9531 11943 9537
rect 11992 9540 12572 9568
rect 10505 9503 10563 9509
rect 10505 9500 10517 9503
rect 9180 9472 10517 9500
rect 9180 9460 9186 9472
rect 10505 9469 10517 9472
rect 10551 9469 10563 9503
rect 11992 9500 12020 9540
rect 10505 9463 10563 9469
rect 10971 9472 12020 9500
rect 2308 9435 2366 9441
rect 2308 9401 2320 9435
rect 2354 9432 2366 9435
rect 2498 9432 2504 9444
rect 2354 9404 2504 9432
rect 2354 9401 2366 9404
rect 2308 9395 2366 9401
rect 2498 9392 2504 9404
rect 2556 9392 2562 9444
rect 4338 9392 4344 9444
rect 4396 9432 4402 9444
rect 5169 9435 5227 9441
rect 5169 9432 5181 9435
rect 4396 9404 5181 9432
rect 4396 9392 4402 9404
rect 5169 9401 5181 9404
rect 5215 9432 5227 9435
rect 5258 9432 5264 9444
rect 5215 9404 5264 9432
rect 5215 9401 5227 9404
rect 5169 9395 5227 9401
rect 5258 9392 5264 9404
rect 5316 9392 5322 9444
rect 6089 9435 6147 9441
rect 6089 9401 6101 9435
rect 6135 9432 6147 9435
rect 6135 9404 7696 9432
rect 6135 9401 6147 9404
rect 6089 9395 6147 9401
rect 1673 9367 1731 9373
rect 1673 9333 1685 9367
rect 1719 9364 1731 9367
rect 3050 9364 3056 9376
rect 1719 9336 3056 9364
rect 1719 9333 1731 9336
rect 1673 9327 1731 9333
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 3421 9367 3479 9373
rect 3421 9333 3433 9367
rect 3467 9364 3479 9367
rect 3510 9364 3516 9376
rect 3467 9336 3516 9364
rect 3467 9333 3479 9336
rect 3421 9327 3479 9333
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 4157 9367 4215 9373
rect 4157 9333 4169 9367
rect 4203 9364 4215 9367
rect 4709 9367 4767 9373
rect 4709 9364 4721 9367
rect 4203 9336 4721 9364
rect 4203 9333 4215 9336
rect 4157 9327 4215 9333
rect 4709 9333 4721 9336
rect 4755 9333 4767 9367
rect 4709 9327 4767 9333
rect 4798 9324 4804 9376
rect 4856 9364 4862 9376
rect 5077 9367 5135 9373
rect 5077 9364 5089 9367
rect 4856 9336 5089 9364
rect 4856 9324 4862 9336
rect 5077 9333 5089 9336
rect 5123 9364 5135 9367
rect 5626 9364 5632 9376
rect 5123 9336 5632 9364
rect 5123 9333 5135 9336
rect 5077 9327 5135 9333
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 6181 9367 6239 9373
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 6825 9367 6883 9373
rect 6825 9364 6837 9367
rect 6227 9336 6837 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 6825 9333 6837 9336
rect 6871 9333 6883 9367
rect 6825 9327 6883 9333
rect 7193 9367 7251 9373
rect 7193 9333 7205 9367
rect 7239 9364 7251 9367
rect 7282 9364 7288 9376
rect 7239 9336 7288 9364
rect 7239 9333 7251 9336
rect 7193 9327 7251 9333
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 7668 9373 7696 9404
rect 7926 9392 7932 9444
rect 7984 9432 7990 9444
rect 9677 9435 9735 9441
rect 9677 9432 9689 9435
rect 7984 9404 8432 9432
rect 7984 9392 7990 9404
rect 8404 9376 8432 9404
rect 9232 9404 9689 9432
rect 7653 9367 7711 9373
rect 7653 9333 7665 9367
rect 7699 9333 7711 9367
rect 7653 9327 7711 9333
rect 8018 9324 8024 9376
rect 8076 9364 8082 9376
rect 8113 9367 8171 9373
rect 8113 9364 8125 9367
rect 8076 9336 8125 9364
rect 8076 9324 8082 9336
rect 8113 9333 8125 9336
rect 8159 9333 8171 9367
rect 8113 9327 8171 9333
rect 8386 9324 8392 9376
rect 8444 9324 8450 9376
rect 8481 9367 8539 9373
rect 8481 9333 8493 9367
rect 8527 9364 8539 9367
rect 9232 9364 9260 9404
rect 9677 9401 9689 9404
rect 9723 9401 9735 9435
rect 9677 9395 9735 9401
rect 9858 9392 9864 9444
rect 9916 9432 9922 9444
rect 10410 9432 10416 9444
rect 9916 9404 10416 9432
rect 9916 9392 9922 9404
rect 10410 9392 10416 9404
rect 10468 9392 10474 9444
rect 8527 9336 9260 9364
rect 8527 9333 8539 9336
rect 8481 9327 8539 9333
rect 9490 9324 9496 9376
rect 9548 9364 9554 9376
rect 10597 9367 10655 9373
rect 10597 9364 10609 9367
rect 9548 9336 10609 9364
rect 9548 9324 9554 9336
rect 10597 9333 10609 9336
rect 10643 9333 10655 9367
rect 10597 9327 10655 9333
rect 10870 9324 10876 9376
rect 10928 9364 10934 9376
rect 10971 9364 10999 9472
rect 12342 9460 12348 9512
rect 12400 9500 12406 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 12400 9472 12449 9500
rect 12400 9460 12406 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12544 9500 12572 9540
rect 14185 9537 14197 9571
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9568 17095 9571
rect 17678 9568 17684 9580
rect 17083 9540 17684 9568
rect 17083 9537 17095 9540
rect 17037 9531 17095 9537
rect 17678 9528 17684 9540
rect 17736 9528 17742 9580
rect 14452 9503 14510 9509
rect 12544 9472 12848 9500
rect 12437 9463 12495 9469
rect 11701 9435 11759 9441
rect 11701 9401 11713 9435
rect 11747 9432 11759 9435
rect 11882 9432 11888 9444
rect 11747 9404 11888 9432
rect 11747 9401 11759 9404
rect 11701 9395 11759 9401
rect 11882 9392 11888 9404
rect 11940 9392 11946 9444
rect 12161 9435 12219 9441
rect 12161 9401 12173 9435
rect 12207 9432 12219 9435
rect 12250 9432 12256 9444
rect 12207 9404 12256 9432
rect 12207 9401 12219 9404
rect 12161 9395 12219 9401
rect 12250 9392 12256 9404
rect 12308 9392 12314 9444
rect 12710 9441 12716 9444
rect 12704 9432 12716 9441
rect 12671 9404 12716 9432
rect 12704 9395 12716 9404
rect 12710 9392 12716 9395
rect 12768 9392 12774 9444
rect 12820 9432 12848 9472
rect 14452 9469 14464 9503
rect 14498 9500 14510 9503
rect 14826 9500 14832 9512
rect 14498 9472 14832 9500
rect 14498 9469 14510 9472
rect 14452 9463 14510 9469
rect 14826 9460 14832 9472
rect 14884 9460 14890 9512
rect 15010 9460 15016 9512
rect 15068 9500 15074 9512
rect 16761 9503 16819 9509
rect 16761 9500 16773 9503
rect 15068 9472 16773 9500
rect 15068 9460 15074 9472
rect 16761 9469 16773 9472
rect 16807 9469 16819 9503
rect 16761 9463 16819 9469
rect 15654 9432 15660 9444
rect 12820 9404 15660 9432
rect 15654 9392 15660 9404
rect 15712 9392 15718 9444
rect 16114 9392 16120 9444
rect 16172 9432 16178 9444
rect 18138 9432 18144 9444
rect 16172 9404 18144 9432
rect 16172 9392 16178 9404
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 11330 9364 11336 9376
rect 10928 9336 10999 9364
rect 11291 9336 11336 9364
rect 10928 9324 10934 9336
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 11793 9367 11851 9373
rect 11793 9333 11805 9367
rect 11839 9364 11851 9367
rect 12434 9364 12440 9376
rect 11839 9336 12440 9364
rect 11839 9333 11851 9336
rect 11793 9327 11851 9333
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 14826 9324 14832 9376
rect 14884 9364 14890 9376
rect 15565 9367 15623 9373
rect 15565 9364 15577 9367
rect 14884 9336 15577 9364
rect 14884 9324 14890 9336
rect 15565 9333 15577 9336
rect 15611 9333 15623 9367
rect 15565 9327 15623 9333
rect 16393 9367 16451 9373
rect 16393 9333 16405 9367
rect 16439 9364 16451 9367
rect 16666 9364 16672 9376
rect 16439 9336 16672 9364
rect 16439 9333 16451 9336
rect 16393 9327 16451 9333
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 16850 9324 16856 9376
rect 16908 9364 16914 9376
rect 16908 9336 16953 9364
rect 16908 9324 16914 9336
rect 1104 9274 18860 9296
rect 1104 9222 6912 9274
rect 6964 9222 6976 9274
rect 7028 9222 7040 9274
rect 7092 9222 7104 9274
rect 7156 9222 12843 9274
rect 12895 9222 12907 9274
rect 12959 9222 12971 9274
rect 13023 9222 13035 9274
rect 13087 9222 18860 9274
rect 1104 9200 18860 9222
rect 7285 9163 7343 9169
rect 1412 9132 7236 9160
rect 1412 9033 1440 9132
rect 2409 9095 2467 9101
rect 2409 9061 2421 9095
rect 2455 9092 2467 9095
rect 2498 9092 2504 9104
rect 2455 9064 2504 9092
rect 2455 9061 2467 9064
rect 2409 9055 2467 9061
rect 2498 9052 2504 9064
rect 2556 9052 2562 9104
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 4706 9092 4712 9104
rect 4120 9064 4712 9092
rect 4120 9052 4126 9064
rect 4706 9052 4712 9064
rect 4764 9092 4770 9104
rect 5258 9092 5264 9104
rect 4764 9064 5264 9092
rect 4764 9052 4770 9064
rect 5258 9052 5264 9064
rect 5316 9052 5322 9104
rect 5902 9052 5908 9104
rect 5960 9101 5966 9104
rect 5960 9095 6024 9101
rect 5960 9061 5978 9095
rect 6012 9061 6024 9095
rect 7208 9092 7236 9132
rect 7285 9129 7297 9163
rect 7331 9160 7343 9163
rect 7466 9160 7472 9172
rect 7331 9132 7472 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 8202 9120 8208 9172
rect 8260 9160 8266 9172
rect 8757 9163 8815 9169
rect 8757 9160 8769 9163
rect 8260 9132 8769 9160
rect 8260 9120 8266 9132
rect 8757 9129 8769 9132
rect 8803 9129 8815 9163
rect 10045 9163 10103 9169
rect 10045 9160 10057 9163
rect 8757 9123 8815 9129
rect 8864 9132 10057 9160
rect 7208 9064 7512 9092
rect 5960 9055 6024 9061
rect 5960 9052 5966 9055
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 8993 1455 9027
rect 1397 8987 1455 8993
rect 2314 8984 2320 9036
rect 2372 9024 2378 9036
rect 2372 8996 2417 9024
rect 2372 8984 2378 8996
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 3329 9027 3387 9033
rect 3329 9024 3341 9027
rect 2832 8996 3341 9024
rect 2832 8984 2838 8996
rect 3329 8993 3341 8996
rect 3375 8993 3387 9027
rect 4321 9027 4379 9033
rect 4321 9024 4333 9027
rect 3329 8987 3387 8993
rect 3528 8996 4333 9024
rect 3528 8968 3556 8996
rect 4321 8993 4333 8996
rect 4367 8993 4379 9027
rect 4321 8987 4379 8993
rect 5721 9027 5779 9033
rect 5721 8993 5733 9027
rect 5767 9024 5779 9027
rect 7285 9027 7343 9033
rect 7285 9024 7297 9027
rect 5767 8996 7297 9024
rect 5767 8993 5779 8996
rect 5721 8987 5779 8993
rect 7285 8993 7297 8996
rect 7331 9024 7343 9027
rect 7377 9027 7435 9033
rect 7377 9024 7389 9027
rect 7331 8996 7389 9024
rect 7331 8993 7343 8996
rect 7285 8987 7343 8993
rect 7377 8993 7389 8996
rect 7423 8993 7435 9027
rect 7484 9024 7512 9064
rect 7558 9052 7564 9104
rect 7616 9101 7622 9104
rect 7616 9095 7680 9101
rect 7616 9061 7634 9095
rect 7668 9061 7680 9095
rect 7616 9055 7680 9061
rect 7616 9052 7622 9055
rect 8018 9052 8024 9104
rect 8076 9092 8082 9104
rect 8864 9092 8892 9132
rect 10045 9129 10057 9132
rect 10091 9160 10103 9163
rect 10091 9132 11284 9160
rect 10091 9129 10103 9132
rect 10045 9123 10103 9129
rect 10137 9095 10195 9101
rect 10137 9092 10149 9095
rect 8076 9064 8892 9092
rect 10060 9064 10149 9092
rect 8076 9052 8082 9064
rect 10060 9036 10088 9064
rect 10137 9061 10149 9064
rect 10183 9061 10195 9095
rect 11146 9092 11152 9104
rect 10137 9055 10195 9061
rect 10520 9064 11152 9092
rect 7484 8996 8432 9024
rect 7377 8987 7435 8993
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8925 2559 8959
rect 3418 8956 3424 8968
rect 3379 8928 3424 8956
rect 2501 8919 2559 8925
rect 1581 8891 1639 8897
rect 1581 8857 1593 8891
rect 1627 8888 1639 8891
rect 1627 8860 2176 8888
rect 1627 8857 1639 8860
rect 1581 8851 1639 8857
rect 1946 8820 1952 8832
rect 1907 8792 1952 8820
rect 1946 8780 1952 8792
rect 2004 8780 2010 8832
rect 2148 8820 2176 8860
rect 2406 8848 2412 8900
rect 2464 8888 2470 8900
rect 2516 8888 2544 8919
rect 3418 8916 3424 8928
rect 3476 8916 3482 8968
rect 3510 8916 3516 8968
rect 3568 8956 3574 8968
rect 4065 8959 4123 8965
rect 3568 8928 3613 8956
rect 3568 8916 3574 8928
rect 4065 8925 4077 8959
rect 4111 8925 4123 8959
rect 8404 8956 8432 8996
rect 8478 8984 8484 9036
rect 8536 9024 8542 9036
rect 9582 9024 9588 9036
rect 8536 8996 9588 9024
rect 8536 8984 8542 8996
rect 9582 8984 9588 8996
rect 9640 8984 9646 9036
rect 10042 8984 10048 9036
rect 10100 8984 10106 9036
rect 10520 9024 10548 9064
rect 11146 9052 11152 9064
rect 11204 9052 11210 9104
rect 10152 8996 10548 9024
rect 10152 8956 10180 8996
rect 10686 8984 10692 9036
rect 10744 9024 10750 9036
rect 10870 9024 10876 9036
rect 10744 8996 10876 9024
rect 10744 8984 10750 8996
rect 10870 8984 10876 8996
rect 10928 8984 10934 9036
rect 11256 9024 11284 9132
rect 11330 9120 11336 9172
rect 11388 9160 11394 9172
rect 11793 9163 11851 9169
rect 11793 9160 11805 9163
rect 11388 9132 11805 9160
rect 11388 9120 11394 9132
rect 11793 9129 11805 9132
rect 11839 9129 11851 9163
rect 11793 9123 11851 9129
rect 11882 9120 11888 9172
rect 11940 9160 11946 9172
rect 12345 9163 12403 9169
rect 12345 9160 12357 9163
rect 11940 9132 12357 9160
rect 11940 9120 11946 9132
rect 12345 9129 12357 9132
rect 12391 9129 12403 9163
rect 12345 9123 12403 9129
rect 12713 9163 12771 9169
rect 12713 9129 12725 9163
rect 12759 9160 12771 9163
rect 13173 9163 13231 9169
rect 13173 9160 13185 9163
rect 12759 9132 13185 9160
rect 12759 9129 12771 9132
rect 12713 9123 12771 9129
rect 13173 9129 13185 9132
rect 13219 9129 13231 9163
rect 13173 9123 13231 9129
rect 14645 9163 14703 9169
rect 14645 9129 14657 9163
rect 14691 9160 14703 9163
rect 15286 9160 15292 9172
rect 14691 9132 15292 9160
rect 14691 9129 14703 9132
rect 14645 9123 14703 9129
rect 11701 9095 11759 9101
rect 11701 9061 11713 9095
rect 11747 9092 11759 9095
rect 12526 9092 12532 9104
rect 11747 9064 12532 9092
rect 11747 9061 11759 9064
rect 11701 9055 11759 9061
rect 12526 9052 12532 9064
rect 12584 9052 12590 9104
rect 12728 9024 12756 9123
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 16298 9120 16304 9172
rect 16356 9120 16362 9172
rect 17494 9160 17500 9172
rect 17455 9132 17500 9160
rect 17494 9120 17500 9132
rect 17552 9120 17558 9172
rect 12805 9095 12863 9101
rect 12805 9061 12817 9095
rect 12851 9092 12863 9095
rect 15010 9092 15016 9104
rect 12851 9064 15016 9092
rect 12851 9061 12863 9064
rect 12805 9055 12863 9061
rect 11256 8996 12756 9024
rect 10318 8956 10324 8968
rect 8404 8928 10180 8956
rect 10279 8928 10324 8956
rect 4065 8919 4123 8925
rect 2464 8860 2544 8888
rect 2464 8848 2470 8860
rect 2590 8848 2596 8900
rect 2648 8888 2654 8900
rect 4080 8888 4108 8919
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 10410 8916 10416 8968
rect 10468 8956 10474 8968
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 10468 8928 10977 8956
rect 10468 8916 10474 8928
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 11146 8956 11152 8968
rect 11107 8928 11152 8956
rect 10965 8919 11023 8925
rect 11146 8916 11152 8928
rect 11204 8916 11210 8968
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8956 12035 8959
rect 12066 8956 12072 8968
rect 12023 8928 12072 8956
rect 12023 8925 12035 8928
rect 11977 8919 12035 8925
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 12342 8916 12348 8968
rect 12400 8956 12406 8968
rect 12820 8956 12848 9055
rect 15010 9052 15016 9064
rect 15068 9052 15074 9104
rect 16316 9092 16344 9120
rect 16132 9064 16344 9092
rect 16132 9036 16160 9064
rect 13998 8984 14004 9036
rect 14056 9024 14062 9036
rect 14182 9024 14188 9036
rect 14056 8996 14188 9024
rect 14056 8984 14062 8996
rect 14182 8984 14188 8996
rect 14240 9024 14246 9036
rect 14553 9027 14611 9033
rect 14553 9024 14565 9027
rect 14240 8996 14565 9024
rect 14240 8984 14246 8996
rect 14553 8993 14565 8996
rect 14599 8993 14611 9027
rect 16114 9024 16120 9036
rect 16027 8996 16120 9024
rect 14553 8987 14611 8993
rect 16114 8984 16120 8996
rect 16172 8984 16178 9036
rect 16384 9027 16442 9033
rect 16384 8993 16396 9027
rect 16430 9024 16442 9027
rect 17126 9024 17132 9036
rect 16430 8996 17132 9024
rect 16430 8993 16442 8996
rect 16384 8987 16442 8993
rect 17126 8984 17132 8996
rect 17184 8984 17190 9036
rect 12400 8928 12848 8956
rect 12897 8959 12955 8965
rect 12400 8916 12406 8928
rect 12897 8925 12909 8959
rect 12943 8925 12955 8959
rect 13354 8956 13360 8968
rect 13315 8928 13360 8956
rect 12897 8919 12955 8925
rect 2648 8860 4108 8888
rect 2648 8848 2654 8860
rect 2866 8820 2872 8832
rect 2148 8792 2872 8820
rect 2866 8780 2872 8792
rect 2924 8780 2930 8832
rect 2961 8823 3019 8829
rect 2961 8789 2973 8823
rect 3007 8820 3019 8823
rect 3510 8820 3516 8832
rect 3007 8792 3516 8820
rect 3007 8789 3019 8792
rect 2961 8783 3019 8789
rect 3510 8780 3516 8792
rect 3568 8780 3574 8832
rect 4080 8820 4108 8860
rect 7101 8891 7159 8897
rect 7101 8857 7113 8891
rect 7147 8888 7159 8891
rect 7374 8888 7380 8900
rect 7147 8860 7380 8888
rect 7147 8857 7159 8860
rect 7101 8851 7159 8857
rect 7374 8848 7380 8860
rect 7432 8848 7438 8900
rect 9677 8891 9735 8897
rect 9677 8857 9689 8891
rect 9723 8888 9735 8891
rect 9858 8888 9864 8900
rect 9723 8860 9864 8888
rect 9723 8857 9735 8860
rect 9677 8851 9735 8857
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 10502 8888 10508 8900
rect 10463 8860 10508 8888
rect 10502 8848 10508 8860
rect 10560 8848 10566 8900
rect 11333 8891 11391 8897
rect 11333 8857 11345 8891
rect 11379 8888 11391 8891
rect 11606 8888 11612 8900
rect 11379 8860 11612 8888
rect 11379 8857 11391 8860
rect 11333 8851 11391 8857
rect 11606 8848 11612 8860
rect 11664 8848 11670 8900
rect 12710 8848 12716 8900
rect 12768 8888 12774 8900
rect 12912 8888 12940 8919
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 14826 8956 14832 8968
rect 14787 8928 14832 8956
rect 14826 8916 14832 8928
rect 14884 8916 14890 8968
rect 15286 8956 15292 8968
rect 15247 8928 15292 8956
rect 15286 8916 15292 8928
rect 15344 8916 15350 8968
rect 12768 8860 12940 8888
rect 13173 8891 13231 8897
rect 12768 8848 12774 8860
rect 13173 8857 13185 8891
rect 13219 8888 13231 8891
rect 13219 8860 14320 8888
rect 13219 8857 13231 8860
rect 13173 8851 13231 8857
rect 4430 8820 4436 8832
rect 4080 8792 4436 8820
rect 4430 8780 4436 8792
rect 4488 8780 4494 8832
rect 4706 8780 4712 8832
rect 4764 8820 4770 8832
rect 5445 8823 5503 8829
rect 5445 8820 5457 8823
rect 4764 8792 5457 8820
rect 4764 8780 4770 8792
rect 5445 8789 5457 8792
rect 5491 8789 5503 8823
rect 5445 8783 5503 8789
rect 5626 8780 5632 8832
rect 5684 8820 5690 8832
rect 9398 8820 9404 8832
rect 5684 8792 9404 8820
rect 5684 8780 5690 8792
rect 9398 8780 9404 8792
rect 9456 8820 9462 8832
rect 13906 8820 13912 8832
rect 9456 8792 13912 8820
rect 9456 8780 9462 8792
rect 13906 8780 13912 8792
rect 13964 8780 13970 8832
rect 13998 8780 14004 8832
rect 14056 8820 14062 8832
rect 14185 8823 14243 8829
rect 14185 8820 14197 8823
rect 14056 8792 14197 8820
rect 14056 8780 14062 8792
rect 14185 8789 14197 8792
rect 14231 8789 14243 8823
rect 14292 8820 14320 8860
rect 14918 8848 14924 8900
rect 14976 8888 14982 8900
rect 15562 8888 15568 8900
rect 14976 8860 15568 8888
rect 14976 8848 14982 8860
rect 15562 8848 15568 8860
rect 15620 8848 15626 8900
rect 15194 8820 15200 8832
rect 14292 8792 15200 8820
rect 14185 8783 14243 8789
rect 15194 8780 15200 8792
rect 15252 8820 15258 8832
rect 16482 8820 16488 8832
rect 15252 8792 16488 8820
rect 15252 8780 15258 8792
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 1104 8730 18860 8752
rect 1104 8678 3947 8730
rect 3999 8678 4011 8730
rect 4063 8678 4075 8730
rect 4127 8678 4139 8730
rect 4191 8678 9878 8730
rect 9930 8678 9942 8730
rect 9994 8678 10006 8730
rect 10058 8678 10070 8730
rect 10122 8678 15808 8730
rect 15860 8678 15872 8730
rect 15924 8678 15936 8730
rect 15988 8678 16000 8730
rect 16052 8678 18860 8730
rect 1104 8656 18860 8678
rect 2038 8616 2044 8628
rect 1412 8588 2044 8616
rect 1412 8489 1440 8588
rect 2038 8576 2044 8588
rect 2096 8616 2102 8628
rect 2590 8616 2596 8628
rect 2096 8588 2596 8616
rect 2096 8576 2102 8588
rect 2590 8576 2596 8588
rect 2648 8576 2654 8628
rect 5902 8576 5908 8628
rect 5960 8616 5966 8628
rect 6273 8619 6331 8625
rect 6273 8616 6285 8619
rect 5960 8588 6285 8616
rect 5960 8576 5966 8588
rect 6273 8585 6285 8588
rect 6319 8585 6331 8619
rect 10505 8619 10563 8625
rect 10505 8616 10517 8619
rect 6273 8579 6331 8585
rect 7107 8588 10517 8616
rect 2406 8508 2412 8560
rect 2464 8548 2470 8560
rect 2777 8551 2835 8557
rect 2777 8548 2789 8551
rect 2464 8520 2789 8548
rect 2464 8508 2470 8520
rect 2777 8517 2789 8520
rect 2823 8517 2835 8551
rect 2777 8511 2835 8517
rect 3053 8551 3111 8557
rect 3053 8517 3065 8551
rect 3099 8517 3111 8551
rect 3053 8511 3111 8517
rect 1397 8483 1455 8489
rect 1397 8449 1409 8483
rect 1443 8449 1455 8483
rect 1397 8443 1455 8449
rect 2498 8440 2504 8492
rect 2556 8480 2562 8492
rect 3068 8480 3096 8511
rect 3326 8508 3332 8560
rect 3384 8548 3390 8560
rect 4249 8551 4307 8557
rect 4249 8548 4261 8551
rect 3384 8520 4261 8548
rect 3384 8508 3390 8520
rect 4249 8517 4261 8520
rect 4295 8517 4307 8551
rect 4249 8511 4307 8517
rect 6638 8508 6644 8560
rect 6696 8548 6702 8560
rect 7009 8551 7067 8557
rect 7009 8548 7021 8551
rect 6696 8520 7021 8548
rect 6696 8508 6702 8520
rect 7009 8517 7021 8520
rect 7055 8517 7067 8551
rect 7009 8511 7067 8517
rect 3510 8480 3516 8492
rect 2556 8452 3096 8480
rect 3471 8452 3516 8480
rect 2556 8440 2562 8452
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8480 3755 8483
rect 4706 8480 4712 8492
rect 3743 8452 4712 8480
rect 3743 8449 3755 8452
rect 3697 8443 3755 8449
rect 1664 8415 1722 8421
rect 1664 8381 1676 8415
rect 1710 8412 1722 8415
rect 3712 8412 3740 8443
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 1710 8384 3740 8412
rect 4065 8415 4123 8421
rect 1710 8381 1722 8384
rect 1664 8375 1722 8381
rect 4065 8381 4077 8415
rect 4111 8381 4123 8415
rect 4065 8375 4123 8381
rect 3694 8304 3700 8356
rect 3752 8344 3758 8356
rect 4080 8344 4108 8375
rect 4430 8372 4436 8424
rect 4488 8412 4494 8424
rect 4893 8415 4951 8421
rect 4893 8412 4905 8415
rect 4488 8384 4905 8412
rect 4488 8372 4494 8384
rect 4893 8381 4905 8384
rect 4939 8381 4951 8415
rect 7107 8412 7135 8588
rect 10505 8585 10517 8588
rect 10551 8616 10563 8619
rect 10870 8616 10876 8628
rect 10551 8588 10876 8616
rect 10551 8585 10563 8588
rect 10505 8579 10563 8585
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 16114 8616 16120 8628
rect 12492 8588 12537 8616
rect 13464 8588 15792 8616
rect 12492 8576 12498 8588
rect 9214 8508 9220 8560
rect 9272 8548 9278 8560
rect 9582 8548 9588 8560
rect 9272 8520 9588 8548
rect 9272 8508 9278 8520
rect 9582 8508 9588 8520
rect 9640 8548 9646 8560
rect 10318 8548 10324 8560
rect 9640 8520 10324 8548
rect 9640 8508 9646 8520
rect 10318 8508 10324 8520
rect 10376 8508 10382 8560
rect 11149 8551 11207 8557
rect 11149 8517 11161 8551
rect 11195 8548 11207 8551
rect 13262 8548 13268 8560
rect 11195 8520 13268 8548
rect 11195 8517 11207 8520
rect 11149 8511 11207 8517
rect 13262 8508 13268 8520
rect 13320 8508 13326 8560
rect 11698 8480 11704 8492
rect 11659 8452 11704 8480
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 12710 8440 12716 8492
rect 12768 8480 12774 8492
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12768 8452 13001 8480
rect 12768 8440 12774 8452
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 13464 8480 13492 8588
rect 13541 8551 13599 8557
rect 13541 8517 13553 8551
rect 13587 8548 13599 8551
rect 15562 8548 15568 8560
rect 13587 8520 14504 8548
rect 13587 8517 13599 8520
rect 13541 8511 13599 8517
rect 13998 8480 14004 8492
rect 13464 8452 13584 8480
rect 13959 8452 14004 8480
rect 12989 8443 13047 8449
rect 7169 8415 7227 8421
rect 7169 8412 7181 8415
rect 7107 8384 7181 8412
rect 4893 8375 4951 8381
rect 7169 8381 7181 8384
rect 7215 8381 7227 8415
rect 7169 8375 7227 8381
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8412 7619 8415
rect 7650 8412 7656 8424
rect 7607 8384 7656 8412
rect 7607 8381 7619 8384
rect 7561 8375 7619 8381
rect 7650 8372 7656 8384
rect 7708 8372 7714 8424
rect 7828 8415 7886 8421
rect 7828 8381 7840 8415
rect 7874 8412 7886 8415
rect 11054 8412 11060 8424
rect 7874 8384 11060 8412
rect 7874 8381 7886 8384
rect 7828 8375 7886 8381
rect 11054 8372 11060 8384
rect 11112 8372 11118 8424
rect 11517 8415 11575 8421
rect 11517 8381 11529 8415
rect 11563 8412 11575 8415
rect 13446 8412 13452 8424
rect 11563 8384 13452 8412
rect 11563 8381 11575 8384
rect 11517 8375 11575 8381
rect 13446 8372 13452 8384
rect 13504 8372 13510 8424
rect 5166 8353 5172 8356
rect 5160 8344 5172 8353
rect 3752 8316 4108 8344
rect 5127 8316 5172 8344
rect 3752 8304 3758 8316
rect 5160 8307 5172 8316
rect 5166 8304 5172 8307
rect 5224 8304 5230 8356
rect 8110 8304 8116 8356
rect 8168 8344 8174 8356
rect 9217 8347 9275 8353
rect 9217 8344 9229 8347
rect 8168 8316 9229 8344
rect 8168 8304 8174 8316
rect 9217 8313 9229 8316
rect 9263 8313 9275 8347
rect 9217 8307 9275 8313
rect 9490 8304 9496 8356
rect 9548 8344 9554 8356
rect 11606 8344 11612 8356
rect 9548 8316 11468 8344
rect 11567 8316 11612 8344
rect 9548 8304 9554 8316
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 3421 8279 3479 8285
rect 3421 8276 3433 8279
rect 3016 8248 3433 8276
rect 3016 8236 3022 8248
rect 3421 8245 3433 8248
rect 3467 8276 3479 8279
rect 3510 8276 3516 8288
rect 3467 8248 3516 8276
rect 3467 8245 3479 8248
rect 3421 8239 3479 8245
rect 3510 8236 3516 8248
rect 3568 8236 3574 8288
rect 6730 8236 6736 8288
rect 6788 8276 6794 8288
rect 7558 8276 7564 8288
rect 6788 8248 7564 8276
rect 6788 8236 6794 8248
rect 7558 8236 7564 8248
rect 7616 8236 7622 8288
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 8941 8279 8999 8285
rect 8941 8276 8953 8279
rect 8812 8248 8953 8276
rect 8812 8236 8818 8248
rect 8941 8245 8953 8248
rect 8987 8245 8999 8279
rect 11440 8276 11468 8316
rect 11606 8304 11612 8316
rect 11664 8304 11670 8356
rect 12897 8347 12955 8353
rect 12897 8344 12909 8347
rect 11716 8316 12909 8344
rect 11716 8276 11744 8316
rect 12897 8313 12909 8316
rect 12943 8344 12955 8347
rect 13556 8344 13584 8452
rect 13998 8440 14004 8452
rect 14056 8440 14062 8492
rect 14185 8483 14243 8489
rect 14185 8449 14197 8483
rect 14231 8449 14243 8483
rect 14476 8480 14504 8520
rect 14752 8520 15568 8548
rect 14752 8480 14780 8520
rect 15562 8508 15568 8520
rect 15620 8508 15626 8560
rect 14476 8452 14780 8480
rect 14185 8443 14243 8449
rect 14200 8412 14228 8443
rect 14826 8440 14832 8492
rect 14884 8480 14890 8492
rect 15105 8483 15163 8489
rect 15105 8480 15117 8483
rect 14884 8452 15117 8480
rect 14884 8440 14890 8452
rect 15105 8449 15117 8452
rect 15151 8449 15163 8483
rect 15105 8443 15163 8449
rect 15764 8412 15792 8588
rect 15856 8588 16120 8616
rect 15856 8489 15884 8588
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 16206 8576 16212 8628
rect 16264 8616 16270 8628
rect 17126 8616 17132 8628
rect 16264 8588 17132 8616
rect 16264 8576 16270 8588
rect 17126 8576 17132 8588
rect 17184 8616 17190 8628
rect 17221 8619 17279 8625
rect 17221 8616 17233 8619
rect 17184 8588 17233 8616
rect 17184 8576 17190 8588
rect 17221 8585 17233 8588
rect 17267 8585 17279 8619
rect 17221 8579 17279 8585
rect 17862 8508 17868 8560
rect 17920 8548 17926 8560
rect 18233 8551 18291 8557
rect 18233 8548 18245 8551
rect 17920 8520 18245 8548
rect 17920 8508 17926 8520
rect 18233 8517 18245 8520
rect 18279 8517 18291 8551
rect 18233 8511 18291 8517
rect 15841 8483 15899 8489
rect 15841 8449 15853 8483
rect 15887 8449 15899 8483
rect 15841 8443 15899 8449
rect 17126 8412 17132 8424
rect 14200 8384 15700 8412
rect 15764 8384 17132 8412
rect 12943 8316 13584 8344
rect 13909 8347 13967 8353
rect 12943 8313 12955 8316
rect 12897 8307 12955 8313
rect 13909 8313 13921 8347
rect 13955 8344 13967 8347
rect 15013 8347 15071 8353
rect 13955 8316 14596 8344
rect 13955 8313 13967 8316
rect 13909 8307 13967 8313
rect 11440 8248 11744 8276
rect 8941 8239 8999 8245
rect 12250 8236 12256 8288
rect 12308 8276 12314 8288
rect 12805 8279 12863 8285
rect 12805 8276 12817 8279
rect 12308 8248 12817 8276
rect 12308 8236 12314 8248
rect 12805 8245 12817 8248
rect 12851 8276 12863 8279
rect 13538 8276 13544 8288
rect 12851 8248 13544 8276
rect 12851 8245 12863 8248
rect 12805 8239 12863 8245
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 14568 8285 14596 8316
rect 15013 8313 15025 8347
rect 15059 8344 15071 8347
rect 15102 8344 15108 8356
rect 15059 8316 15108 8344
rect 15059 8313 15071 8316
rect 15013 8307 15071 8313
rect 15102 8304 15108 8316
rect 15160 8304 15166 8356
rect 15672 8344 15700 8384
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 18046 8412 18052 8424
rect 18007 8384 18052 8412
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 16086 8347 16144 8353
rect 16086 8344 16098 8347
rect 15672 8316 16098 8344
rect 16086 8313 16098 8316
rect 16132 8344 16144 8347
rect 16482 8344 16488 8356
rect 16132 8316 16488 8344
rect 16132 8313 16144 8316
rect 16086 8307 16144 8313
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 14553 8279 14611 8285
rect 14553 8245 14565 8279
rect 14599 8245 14611 8279
rect 14918 8276 14924 8288
rect 14879 8248 14924 8276
rect 14553 8239 14611 8245
rect 14918 8236 14924 8248
rect 14976 8236 14982 8288
rect 1104 8186 18860 8208
rect 1104 8134 6912 8186
rect 6964 8134 6976 8186
rect 7028 8134 7040 8186
rect 7092 8134 7104 8186
rect 7156 8134 12843 8186
rect 12895 8134 12907 8186
rect 12959 8134 12971 8186
rect 13023 8134 13035 8186
rect 13087 8134 18860 8186
rect 1104 8112 18860 8134
rect 2317 8075 2375 8081
rect 2317 8041 2329 8075
rect 2363 8072 2375 8075
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 2363 8044 4077 8072
rect 2363 8041 2375 8044
rect 2317 8035 2375 8041
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 4065 8035 4123 8041
rect 4433 8075 4491 8081
rect 4433 8041 4445 8075
rect 4479 8072 4491 8075
rect 4614 8072 4620 8084
rect 4479 8044 4620 8072
rect 4479 8041 4491 8044
rect 4433 8035 4491 8041
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 5077 8075 5135 8081
rect 5077 8041 5089 8075
rect 5123 8072 5135 8075
rect 5350 8072 5356 8084
rect 5123 8044 5356 8072
rect 5123 8041 5135 8044
rect 5077 8035 5135 8041
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 6089 8075 6147 8081
rect 6089 8041 6101 8075
rect 6135 8041 6147 8075
rect 6089 8035 6147 8041
rect 6457 8075 6515 8081
rect 6457 8041 6469 8075
rect 6503 8072 6515 8075
rect 7653 8075 7711 8081
rect 7653 8072 7665 8075
rect 6503 8044 7665 8072
rect 6503 8041 6515 8044
rect 6457 8035 6515 8041
rect 7653 8041 7665 8044
rect 7699 8041 7711 8075
rect 7653 8035 7711 8041
rect 2958 7964 2964 8016
rect 3016 8004 3022 8016
rect 3237 8007 3295 8013
rect 3237 8004 3249 8007
rect 3016 7976 3249 8004
rect 3016 7964 3022 7976
rect 3237 7973 3249 7976
rect 3283 7973 3295 8007
rect 3237 7967 3295 7973
rect 3602 7964 3608 8016
rect 3660 8004 3666 8016
rect 5445 8007 5503 8013
rect 5445 8004 5457 8007
rect 3660 7976 5457 8004
rect 3660 7964 3666 7976
rect 5445 7973 5457 7976
rect 5491 7973 5503 8007
rect 6104 8004 6132 8035
rect 8570 8032 8576 8084
rect 8628 8072 8634 8084
rect 8665 8075 8723 8081
rect 8665 8072 8677 8075
rect 8628 8044 8677 8072
rect 8628 8032 8634 8044
rect 8665 8041 8677 8044
rect 8711 8041 8723 8075
rect 8665 8035 8723 8041
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 12710 8072 12716 8084
rect 8904 8044 11836 8072
rect 12671 8044 12716 8072
rect 8904 8032 8910 8044
rect 7374 8004 7380 8016
rect 6104 7976 7380 8004
rect 5445 7967 5503 7973
rect 7374 7964 7380 7976
rect 7432 7964 7438 8016
rect 8021 8007 8079 8013
rect 8021 7973 8033 8007
rect 8067 8004 8079 8007
rect 9674 8004 9680 8016
rect 8067 7976 9680 8004
rect 8067 7973 8079 7976
rect 8021 7967 8079 7973
rect 9674 7964 9680 7976
rect 9732 7964 9738 8016
rect 10042 7964 10048 8016
rect 10100 8004 10106 8016
rect 10100 7976 10145 8004
rect 10100 7964 10106 7976
rect 10410 7964 10416 8016
rect 10468 8004 10474 8016
rect 10686 8004 10692 8016
rect 10468 7976 10692 8004
rect 10468 7964 10474 7976
rect 10686 7964 10692 7976
rect 10744 7964 10750 8016
rect 11600 8007 11658 8013
rect 11600 7973 11612 8007
rect 11646 8004 11658 8007
rect 11698 8004 11704 8016
rect 11646 7976 11704 8004
rect 11646 7973 11658 7976
rect 11600 7967 11658 7973
rect 11698 7964 11704 7976
rect 11756 7964 11762 8016
rect 2222 7936 2228 7948
rect 2183 7908 2228 7936
rect 2222 7896 2228 7908
rect 2280 7896 2286 7948
rect 3329 7939 3387 7945
rect 3329 7905 3341 7939
rect 3375 7936 3387 7939
rect 6086 7936 6092 7948
rect 3375 7908 6092 7936
rect 3375 7905 3387 7908
rect 3329 7899 3387 7905
rect 2406 7868 2412 7880
rect 2367 7840 2412 7868
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2314 7760 2320 7812
rect 2372 7800 2378 7812
rect 2869 7803 2927 7809
rect 2869 7800 2881 7803
rect 2372 7772 2881 7800
rect 2372 7760 2378 7772
rect 2869 7769 2881 7772
rect 2915 7769 2927 7803
rect 2869 7763 2927 7769
rect 3234 7760 3240 7812
rect 3292 7800 3298 7812
rect 3344 7800 3372 7899
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 7101 7939 7159 7945
rect 7101 7905 7113 7939
rect 7147 7905 7159 7939
rect 7101 7899 7159 7905
rect 8113 7939 8171 7945
rect 8113 7905 8125 7939
rect 8159 7936 8171 7939
rect 9766 7936 9772 7948
rect 8159 7908 9772 7936
rect 8159 7905 8171 7908
rect 8113 7899 8171 7905
rect 3513 7871 3571 7877
rect 3513 7837 3525 7871
rect 3559 7868 3571 7871
rect 4522 7868 4528 7880
rect 3559 7840 3832 7868
rect 4483 7840 4528 7868
rect 3559 7837 3571 7840
rect 3513 7831 3571 7837
rect 3292 7772 3372 7800
rect 3804 7800 3832 7840
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 4706 7868 4712 7880
rect 4667 7840 4712 7868
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7837 5595 7871
rect 5718 7868 5724 7880
rect 5679 7840 5724 7868
rect 5537 7831 5595 7837
rect 4724 7800 4752 7828
rect 3804 7772 4752 7800
rect 5552 7800 5580 7831
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 6546 7868 6552 7880
rect 6507 7840 6552 7868
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 6730 7868 6736 7880
rect 6691 7840 6736 7868
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 7116 7868 7144 7899
rect 9766 7896 9772 7908
rect 9824 7896 9830 7948
rect 9858 7896 9864 7948
rect 9916 7936 9922 7948
rect 10134 7936 10140 7948
rect 9916 7908 10140 7936
rect 9916 7896 9922 7908
rect 10134 7896 10140 7908
rect 10192 7896 10198 7948
rect 10318 7896 10324 7948
rect 10376 7936 10382 7948
rect 11333 7939 11391 7945
rect 11333 7936 11345 7939
rect 10376 7908 11345 7936
rect 10376 7896 10382 7908
rect 11333 7905 11345 7908
rect 11379 7905 11391 7939
rect 11808 7936 11836 8044
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 13354 8072 13360 8084
rect 13315 8044 13360 8072
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 14366 8032 14372 8084
rect 14424 8072 14430 8084
rect 14645 8075 14703 8081
rect 14645 8072 14657 8075
rect 14424 8044 14657 8072
rect 14424 8032 14430 8044
rect 14645 8041 14657 8044
rect 14691 8041 14703 8075
rect 14645 8035 14703 8041
rect 16482 8032 16488 8084
rect 16540 8072 16546 8084
rect 16669 8075 16727 8081
rect 16669 8072 16681 8075
rect 16540 8044 16681 8072
rect 16540 8032 16546 8044
rect 16669 8041 16681 8044
rect 16715 8041 16727 8075
rect 16669 8035 16727 8041
rect 16850 8032 16856 8084
rect 16908 8072 16914 8084
rect 16945 8075 17003 8081
rect 16945 8072 16957 8075
rect 16908 8044 16957 8072
rect 16908 8032 16914 8044
rect 16945 8041 16957 8044
rect 16991 8041 17003 8075
rect 17310 8072 17316 8084
rect 17271 8044 17316 8072
rect 16945 8035 17003 8041
rect 17310 8032 17316 8044
rect 17368 8032 17374 8084
rect 13906 7964 13912 8016
rect 13964 8004 13970 8016
rect 14553 8007 14611 8013
rect 14553 8004 14565 8007
rect 13964 7976 14565 8004
rect 13964 7964 13970 7976
rect 14553 7973 14565 7976
rect 14599 8004 14611 8007
rect 14599 7976 18000 8004
rect 14599 7973 14611 7976
rect 14553 7967 14611 7973
rect 13354 7936 13360 7948
rect 11808 7908 13360 7936
rect 11333 7899 11391 7905
rect 13354 7896 13360 7908
rect 13412 7896 13418 7948
rect 13630 7936 13636 7948
rect 13464 7908 13636 7936
rect 8202 7868 8208 7880
rect 7116 7840 8064 7868
rect 8163 7840 8208 7868
rect 7098 7800 7104 7812
rect 5552 7772 7104 7800
rect 3292 7760 3298 7772
rect 7098 7760 7104 7772
rect 7156 7760 7162 7812
rect 8036 7800 8064 7840
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 8938 7828 8944 7880
rect 8996 7868 9002 7880
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 8996 7840 10241 7868
rect 8996 7828 9002 7840
rect 10229 7837 10241 7840
rect 10275 7837 10287 7871
rect 10686 7868 10692 7880
rect 10647 7840 10692 7868
rect 10229 7831 10287 7837
rect 10686 7828 10692 7840
rect 10744 7828 10750 7880
rect 13464 7877 13492 7908
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 17972 7945 18000 7976
rect 15545 7939 15603 7945
rect 15545 7936 15557 7939
rect 14844 7908 15557 7936
rect 14844 7880 14872 7908
rect 15545 7905 15557 7908
rect 15591 7905 15603 7939
rect 15545 7899 15603 7905
rect 17957 7939 18015 7945
rect 17957 7905 17969 7939
rect 18003 7905 18015 7939
rect 17957 7899 18015 7905
rect 13449 7871 13507 7877
rect 13449 7868 13461 7871
rect 12360 7840 13461 7868
rect 8036 7772 11376 7800
rect 1854 7732 1860 7744
rect 1815 7704 1860 7732
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 3786 7692 3792 7744
rect 3844 7732 3850 7744
rect 7285 7735 7343 7741
rect 7285 7732 7297 7735
rect 3844 7704 7297 7732
rect 3844 7692 3850 7704
rect 7285 7701 7297 7704
rect 7331 7701 7343 7735
rect 7285 7695 7343 7701
rect 8018 7692 8024 7744
rect 8076 7732 8082 7744
rect 8202 7732 8208 7744
rect 8076 7704 8208 7732
rect 8076 7692 8082 7704
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8294 7692 8300 7744
rect 8352 7732 8358 7744
rect 9677 7735 9735 7741
rect 9677 7732 9689 7735
rect 8352 7704 9689 7732
rect 8352 7692 8358 7704
rect 9677 7701 9689 7704
rect 9723 7701 9735 7735
rect 11348 7732 11376 7772
rect 12360 7732 12388 7840
rect 13449 7837 13461 7840
rect 13495 7837 13507 7871
rect 13449 7831 13507 7837
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7837 13599 7871
rect 14826 7868 14832 7880
rect 14787 7840 14832 7868
rect 13541 7831 13599 7837
rect 13170 7760 13176 7812
rect 13228 7800 13234 7812
rect 13556 7800 13584 7831
rect 14826 7828 14832 7840
rect 14884 7828 14890 7880
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 13228 7772 13584 7800
rect 13228 7760 13234 7772
rect 13630 7760 13636 7812
rect 13688 7800 13694 7812
rect 15304 7800 15332 7831
rect 17126 7828 17132 7880
rect 17184 7868 17190 7880
rect 17405 7871 17463 7877
rect 17405 7868 17417 7871
rect 17184 7840 17417 7868
rect 17184 7828 17190 7840
rect 17405 7837 17417 7840
rect 17451 7837 17463 7871
rect 17405 7831 17463 7837
rect 17494 7828 17500 7880
rect 17552 7868 17558 7880
rect 17552 7840 17597 7868
rect 17552 7828 17558 7840
rect 18138 7800 18144 7812
rect 13688 7772 15332 7800
rect 18099 7772 18144 7800
rect 13688 7760 13694 7772
rect 18138 7760 18144 7772
rect 18196 7760 18202 7812
rect 11348 7704 12388 7732
rect 12989 7735 13047 7741
rect 9677 7695 9735 7701
rect 12989 7701 13001 7735
rect 13035 7732 13047 7735
rect 13814 7732 13820 7744
rect 13035 7704 13820 7732
rect 13035 7701 13047 7704
rect 12989 7695 13047 7701
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 14185 7735 14243 7741
rect 14185 7701 14197 7735
rect 14231 7732 14243 7735
rect 15654 7732 15660 7744
rect 14231 7704 15660 7732
rect 14231 7701 14243 7704
rect 14185 7695 14243 7701
rect 15654 7692 15660 7704
rect 15712 7692 15718 7744
rect 1104 7642 18860 7664
rect 1104 7590 3947 7642
rect 3999 7590 4011 7642
rect 4063 7590 4075 7642
rect 4127 7590 4139 7642
rect 4191 7590 9878 7642
rect 9930 7590 9942 7642
rect 9994 7590 10006 7642
rect 10058 7590 10070 7642
rect 10122 7590 15808 7642
rect 15860 7590 15872 7642
rect 15924 7590 15936 7642
rect 15988 7590 16000 7642
rect 16052 7590 18860 7642
rect 1104 7568 18860 7590
rect 2222 7488 2228 7540
rect 2280 7528 2286 7540
rect 3697 7531 3755 7537
rect 3697 7528 3709 7531
rect 2280 7500 3709 7528
rect 2280 7488 2286 7500
rect 3697 7497 3709 7500
rect 3743 7497 3755 7531
rect 3697 7491 3755 7497
rect 5166 7488 5172 7540
rect 5224 7528 5230 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 5224 7500 6377 7528
rect 5224 7488 5230 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 7098 7528 7104 7540
rect 7059 7500 7104 7528
rect 6365 7491 6423 7497
rect 7098 7488 7104 7500
rect 7156 7488 7162 7540
rect 11698 7528 11704 7540
rect 7208 7500 11284 7528
rect 11659 7500 11704 7528
rect 6178 7420 6184 7472
rect 6236 7460 6242 7472
rect 7208 7460 7236 7500
rect 6236 7432 7236 7460
rect 11256 7460 11284 7500
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 11977 7531 12035 7537
rect 11977 7497 11989 7531
rect 12023 7528 12035 7531
rect 12158 7528 12164 7540
rect 12023 7500 12164 7528
rect 12023 7497 12035 7500
rect 11977 7491 12035 7497
rect 12158 7488 12164 7500
rect 12216 7488 12222 7540
rect 12342 7488 12348 7540
rect 12400 7528 12406 7540
rect 16390 7528 16396 7540
rect 12400 7500 16396 7528
rect 12400 7488 12406 7500
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 16577 7531 16635 7537
rect 16577 7497 16589 7531
rect 16623 7528 16635 7531
rect 16758 7528 16764 7540
rect 16623 7500 16764 7528
rect 16623 7497 16635 7500
rect 16577 7491 16635 7497
rect 16758 7488 16764 7500
rect 16816 7488 16822 7540
rect 12360 7460 12388 7488
rect 13446 7460 13452 7472
rect 11256 7432 12388 7460
rect 13407 7432 13452 7460
rect 6236 7420 6242 7432
rect 13446 7420 13452 7432
rect 13504 7420 13510 7472
rect 18230 7460 18236 7472
rect 13556 7432 14044 7460
rect 18191 7432 18236 7460
rect 2682 7352 2688 7404
rect 2740 7392 2746 7404
rect 3142 7392 3148 7404
rect 2740 7364 3148 7392
rect 2740 7352 2746 7364
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 4706 7392 4712 7404
rect 4387 7364 4712 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 4798 7352 4804 7404
rect 4856 7392 4862 7404
rect 4985 7395 5043 7401
rect 4985 7392 4997 7395
rect 4856 7364 4997 7392
rect 4856 7352 4862 7364
rect 4985 7361 4997 7364
rect 5031 7361 5043 7395
rect 7650 7392 7656 7404
rect 7611 7364 7656 7392
rect 4985 7355 5043 7361
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 10318 7392 10324 7404
rect 10279 7364 10324 7392
rect 10318 7352 10324 7364
rect 10376 7352 10382 7404
rect 11330 7352 11336 7404
rect 11388 7392 11394 7404
rect 11790 7392 11796 7404
rect 11388 7364 11796 7392
rect 11388 7352 11394 7364
rect 11790 7352 11796 7364
rect 11848 7392 11854 7404
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 11848 7364 12909 7392
rect 11848 7352 11854 7364
rect 12897 7361 12909 7364
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 13170 7392 13176 7404
rect 13127 7364 13176 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 1581 7327 1639 7333
rect 1581 7293 1593 7327
rect 1627 7293 1639 7327
rect 1581 7287 1639 7293
rect 1848 7327 1906 7333
rect 1848 7293 1860 7327
rect 1894 7324 1906 7327
rect 2406 7324 2412 7336
rect 1894 7296 2412 7324
rect 1894 7293 1906 7296
rect 1848 7287 1906 7293
rect 1596 7256 1624 7287
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 3694 7284 3700 7336
rect 3752 7324 3758 7336
rect 4893 7327 4951 7333
rect 3752 7296 4200 7324
rect 3752 7284 3758 7296
rect 2314 7256 2320 7268
rect 1596 7228 2320 7256
rect 2314 7216 2320 7228
rect 2372 7216 2378 7268
rect 4172 7265 4200 7296
rect 4893 7293 4905 7327
rect 4939 7293 4951 7327
rect 6638 7324 6644 7336
rect 4893 7287 4951 7293
rect 5184 7296 6644 7324
rect 3237 7259 3295 7265
rect 3237 7225 3249 7259
rect 3283 7256 3295 7259
rect 4065 7259 4123 7265
rect 4065 7256 4077 7259
rect 3283 7228 4077 7256
rect 3283 7225 3295 7228
rect 3237 7219 3295 7225
rect 4065 7225 4077 7228
rect 4111 7225 4123 7259
rect 4065 7219 4123 7225
rect 4157 7259 4215 7265
rect 4157 7225 4169 7259
rect 4203 7256 4215 7259
rect 4908 7256 4936 7287
rect 5184 7256 5212 7296
rect 6638 7284 6644 7296
rect 6696 7284 6702 7336
rect 7190 7284 7196 7336
rect 7248 7324 7254 7336
rect 7469 7327 7527 7333
rect 7469 7324 7481 7327
rect 7248 7296 7481 7324
rect 7248 7284 7254 7296
rect 7469 7293 7481 7296
rect 7515 7293 7527 7327
rect 7469 7287 7527 7293
rect 7561 7327 7619 7333
rect 7561 7293 7573 7327
rect 7607 7324 7619 7327
rect 7742 7324 7748 7336
rect 7607 7296 7748 7324
rect 7607 7293 7619 7296
rect 7561 7287 7619 7293
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 8478 7324 8484 7336
rect 8439 7296 8484 7324
rect 8478 7284 8484 7296
rect 8536 7284 8542 7336
rect 8754 7333 8760 7336
rect 8748 7324 8760 7333
rect 8715 7296 8760 7324
rect 8748 7287 8760 7296
rect 8812 7324 8818 7336
rect 10226 7324 10232 7336
rect 8812 7296 10232 7324
rect 8754 7284 8760 7287
rect 8812 7284 8818 7296
rect 10226 7284 10232 7296
rect 10284 7284 10290 7336
rect 10870 7284 10876 7336
rect 10928 7324 10934 7336
rect 12161 7327 12219 7333
rect 12161 7324 12173 7327
rect 10928 7296 12173 7324
rect 10928 7284 10934 7296
rect 12161 7293 12173 7296
rect 12207 7293 12219 7327
rect 12161 7287 12219 7293
rect 12250 7284 12256 7336
rect 12308 7324 12314 7336
rect 13556 7324 13584 7432
rect 14016 7401 14044 7432
rect 18230 7420 18236 7432
rect 18288 7420 18294 7472
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 12308 7296 13584 7324
rect 13648 7364 13921 7392
rect 12308 7284 12314 7296
rect 4203 7228 4844 7256
rect 4908 7228 5212 7256
rect 5252 7259 5310 7265
rect 4203 7225 4215 7228
rect 4157 7219 4215 7225
rect 2958 7188 2964 7200
rect 2919 7160 2964 7188
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 4706 7188 4712 7200
rect 4667 7160 4712 7188
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 4816 7188 4844 7228
rect 5252 7225 5264 7259
rect 5298 7256 5310 7259
rect 5718 7256 5724 7268
rect 5298 7228 5724 7256
rect 5298 7225 5310 7228
rect 5252 7219 5310 7225
rect 5718 7216 5724 7228
rect 5776 7256 5782 7268
rect 8938 7256 8944 7268
rect 5776 7228 8944 7256
rect 5776 7216 5782 7228
rect 8938 7216 8944 7228
rect 8996 7216 9002 7268
rect 9674 7216 9680 7268
rect 9732 7256 9738 7268
rect 10588 7259 10646 7265
rect 9732 7228 10548 7256
rect 9732 7216 9738 7228
rect 10520 7200 10548 7228
rect 10588 7225 10600 7259
rect 10634 7256 10646 7259
rect 12268 7256 12296 7284
rect 13648 7256 13676 7364
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 14001 7395 14059 7401
rect 14001 7361 14013 7395
rect 14047 7361 14059 7395
rect 14001 7355 14059 7361
rect 14826 7352 14832 7404
rect 14884 7392 14890 7404
rect 15105 7395 15163 7401
rect 15105 7392 15117 7395
rect 14884 7364 15117 7392
rect 14884 7352 14890 7364
rect 15105 7361 15117 7364
rect 15151 7361 15163 7395
rect 15105 7355 15163 7361
rect 15654 7352 15660 7404
rect 15712 7392 15718 7404
rect 16025 7395 16083 7401
rect 16025 7392 16037 7395
rect 15712 7364 16037 7392
rect 15712 7352 15718 7364
rect 16025 7361 16037 7364
rect 16071 7361 16083 7395
rect 16025 7355 16083 7361
rect 16209 7395 16267 7401
rect 16209 7361 16221 7395
rect 16255 7392 16267 7395
rect 16482 7392 16488 7404
rect 16255 7364 16488 7392
rect 16255 7361 16267 7364
rect 16209 7355 16267 7361
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 16666 7352 16672 7404
rect 16724 7392 16730 7404
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 16724 7364 17049 7392
rect 16724 7352 16730 7364
rect 17037 7361 17049 7364
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 17221 7395 17279 7401
rect 17221 7361 17233 7395
rect 17267 7392 17279 7395
rect 17586 7392 17592 7404
rect 17267 7364 17592 7392
rect 17267 7361 17279 7364
rect 17221 7355 17279 7361
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 14921 7327 14979 7333
rect 14921 7293 14933 7327
rect 14967 7324 14979 7327
rect 15286 7324 15292 7336
rect 14967 7296 15292 7324
rect 14967 7293 14979 7296
rect 14921 7287 14979 7293
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 16942 7324 16948 7336
rect 16903 7296 16948 7324
rect 16942 7284 16948 7296
rect 17000 7284 17006 7336
rect 17954 7284 17960 7336
rect 18012 7324 18018 7336
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 18012 7296 18061 7324
rect 18012 7284 18018 7296
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 13814 7256 13820 7268
rect 10634 7228 12296 7256
rect 12452 7228 13676 7256
rect 13775 7228 13820 7256
rect 10634 7225 10646 7228
rect 10588 7219 10646 7225
rect 6178 7188 6184 7200
rect 4816 7160 6184 7188
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 7558 7148 7564 7200
rect 7616 7188 7622 7200
rect 7742 7188 7748 7200
rect 7616 7160 7748 7188
rect 7616 7148 7622 7160
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 9398 7148 9404 7200
rect 9456 7188 9462 7200
rect 9861 7191 9919 7197
rect 9861 7188 9873 7191
rect 9456 7160 9873 7188
rect 9456 7148 9462 7160
rect 9861 7157 9873 7160
rect 9907 7157 9919 7191
rect 9861 7151 9919 7157
rect 10502 7148 10508 7200
rect 10560 7148 10566 7200
rect 12452 7197 12480 7228
rect 13814 7216 13820 7228
rect 13872 7216 13878 7268
rect 15933 7259 15991 7265
rect 15933 7256 15945 7259
rect 14568 7228 15945 7256
rect 12437 7191 12495 7197
rect 12437 7157 12449 7191
rect 12483 7157 12495 7191
rect 12437 7151 12495 7157
rect 12805 7191 12863 7197
rect 12805 7157 12817 7191
rect 12851 7188 12863 7191
rect 14090 7188 14096 7200
rect 12851 7160 14096 7188
rect 12851 7157 12863 7160
rect 12805 7151 12863 7157
rect 14090 7148 14096 7160
rect 14148 7148 14154 7200
rect 14568 7197 14596 7228
rect 15933 7225 15945 7228
rect 15979 7225 15991 7259
rect 15933 7219 15991 7225
rect 14553 7191 14611 7197
rect 14553 7157 14565 7191
rect 14599 7157 14611 7191
rect 14553 7151 14611 7157
rect 14642 7148 14648 7200
rect 14700 7188 14706 7200
rect 15013 7191 15071 7197
rect 15013 7188 15025 7191
rect 14700 7160 15025 7188
rect 14700 7148 14706 7160
rect 15013 7157 15025 7160
rect 15059 7157 15071 7191
rect 15013 7151 15071 7157
rect 15565 7191 15623 7197
rect 15565 7157 15577 7191
rect 15611 7188 15623 7191
rect 15654 7188 15660 7200
rect 15611 7160 15660 7188
rect 15611 7157 15623 7160
rect 15565 7151 15623 7157
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 1104 7098 18860 7120
rect 1104 7046 6912 7098
rect 6964 7046 6976 7098
rect 7028 7046 7040 7098
rect 7092 7046 7104 7098
rect 7156 7046 12843 7098
rect 12895 7046 12907 7098
rect 12959 7046 12971 7098
rect 13023 7046 13035 7098
rect 13087 7046 18860 7098
rect 1104 7024 18860 7046
rect 2314 6944 2320 6996
rect 2372 6984 2378 6996
rect 3881 6987 3939 6993
rect 3881 6984 3893 6987
rect 2372 6956 3893 6984
rect 2372 6944 2378 6956
rect 3881 6953 3893 6956
rect 3927 6984 3939 6987
rect 4798 6984 4804 6996
rect 3927 6956 4804 6984
rect 3927 6953 3939 6956
rect 3881 6947 3939 6953
rect 4798 6944 4804 6956
rect 4856 6944 4862 6996
rect 6365 6987 6423 6993
rect 6365 6953 6377 6987
rect 6411 6984 6423 6987
rect 6546 6984 6552 6996
rect 6411 6956 6552 6984
rect 6411 6953 6423 6956
rect 6365 6947 6423 6953
rect 6546 6944 6552 6956
rect 6604 6944 6610 6996
rect 7193 6987 7251 6993
rect 7193 6953 7205 6987
rect 7239 6984 7251 6987
rect 8018 6984 8024 6996
rect 7239 6956 8024 6984
rect 7239 6953 7251 6956
rect 7193 6947 7251 6953
rect 8018 6944 8024 6956
rect 8076 6944 8082 6996
rect 8757 6987 8815 6993
rect 8757 6953 8769 6987
rect 8803 6984 8815 6987
rect 8938 6984 8944 6996
rect 8803 6956 8944 6984
rect 8803 6953 8815 6956
rect 8757 6947 8815 6953
rect 8938 6944 8944 6956
rect 8996 6944 9002 6996
rect 9582 6944 9588 6996
rect 9640 6984 9646 6996
rect 10134 6984 10140 6996
rect 9640 6956 10140 6984
rect 9640 6944 9646 6956
rect 10134 6944 10140 6956
rect 10192 6944 10198 6996
rect 13170 6944 13176 6996
rect 13228 6984 13234 6996
rect 13357 6987 13415 6993
rect 13357 6984 13369 6987
rect 13228 6956 13369 6984
rect 13228 6944 13234 6956
rect 13357 6953 13369 6956
rect 13403 6984 13415 6987
rect 14921 6987 14979 6993
rect 14921 6984 14933 6987
rect 13403 6956 14933 6984
rect 13403 6953 13415 6956
rect 13357 6947 13415 6953
rect 14921 6953 14933 6956
rect 14967 6953 14979 6987
rect 15654 6984 15660 6996
rect 15615 6956 15660 6984
rect 14921 6947 14979 6953
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 3970 6916 3976 6928
rect 1688 6888 3976 6916
rect 1688 6857 1716 6888
rect 3970 6876 3976 6888
rect 4028 6876 4034 6928
rect 4614 6876 4620 6928
rect 4672 6916 4678 6928
rect 6733 6919 6791 6925
rect 4672 6888 5580 6916
rect 4672 6876 4678 6888
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6817 1731 6851
rect 2314 6848 2320 6860
rect 2275 6820 2320 6848
rect 1673 6811 1731 6817
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 2584 6851 2642 6857
rect 2584 6817 2596 6851
rect 2630 6848 2642 6851
rect 2958 6848 2964 6860
rect 2630 6820 2964 6848
rect 2630 6817 2642 6820
rect 2584 6811 2642 6817
rect 2958 6808 2964 6820
rect 3016 6808 3022 6860
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 4072 6851 4130 6857
rect 4072 6848 4084 6851
rect 3927 6820 4084 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 4072 6817 4084 6820
rect 4118 6817 4130 6851
rect 4332 6851 4390 6857
rect 4332 6848 4344 6851
rect 4072 6811 4130 6817
rect 4172 6820 4344 6848
rect 4172 6780 4200 6820
rect 4332 6817 4344 6820
rect 4378 6848 4390 6851
rect 5258 6848 5264 6860
rect 4378 6820 5264 6848
rect 4378 6817 4390 6820
rect 4332 6811 4390 6817
rect 5258 6808 5264 6820
rect 5316 6808 5322 6860
rect 3712 6752 4200 6780
rect 5552 6780 5580 6888
rect 6733 6885 6745 6919
rect 6779 6916 6791 6919
rect 8846 6916 8852 6928
rect 6779 6888 8852 6916
rect 6779 6885 6791 6888
rect 6733 6879 6791 6885
rect 8846 6876 8852 6888
rect 8904 6876 8910 6928
rect 10318 6916 10324 6928
rect 9784 6888 10324 6916
rect 5721 6851 5779 6857
rect 5721 6817 5733 6851
rect 5767 6848 5779 6851
rect 7098 6848 7104 6860
rect 5767 6820 7104 6848
rect 5767 6817 5779 6820
rect 5721 6811 5779 6817
rect 7098 6808 7104 6820
rect 7156 6808 7162 6860
rect 7377 6851 7435 6857
rect 7377 6817 7389 6851
rect 7423 6848 7435 6851
rect 7466 6848 7472 6860
rect 7423 6820 7472 6848
rect 7423 6817 7435 6820
rect 7377 6811 7435 6817
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 7650 6857 7656 6860
rect 7644 6848 7656 6857
rect 7563 6820 7656 6848
rect 7644 6811 7656 6820
rect 7708 6848 7714 6860
rect 8202 6848 8208 6860
rect 7708 6820 8208 6848
rect 7650 6808 7656 6811
rect 7708 6808 7714 6820
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 9784 6857 9812 6888
rect 10318 6876 10324 6888
rect 10376 6876 10382 6928
rect 10686 6876 10692 6928
rect 10744 6916 10750 6928
rect 16669 6919 16727 6925
rect 16669 6916 16681 6919
rect 10744 6888 16681 6916
rect 10744 6876 10750 6888
rect 16669 6885 16681 6888
rect 16715 6885 16727 6919
rect 16669 6879 16727 6885
rect 9769 6851 9827 6857
rect 9769 6817 9781 6851
rect 9815 6817 9827 6851
rect 9769 6811 9827 6817
rect 10036 6851 10094 6857
rect 10036 6817 10048 6851
rect 10082 6848 10094 6851
rect 11698 6848 11704 6860
rect 10082 6820 11704 6848
rect 10082 6817 10094 6820
rect 10036 6811 10094 6817
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 11882 6848 11888 6860
rect 11843 6820 11888 6848
rect 11882 6808 11888 6820
rect 11940 6808 11946 6860
rect 12066 6808 12072 6860
rect 12124 6848 12130 6860
rect 12894 6848 12900 6860
rect 12124 6820 12756 6848
rect 12855 6820 12900 6848
rect 12124 6808 12130 6820
rect 6546 6780 6552 6792
rect 5552 6752 6552 6780
rect 3712 6721 3740 6752
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6749 6883 6783
rect 6825 6743 6883 6749
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6780 7067 6783
rect 7193 6783 7251 6789
rect 7193 6780 7205 6783
rect 7055 6752 7205 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 7193 6749 7205 6752
rect 7239 6749 7251 6783
rect 7193 6743 7251 6749
rect 9033 6783 9091 6789
rect 9033 6749 9045 6783
rect 9079 6780 9091 6783
rect 9674 6780 9680 6792
rect 9079 6752 9680 6780
rect 9079 6749 9091 6752
rect 9033 6743 9091 6749
rect 3697 6715 3755 6721
rect 3697 6681 3709 6715
rect 3743 6681 3755 6715
rect 3697 6675 3755 6681
rect 5074 6672 5080 6724
rect 5132 6712 5138 6724
rect 5905 6715 5963 6721
rect 5905 6712 5917 6715
rect 5132 6684 5917 6712
rect 5132 6672 5138 6684
rect 5905 6681 5917 6684
rect 5951 6681 5963 6715
rect 5905 6675 5963 6681
rect 1394 6604 1400 6656
rect 1452 6644 1458 6656
rect 1857 6647 1915 6653
rect 1857 6644 1869 6647
rect 1452 6616 1869 6644
rect 1452 6604 1458 6616
rect 1857 6613 1869 6616
rect 1903 6613 1915 6647
rect 1857 6607 1915 6613
rect 4338 6604 4344 6656
rect 4396 6644 4402 6656
rect 5445 6647 5503 6653
rect 5445 6644 5457 6647
rect 4396 6616 5457 6644
rect 4396 6604 4402 6616
rect 5445 6613 5457 6616
rect 5491 6613 5503 6647
rect 6840 6644 6868 6743
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 12161 6783 12219 6789
rect 12161 6749 12173 6783
rect 12207 6780 12219 6783
rect 12250 6780 12256 6792
rect 12207 6752 12256 6780
rect 12207 6749 12219 6752
rect 12161 6743 12219 6749
rect 11517 6715 11575 6721
rect 11517 6681 11529 6715
rect 11563 6712 11575 6715
rect 11606 6712 11612 6724
rect 11563 6684 11612 6712
rect 11563 6681 11575 6684
rect 11517 6675 11575 6681
rect 11606 6672 11612 6684
rect 11664 6672 11670 6724
rect 11992 6712 12020 6743
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 12529 6715 12587 6721
rect 12529 6712 12541 6715
rect 11992 6684 12541 6712
rect 12529 6681 12541 6684
rect 12575 6681 12587 6715
rect 12529 6675 12587 6681
rect 8570 6644 8576 6656
rect 6840 6616 8576 6644
rect 5445 6607 5503 6613
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 11149 6647 11207 6653
rect 11149 6613 11161 6647
rect 11195 6644 11207 6647
rect 12250 6644 12256 6656
rect 11195 6616 12256 6644
rect 11195 6613 11207 6616
rect 11149 6607 11207 6613
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 12728 6644 12756 6820
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 13446 6808 13452 6860
rect 13504 6848 13510 6860
rect 13814 6857 13820 6860
rect 13541 6851 13599 6857
rect 13541 6848 13553 6851
rect 13504 6820 13553 6848
rect 13504 6808 13510 6820
rect 13541 6817 13553 6820
rect 13587 6817 13599 6851
rect 13808 6848 13820 6857
rect 13775 6820 13820 6848
rect 13541 6811 13599 6817
rect 13808 6811 13820 6820
rect 13814 6808 13820 6811
rect 13872 6808 13878 6860
rect 14090 6808 14096 6860
rect 14148 6848 14154 6860
rect 14148 6820 14596 6848
rect 14148 6808 14154 6820
rect 12986 6780 12992 6792
rect 12947 6752 12992 6780
rect 12986 6740 12992 6752
rect 13044 6740 13050 6792
rect 13078 6740 13084 6792
rect 13136 6780 13142 6792
rect 13173 6783 13231 6789
rect 13173 6780 13185 6783
rect 13136 6752 13185 6780
rect 13136 6740 13142 6752
rect 13173 6749 13185 6752
rect 13219 6780 13231 6783
rect 13357 6783 13415 6789
rect 13357 6780 13369 6783
rect 13219 6752 13369 6780
rect 13219 6749 13231 6752
rect 13173 6743 13231 6749
rect 13357 6749 13369 6752
rect 13403 6749 13415 6783
rect 14568 6780 14596 6820
rect 15562 6808 15568 6860
rect 15620 6848 15626 6860
rect 15749 6851 15807 6857
rect 15749 6848 15761 6851
rect 15620 6820 15761 6848
rect 15620 6808 15626 6820
rect 15749 6817 15761 6820
rect 15795 6817 15807 6851
rect 17865 6851 17923 6857
rect 17865 6848 17877 6851
rect 15749 6811 15807 6817
rect 15856 6820 17877 6848
rect 15856 6780 15884 6820
rect 17865 6817 17877 6820
rect 17911 6817 17923 6851
rect 17865 6811 17923 6817
rect 14568 6752 15884 6780
rect 15933 6783 15991 6789
rect 13357 6743 13415 6749
rect 15933 6749 15945 6783
rect 15979 6780 15991 6783
rect 16206 6780 16212 6792
rect 15979 6752 16212 6780
rect 15979 6749 15991 6752
rect 15933 6743 15991 6749
rect 16206 6740 16212 6752
rect 16264 6740 16270 6792
rect 16574 6740 16580 6792
rect 16632 6780 16638 6792
rect 16761 6783 16819 6789
rect 16761 6780 16773 6783
rect 16632 6752 16773 6780
rect 16632 6740 16638 6752
rect 16761 6749 16773 6752
rect 16807 6749 16819 6783
rect 16761 6743 16819 6749
rect 16853 6783 16911 6789
rect 16853 6749 16865 6783
rect 16899 6749 16911 6783
rect 16853 6743 16911 6749
rect 16868 6712 16896 6743
rect 18046 6712 18052 6724
rect 14476 6684 16896 6712
rect 18007 6684 18052 6712
rect 14476 6644 14504 6684
rect 18046 6672 18052 6684
rect 18104 6672 18110 6724
rect 15286 6644 15292 6656
rect 12728 6616 14504 6644
rect 15247 6616 15292 6644
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 16298 6644 16304 6656
rect 16259 6616 16304 6644
rect 16298 6604 16304 6616
rect 16356 6604 16362 6656
rect 1104 6554 18860 6576
rect 1104 6502 3947 6554
rect 3999 6502 4011 6554
rect 4063 6502 4075 6554
rect 4127 6502 4139 6554
rect 4191 6502 9878 6554
rect 9930 6502 9942 6554
rect 9994 6502 10006 6554
rect 10058 6502 10070 6554
rect 10122 6502 15808 6554
rect 15860 6502 15872 6554
rect 15924 6502 15936 6554
rect 15988 6502 16000 6554
rect 16052 6502 18860 6554
rect 1104 6480 18860 6502
rect 2682 6400 2688 6452
rect 2740 6400 2746 6452
rect 4522 6400 4528 6452
rect 4580 6440 4586 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 4580 6412 6561 6440
rect 4580 6400 4586 6412
rect 6549 6409 6561 6412
rect 6595 6409 6607 6443
rect 6549 6403 6607 6409
rect 7098 6400 7104 6452
rect 7156 6440 7162 6452
rect 8202 6440 8208 6452
rect 7156 6412 8064 6440
rect 8163 6412 8208 6440
rect 7156 6400 7162 6412
rect 2700 6372 2728 6400
rect 4062 6372 4068 6384
rect 1688 6344 4068 6372
rect 1688 6245 1716 6344
rect 4062 6332 4068 6344
rect 4120 6332 4126 6384
rect 4430 6332 4436 6384
rect 4488 6372 4494 6384
rect 5721 6375 5779 6381
rect 5721 6372 5733 6375
rect 4488 6344 5733 6372
rect 4488 6332 4494 6344
rect 5721 6341 5733 6344
rect 5767 6341 5779 6375
rect 5721 6335 5779 6341
rect 1946 6264 1952 6316
rect 2004 6304 2010 6316
rect 2685 6307 2743 6313
rect 2685 6304 2697 6307
rect 2004 6276 2697 6304
rect 2004 6264 2010 6276
rect 2685 6273 2697 6276
rect 2731 6273 2743 6307
rect 2685 6267 2743 6273
rect 2869 6307 2927 6313
rect 2869 6273 2881 6307
rect 2915 6304 2927 6307
rect 2958 6304 2964 6316
rect 2915 6276 2964 6304
rect 2915 6273 2927 6276
rect 2869 6267 2927 6273
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 4338 6304 4344 6316
rect 4299 6276 4344 6304
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 5258 6304 5264 6316
rect 5219 6276 5264 6304
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 6362 6304 6368 6316
rect 6323 6276 6368 6304
rect 6362 6264 6368 6276
rect 6420 6264 6426 6316
rect 8036 6304 8064 6412
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 8352 6412 10088 6440
rect 8352 6400 8358 6412
rect 10060 6372 10088 6412
rect 10318 6400 10324 6452
rect 10376 6440 10382 6452
rect 10781 6443 10839 6449
rect 10781 6440 10793 6443
rect 10376 6412 10793 6440
rect 10376 6400 10382 6412
rect 10781 6409 10793 6412
rect 10827 6409 10839 6443
rect 10781 6403 10839 6409
rect 11333 6443 11391 6449
rect 11333 6409 11345 6443
rect 11379 6440 11391 6443
rect 11882 6440 11888 6452
rect 11379 6412 11888 6440
rect 11379 6409 11391 6412
rect 11333 6403 11391 6409
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12710 6440 12716 6452
rect 11992 6412 12716 6440
rect 10505 6375 10563 6381
rect 10060 6344 10456 6372
rect 10428 6304 10456 6344
rect 10505 6341 10517 6375
rect 10551 6372 10563 6375
rect 11238 6372 11244 6384
rect 10551 6344 11244 6372
rect 10551 6341 10563 6344
rect 10505 6335 10563 6341
rect 11238 6332 11244 6344
rect 11296 6332 11302 6384
rect 11790 6332 11796 6384
rect 11848 6372 11854 6384
rect 11992 6372 12020 6412
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 12894 6400 12900 6452
rect 12952 6440 12958 6452
rect 13541 6443 13599 6449
rect 13541 6440 13553 6443
rect 12952 6412 13553 6440
rect 12952 6400 12958 6412
rect 13541 6409 13553 6412
rect 13587 6409 13599 6443
rect 13541 6403 13599 6409
rect 13722 6400 13728 6452
rect 13780 6440 13786 6452
rect 15654 6440 15660 6452
rect 13780 6412 15660 6440
rect 13780 6400 13786 6412
rect 15654 6400 15660 6412
rect 15712 6400 15718 6452
rect 18230 6440 18236 6452
rect 18191 6412 18236 6440
rect 18230 6400 18236 6412
rect 18288 6400 18294 6452
rect 11848 6344 12020 6372
rect 12161 6375 12219 6381
rect 11848 6332 11854 6344
rect 12161 6341 12173 6375
rect 12207 6372 12219 6375
rect 12618 6372 12624 6384
rect 12207 6344 12624 6372
rect 12207 6341 12219 6344
rect 12161 6335 12219 6341
rect 12618 6332 12624 6344
rect 12676 6332 12682 6384
rect 12986 6332 12992 6384
rect 13044 6372 13050 6384
rect 15565 6375 15623 6381
rect 15565 6372 15577 6375
rect 13044 6344 15577 6372
rect 13044 6332 13050 6344
rect 15565 6341 15577 6344
rect 15611 6341 15623 6375
rect 15565 6335 15623 6341
rect 15930 6332 15936 6384
rect 15988 6372 15994 6384
rect 17954 6372 17960 6384
rect 15988 6344 17960 6372
rect 15988 6332 15994 6344
rect 17954 6332 17960 6344
rect 18012 6332 18018 6384
rect 10597 6307 10655 6313
rect 10597 6304 10609 6307
rect 8036 6276 9260 6304
rect 10428 6276 10609 6304
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6205 1731 6239
rect 1673 6199 1731 6205
rect 1854 6196 1860 6248
rect 1912 6236 1918 6248
rect 2593 6239 2651 6245
rect 2593 6236 2605 6239
rect 1912 6208 2605 6236
rect 1912 6196 1918 6208
rect 2593 6205 2605 6208
rect 2639 6205 2651 6239
rect 2593 6199 2651 6205
rect 3237 6239 3295 6245
rect 3237 6205 3249 6239
rect 3283 6236 3295 6239
rect 4982 6236 4988 6248
rect 3283 6208 4988 6236
rect 3283 6205 3295 6208
rect 3237 6199 3295 6205
rect 4982 6196 4988 6208
rect 5040 6196 5046 6248
rect 5442 6196 5448 6248
rect 5500 6236 5506 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 5500 6208 6837 6236
rect 5500 6196 5506 6208
rect 6825 6205 6837 6208
rect 6871 6236 6883 6239
rect 7466 6236 7472 6248
rect 6871 6208 7472 6236
rect 6871 6205 6883 6208
rect 6825 6199 6883 6205
rect 7466 6196 7472 6208
rect 7524 6236 7530 6248
rect 8478 6236 8484 6248
rect 7524 6208 8484 6236
rect 7524 6196 7530 6208
rect 8478 6196 8484 6208
rect 8536 6236 8542 6248
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 8536 6208 9137 6236
rect 8536 6196 8542 6208
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 9232 6236 9260 6276
rect 10597 6273 10609 6276
rect 10643 6273 10655 6307
rect 11330 6304 11336 6316
rect 10597 6267 10655 6273
rect 10796 6276 11336 6304
rect 10796 6236 10824 6276
rect 11330 6264 11336 6276
rect 11388 6264 11394 6316
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11756 6276 11897 6304
rect 11756 6264 11762 6276
rect 11885 6273 11897 6276
rect 11931 6304 11943 6307
rect 13078 6304 13084 6316
rect 11931 6276 13084 6304
rect 11931 6273 11943 6276
rect 11885 6267 11943 6273
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 13173 6307 13231 6313
rect 13173 6273 13185 6307
rect 13219 6304 13231 6307
rect 13538 6304 13544 6316
rect 13219 6276 13544 6304
rect 13219 6273 13231 6276
rect 13173 6267 13231 6273
rect 13538 6264 13544 6276
rect 13596 6304 13602 6316
rect 13814 6304 13820 6316
rect 13596 6276 13820 6304
rect 13596 6264 13602 6276
rect 13814 6264 13820 6276
rect 13872 6304 13878 6316
rect 14185 6307 14243 6313
rect 14185 6304 14197 6307
rect 13872 6276 14197 6304
rect 13872 6264 13878 6276
rect 14185 6273 14197 6276
rect 14231 6273 14243 6307
rect 15102 6304 15108 6316
rect 15063 6276 15108 6304
rect 14185 6267 14243 6273
rect 10962 6236 10968 6248
rect 9232 6208 10824 6236
rect 10923 6208 10968 6236
rect 9125 6199 9183 6205
rect 10962 6196 10968 6208
rect 11020 6196 11026 6248
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 11440 6208 12173 6236
rect 2958 6168 2964 6180
rect 1872 6140 2964 6168
rect 1872 6109 1900 6140
rect 2958 6128 2964 6140
rect 3016 6128 3022 6180
rect 3602 6128 3608 6180
rect 3660 6168 3666 6180
rect 4065 6171 4123 6177
rect 4065 6168 4077 6171
rect 3660 6140 4077 6168
rect 3660 6128 3666 6140
rect 4065 6137 4077 6140
rect 4111 6137 4123 6171
rect 4065 6131 4123 6137
rect 5902 6128 5908 6180
rect 5960 6168 5966 6180
rect 6181 6171 6239 6177
rect 6181 6168 6193 6171
rect 5960 6140 6193 6168
rect 5960 6128 5966 6140
rect 6181 6137 6193 6140
rect 6227 6137 6239 6171
rect 6181 6131 6239 6137
rect 6730 6128 6736 6180
rect 6788 6168 6794 6180
rect 9398 6177 9404 6180
rect 7070 6171 7128 6177
rect 7070 6168 7082 6171
rect 6788 6140 7082 6168
rect 6788 6128 6794 6140
rect 7070 6137 7082 6140
rect 7116 6137 7128 6171
rect 9392 6168 9404 6177
rect 7070 6131 7128 6137
rect 7208 6140 8616 6168
rect 9359 6140 9404 6168
rect 1857 6103 1915 6109
rect 1857 6069 1869 6103
rect 1903 6069 1915 6103
rect 1857 6063 1915 6069
rect 2225 6103 2283 6109
rect 2225 6069 2237 6103
rect 2271 6100 2283 6103
rect 2314 6100 2320 6112
rect 2271 6072 2320 6100
rect 2271 6069 2283 6072
rect 2225 6063 2283 6069
rect 2314 6060 2320 6072
rect 2372 6060 2378 6112
rect 3694 6100 3700 6112
rect 3655 6072 3700 6100
rect 3694 6060 3700 6072
rect 3752 6060 3758 6112
rect 4157 6103 4215 6109
rect 4157 6069 4169 6103
rect 4203 6100 4215 6103
rect 4709 6103 4767 6109
rect 4709 6100 4721 6103
rect 4203 6072 4721 6100
rect 4203 6069 4215 6072
rect 4157 6063 4215 6069
rect 4709 6069 4721 6072
rect 4755 6069 4767 6103
rect 4709 6063 4767 6069
rect 4890 6060 4896 6112
rect 4948 6100 4954 6112
rect 5077 6103 5135 6109
rect 5077 6100 5089 6103
rect 4948 6072 5089 6100
rect 4948 6060 4954 6072
rect 5077 6069 5089 6072
rect 5123 6069 5135 6103
rect 5077 6063 5135 6069
rect 5169 6103 5227 6109
rect 5169 6069 5181 6103
rect 5215 6100 5227 6103
rect 5258 6100 5264 6112
rect 5215 6072 5264 6100
rect 5215 6069 5227 6072
rect 5169 6063 5227 6069
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 6086 6100 6092 6112
rect 6047 6072 6092 6100
rect 6086 6060 6092 6072
rect 6144 6060 6150 6112
rect 6549 6103 6607 6109
rect 6549 6069 6561 6103
rect 6595 6100 6607 6103
rect 7208 6100 7236 6140
rect 6595 6072 7236 6100
rect 6595 6069 6607 6072
rect 6549 6063 6607 6069
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 8481 6103 8539 6109
rect 8481 6100 8493 6103
rect 7340 6072 8493 6100
rect 7340 6060 7346 6072
rect 8481 6069 8493 6072
rect 8527 6069 8539 6103
rect 8588 6100 8616 6140
rect 9392 6131 9404 6140
rect 9398 6128 9404 6131
rect 9456 6128 9462 6180
rect 10597 6171 10655 6177
rect 10597 6137 10609 6171
rect 10643 6168 10655 6171
rect 11440 6168 11468 6208
rect 12161 6205 12173 6208
rect 12207 6205 12219 6239
rect 12161 6199 12219 6205
rect 12618 6196 12624 6248
rect 12676 6236 12682 6248
rect 13722 6236 13728 6248
rect 12676 6208 13728 6236
rect 12676 6196 12682 6208
rect 13722 6196 13728 6208
rect 13780 6196 13786 6248
rect 13906 6236 13912 6248
rect 13867 6208 13912 6236
rect 13906 6196 13912 6208
rect 13964 6196 13970 6248
rect 14200 6236 14228 6267
rect 15102 6264 15108 6276
rect 15160 6264 15166 6316
rect 16117 6307 16175 6313
rect 16117 6273 16129 6307
rect 16163 6273 16175 6307
rect 16117 6267 16175 6273
rect 16132 6236 16160 6267
rect 14200 6208 16160 6236
rect 17034 6196 17040 6248
rect 17092 6236 17098 6248
rect 17405 6239 17463 6245
rect 17405 6236 17417 6239
rect 17092 6208 17417 6236
rect 17092 6196 17098 6208
rect 17405 6205 17417 6208
rect 17451 6205 17463 6239
rect 17405 6199 17463 6205
rect 17770 6196 17776 6248
rect 17828 6236 17834 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 17828 6208 18061 6236
rect 17828 6196 17834 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 10643 6140 11468 6168
rect 10643 6137 10655 6140
rect 10597 6131 10655 6137
rect 11514 6128 11520 6180
rect 11572 6168 11578 6180
rect 11701 6171 11759 6177
rect 11701 6168 11713 6171
rect 11572 6140 11713 6168
rect 11572 6128 11578 6140
rect 11701 6137 11713 6140
rect 11747 6168 11759 6171
rect 17310 6168 17316 6180
rect 11747 6140 17316 6168
rect 11747 6137 11759 6140
rect 11701 6131 11759 6137
rect 17310 6128 17316 6140
rect 17368 6128 17374 6180
rect 11606 6100 11612 6112
rect 8588 6072 11612 6100
rect 8481 6063 8539 6069
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 11793 6103 11851 6109
rect 11793 6069 11805 6103
rect 11839 6100 11851 6103
rect 12529 6103 12587 6109
rect 12529 6100 12541 6103
rect 11839 6072 12541 6100
rect 11839 6069 11851 6072
rect 11793 6063 11851 6069
rect 12529 6069 12541 6072
rect 12575 6069 12587 6103
rect 12529 6063 12587 6069
rect 12710 6060 12716 6112
rect 12768 6100 12774 6112
rect 12897 6103 12955 6109
rect 12897 6100 12909 6103
rect 12768 6072 12909 6100
rect 12768 6060 12774 6072
rect 12897 6069 12909 6072
rect 12943 6069 12955 6103
rect 12897 6063 12955 6069
rect 12989 6103 13047 6109
rect 12989 6069 13001 6103
rect 13035 6100 13047 6103
rect 13354 6100 13360 6112
rect 13035 6072 13360 6100
rect 13035 6069 13047 6072
rect 12989 6063 13047 6069
rect 13354 6060 13360 6072
rect 13412 6100 13418 6112
rect 13814 6100 13820 6112
rect 13412 6072 13820 6100
rect 13412 6060 13418 6072
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 13906 6060 13912 6112
rect 13964 6100 13970 6112
rect 14001 6103 14059 6109
rect 14001 6100 14013 6103
rect 13964 6072 14013 6100
rect 13964 6060 13970 6072
rect 14001 6069 14013 6072
rect 14047 6100 14059 6103
rect 14182 6100 14188 6112
rect 14047 6072 14188 6100
rect 14047 6069 14059 6072
rect 14001 6063 14059 6069
rect 14182 6060 14188 6072
rect 14240 6060 14246 6112
rect 14550 6100 14556 6112
rect 14511 6072 14556 6100
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 14918 6100 14924 6112
rect 14879 6072 14924 6100
rect 14918 6060 14924 6072
rect 14976 6060 14982 6112
rect 15013 6103 15071 6109
rect 15013 6069 15025 6103
rect 15059 6100 15071 6103
rect 15470 6100 15476 6112
rect 15059 6072 15476 6100
rect 15059 6069 15071 6072
rect 15013 6063 15071 6069
rect 15470 6060 15476 6072
rect 15528 6060 15534 6112
rect 15930 6100 15936 6112
rect 15891 6072 15936 6100
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 16025 6103 16083 6109
rect 16025 6069 16037 6103
rect 16071 6100 16083 6103
rect 16390 6100 16396 6112
rect 16071 6072 16396 6100
rect 16071 6069 16083 6072
rect 16025 6063 16083 6069
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 17586 6100 17592 6112
rect 17547 6072 17592 6100
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 1104 6010 18860 6032
rect 1104 5958 6912 6010
rect 6964 5958 6976 6010
rect 7028 5958 7040 6010
rect 7092 5958 7104 6010
rect 7156 5958 12843 6010
rect 12895 5958 12907 6010
rect 12959 5958 12971 6010
rect 13023 5958 13035 6010
rect 13087 5958 18860 6010
rect 1104 5936 18860 5958
rect 4065 5899 4123 5905
rect 4065 5865 4077 5899
rect 4111 5896 4123 5899
rect 6086 5896 6092 5908
rect 4111 5868 6092 5896
rect 4111 5865 4123 5868
rect 4065 5859 4123 5865
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 6730 5856 6736 5908
rect 6788 5896 6794 5908
rect 6825 5899 6883 5905
rect 6825 5896 6837 5899
rect 6788 5868 6837 5896
rect 6788 5856 6794 5868
rect 6825 5865 6837 5868
rect 6871 5865 6883 5899
rect 6825 5859 6883 5865
rect 6917 5899 6975 5905
rect 6917 5865 6929 5899
rect 6963 5896 6975 5899
rect 8018 5896 8024 5908
rect 6963 5868 8024 5896
rect 6963 5865 6975 5868
rect 6917 5859 6975 5865
rect 8018 5856 8024 5868
rect 8076 5896 8082 5908
rect 9309 5899 9367 5905
rect 9309 5896 9321 5899
rect 8076 5868 9321 5896
rect 8076 5856 8082 5868
rect 9309 5865 9321 5868
rect 9355 5865 9367 5899
rect 9309 5859 9367 5865
rect 10962 5856 10968 5908
rect 11020 5896 11026 5908
rect 11885 5899 11943 5905
rect 11885 5896 11897 5899
rect 11020 5868 11897 5896
rect 11020 5856 11026 5868
rect 11885 5865 11897 5868
rect 11931 5896 11943 5899
rect 14185 5899 14243 5905
rect 11931 5868 14044 5896
rect 11931 5865 11943 5868
rect 11885 5859 11943 5865
rect 1848 5831 1906 5837
rect 1848 5797 1860 5831
rect 1894 5828 1906 5831
rect 4338 5828 4344 5840
rect 1894 5800 4344 5828
rect 1894 5797 1906 5800
rect 1848 5791 1906 5797
rect 4338 5788 4344 5800
rect 4396 5788 4402 5840
rect 4525 5831 4583 5837
rect 4525 5797 4537 5831
rect 4571 5828 4583 5831
rect 5166 5828 5172 5840
rect 4571 5800 5172 5828
rect 4571 5797 4583 5800
rect 4525 5791 4583 5797
rect 2682 5720 2688 5772
rect 2740 5760 2746 5772
rect 3234 5760 3240 5772
rect 2740 5732 3240 5760
rect 2740 5720 2746 5732
rect 3234 5720 3240 5732
rect 3292 5720 3298 5772
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 4212 5732 4445 5760
rect 4212 5720 4218 5732
rect 4433 5729 4445 5732
rect 4479 5729 4491 5763
rect 4433 5723 4491 5729
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1544 5664 1593 5692
rect 1544 5652 1550 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4540 5692 4568 5791
rect 5166 5788 5172 5800
rect 5224 5788 5230 5840
rect 10318 5828 10324 5840
rect 5276 5800 7880 5828
rect 4706 5720 4712 5772
rect 4764 5760 4770 5772
rect 5276 5769 5304 5800
rect 5261 5763 5319 5769
rect 5261 5760 5273 5763
rect 4764 5732 5273 5760
rect 4764 5720 4770 5732
rect 5261 5729 5273 5732
rect 5307 5729 5319 5763
rect 5442 5760 5448 5772
rect 5403 5732 5448 5760
rect 5261 5723 5319 5729
rect 5442 5720 5448 5732
rect 5500 5720 5506 5772
rect 5712 5763 5770 5769
rect 5712 5729 5724 5763
rect 5758 5760 5770 5763
rect 6917 5763 6975 5769
rect 6917 5760 6929 5763
rect 5758 5732 6929 5760
rect 5758 5729 5770 5732
rect 5712 5723 5770 5729
rect 6917 5729 6929 5732
rect 6963 5729 6975 5763
rect 7098 5760 7104 5772
rect 7059 5732 7104 5760
rect 6917 5723 6975 5729
rect 7098 5720 7104 5732
rect 7156 5720 7162 5772
rect 7852 5769 7880 5800
rect 9968 5800 10324 5828
rect 7829 5763 7887 5769
rect 7829 5729 7841 5763
rect 7875 5729 7887 5763
rect 7829 5723 7887 5729
rect 8196 5763 8254 5769
rect 8196 5729 8208 5763
rect 8242 5760 8254 5763
rect 9306 5760 9312 5772
rect 8242 5732 9312 5760
rect 8242 5729 8254 5732
rect 8196 5723 8254 5729
rect 9306 5720 9312 5732
rect 9364 5720 9370 5772
rect 9968 5769 9996 5800
rect 10318 5788 10324 5800
rect 10376 5788 10382 5840
rect 12158 5828 12164 5840
rect 12084 5800 12164 5828
rect 9953 5763 10011 5769
rect 9953 5729 9965 5763
rect 9999 5729 10011 5763
rect 9953 5723 10011 5729
rect 10220 5763 10278 5769
rect 10220 5729 10232 5763
rect 10266 5760 10278 5763
rect 11238 5760 11244 5772
rect 10266 5732 11244 5760
rect 10266 5729 10278 5732
rect 10220 5723 10278 5729
rect 11238 5720 11244 5732
rect 11296 5720 11302 5772
rect 12084 5769 12112 5800
rect 12158 5788 12164 5800
rect 12216 5788 12222 5840
rect 12069 5763 12127 5769
rect 12069 5729 12081 5763
rect 12115 5729 12127 5763
rect 12069 5723 12127 5729
rect 12428 5763 12486 5769
rect 12428 5729 12440 5763
rect 12474 5760 12486 5763
rect 13722 5760 13728 5772
rect 12474 5732 13728 5760
rect 12474 5729 12486 5732
rect 12428 5723 12486 5729
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 14016 5769 14044 5868
rect 14185 5865 14197 5899
rect 14231 5896 14243 5899
rect 14918 5896 14924 5908
rect 14231 5868 14924 5896
rect 14231 5865 14243 5868
rect 14185 5859 14243 5865
rect 14918 5856 14924 5868
rect 14976 5856 14982 5908
rect 18046 5896 18052 5908
rect 18007 5868 18052 5896
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 14090 5788 14096 5840
rect 14148 5828 14154 5840
rect 14642 5828 14648 5840
rect 14148 5800 14648 5828
rect 14148 5788 14154 5800
rect 14642 5788 14648 5800
rect 14700 5788 14706 5840
rect 14001 5763 14059 5769
rect 14001 5729 14013 5763
rect 14047 5729 14059 5763
rect 14001 5723 14059 5729
rect 14553 5763 14611 5769
rect 14553 5729 14565 5763
rect 14599 5760 14611 5763
rect 15289 5763 15347 5769
rect 15289 5760 15301 5763
rect 14599 5732 15301 5760
rect 14599 5729 14611 5732
rect 14553 5723 14611 5729
rect 15289 5729 15301 5732
rect 15335 5729 15347 5763
rect 17310 5760 17316 5772
rect 17271 5732 17316 5760
rect 15289 5723 15347 5729
rect 17310 5720 17316 5732
rect 17368 5720 17374 5772
rect 17865 5763 17923 5769
rect 17865 5729 17877 5763
rect 17911 5729 17923 5763
rect 17865 5723 17923 5729
rect 4120 5664 4568 5692
rect 4617 5695 4675 5701
rect 4120 5652 4126 5664
rect 4617 5661 4629 5695
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 4338 5584 4344 5636
rect 4396 5624 4402 5636
rect 4632 5624 4660 5655
rect 4982 5652 4988 5704
rect 5040 5692 5046 5704
rect 5350 5692 5356 5704
rect 5040 5664 5356 5692
rect 5040 5652 5046 5664
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 7929 5695 7987 5701
rect 7929 5692 7941 5695
rect 7760 5664 7941 5692
rect 4396 5596 4660 5624
rect 4724 5596 5212 5624
rect 4396 5584 4402 5596
rect 2961 5559 3019 5565
rect 2961 5525 2973 5559
rect 3007 5556 3019 5559
rect 3142 5556 3148 5568
rect 3007 5528 3148 5556
rect 3007 5525 3019 5528
rect 2961 5519 3019 5525
rect 3142 5516 3148 5528
rect 3200 5516 3206 5568
rect 3418 5556 3424 5568
rect 3379 5528 3424 5556
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 3786 5516 3792 5568
rect 3844 5556 3850 5568
rect 4724 5556 4752 5596
rect 3844 5528 4752 5556
rect 3844 5516 3850 5528
rect 4798 5516 4804 5568
rect 4856 5556 4862 5568
rect 5077 5559 5135 5565
rect 5077 5556 5089 5559
rect 4856 5528 5089 5556
rect 4856 5516 4862 5528
rect 5077 5525 5089 5528
rect 5123 5525 5135 5559
rect 5184 5556 5212 5596
rect 7760 5568 7788 5664
rect 7929 5661 7941 5664
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 12158 5652 12164 5704
rect 12216 5692 12222 5704
rect 14829 5695 14887 5701
rect 12216 5664 12261 5692
rect 12216 5652 12222 5664
rect 14829 5661 14841 5695
rect 14875 5692 14887 5695
rect 15010 5692 15016 5704
rect 14875 5664 15016 5692
rect 14875 5661 14887 5664
rect 14829 5655 14887 5661
rect 15010 5652 15016 5664
rect 15068 5652 15074 5704
rect 13538 5624 13544 5636
rect 13499 5596 13544 5624
rect 13538 5584 13544 5596
rect 13596 5584 13602 5636
rect 13630 5584 13636 5636
rect 13688 5624 13694 5636
rect 17880 5624 17908 5723
rect 13688 5596 17908 5624
rect 13688 5584 13694 5596
rect 7285 5559 7343 5565
rect 7285 5556 7297 5559
rect 5184 5528 7297 5556
rect 5077 5519 5135 5525
rect 7285 5525 7297 5528
rect 7331 5525 7343 5559
rect 7285 5519 7343 5525
rect 7466 5516 7472 5568
rect 7524 5556 7530 5568
rect 7653 5559 7711 5565
rect 7653 5556 7665 5559
rect 7524 5528 7665 5556
rect 7524 5516 7530 5528
rect 7653 5525 7665 5528
rect 7699 5556 7711 5559
rect 7742 5556 7748 5568
rect 7699 5528 7748 5556
rect 7699 5525 7711 5528
rect 7653 5519 7711 5525
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 11330 5556 11336 5568
rect 11291 5528 11336 5556
rect 11330 5516 11336 5528
rect 11388 5516 11394 5568
rect 12158 5516 12164 5568
rect 12216 5556 12222 5568
rect 12434 5556 12440 5568
rect 12216 5528 12440 5556
rect 12216 5516 12222 5528
rect 12434 5516 12440 5528
rect 12492 5556 12498 5568
rect 13446 5556 13452 5568
rect 12492 5528 13452 5556
rect 12492 5516 12498 5528
rect 13446 5516 13452 5528
rect 13504 5556 13510 5568
rect 13817 5559 13875 5565
rect 13817 5556 13829 5559
rect 13504 5528 13829 5556
rect 13504 5516 13510 5528
rect 13817 5525 13829 5528
rect 13863 5525 13875 5559
rect 17494 5556 17500 5568
rect 17455 5528 17500 5556
rect 13817 5519 13875 5525
rect 17494 5516 17500 5528
rect 17552 5516 17558 5568
rect 1104 5466 18860 5488
rect 1104 5414 3947 5466
rect 3999 5414 4011 5466
rect 4063 5414 4075 5466
rect 4127 5414 4139 5466
rect 4191 5414 9878 5466
rect 9930 5414 9942 5466
rect 9994 5414 10006 5466
rect 10058 5414 10070 5466
rect 10122 5414 15808 5466
rect 15860 5414 15872 5466
rect 15924 5414 15936 5466
rect 15988 5414 16000 5466
rect 16052 5414 18860 5466
rect 1104 5392 18860 5414
rect 3694 5312 3700 5364
rect 3752 5352 3758 5364
rect 4982 5352 4988 5364
rect 3752 5324 4988 5352
rect 3752 5312 3758 5324
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 5074 5312 5080 5364
rect 5132 5352 5138 5364
rect 6181 5355 6239 5361
rect 6181 5352 6193 5355
rect 5132 5324 6193 5352
rect 5132 5312 5138 5324
rect 6181 5321 6193 5324
rect 6227 5321 6239 5355
rect 6181 5315 6239 5321
rect 6362 5312 6368 5364
rect 6420 5352 6426 5364
rect 8846 5352 8852 5364
rect 6420 5324 7420 5352
rect 8807 5324 8852 5352
rect 6420 5312 6426 5324
rect 3973 5287 4031 5293
rect 3973 5253 3985 5287
rect 4019 5284 4031 5287
rect 4019 5256 7328 5284
rect 4019 5253 4031 5256
rect 3973 5247 4031 5253
rect 4338 5176 4344 5228
rect 4396 5216 4402 5228
rect 4525 5219 4583 5225
rect 4525 5216 4537 5219
rect 4396 5188 4537 5216
rect 4396 5176 4402 5188
rect 4525 5185 4537 5188
rect 4571 5216 4583 5219
rect 5537 5219 5595 5225
rect 5537 5216 5549 5219
rect 4571 5188 5549 5216
rect 4571 5185 4583 5188
rect 4525 5179 4583 5185
rect 5537 5185 5549 5188
rect 5583 5185 5595 5219
rect 7098 5216 7104 5228
rect 5537 5179 5595 5185
rect 5920 5188 7104 5216
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 1486 5148 1492 5160
rect 1443 5120 1492 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 1486 5108 1492 5120
rect 1544 5148 1550 5160
rect 2038 5148 2044 5160
rect 1544 5120 2044 5148
rect 1544 5108 1550 5120
rect 2038 5108 2044 5120
rect 2096 5108 2102 5160
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5148 3111 5151
rect 5350 5148 5356 5160
rect 3099 5120 3372 5148
rect 5311 5120 5356 5148
rect 3099 5117 3111 5120
rect 3053 5111 3111 5117
rect 1664 5083 1722 5089
rect 1664 5049 1676 5083
rect 1710 5080 1722 5083
rect 3142 5080 3148 5092
rect 1710 5052 3148 5080
rect 1710 5049 1722 5052
rect 1664 5043 1722 5049
rect 3142 5040 3148 5052
rect 3200 5040 3206 5092
rect 3344 5080 3372 5120
rect 5350 5108 5356 5120
rect 5408 5108 5414 5160
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5148 5503 5151
rect 5920 5148 5948 5188
rect 7098 5176 7104 5188
rect 7156 5176 7162 5228
rect 7300 5225 7328 5256
rect 7392 5225 7420 5324
rect 8846 5312 8852 5324
rect 8904 5312 8910 5364
rect 9582 5352 9588 5364
rect 9140 5324 9588 5352
rect 7466 5244 7472 5296
rect 7524 5284 7530 5296
rect 9140 5284 9168 5324
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 9861 5355 9919 5361
rect 9861 5352 9873 5355
rect 9824 5324 9873 5352
rect 9824 5312 9830 5324
rect 9861 5321 9873 5324
rect 9907 5321 9919 5355
rect 9861 5315 9919 5321
rect 10502 5312 10508 5364
rect 10560 5352 10566 5364
rect 10873 5355 10931 5361
rect 10873 5352 10885 5355
rect 10560 5324 10885 5352
rect 10560 5312 10566 5324
rect 10873 5321 10885 5324
rect 10919 5321 10931 5355
rect 10873 5315 10931 5321
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 11204 5324 13676 5352
rect 11204 5312 11210 5324
rect 7524 5256 9168 5284
rect 7524 5244 7530 5256
rect 9214 5244 9220 5296
rect 9272 5284 9278 5296
rect 12250 5284 12256 5296
rect 9272 5256 12256 5284
rect 9272 5244 9278 5256
rect 12250 5244 12256 5256
rect 12308 5244 12314 5296
rect 13648 5284 13676 5324
rect 13722 5312 13728 5364
rect 13780 5352 13786 5364
rect 13817 5355 13875 5361
rect 13817 5352 13829 5355
rect 13780 5324 13829 5352
rect 13780 5312 13786 5324
rect 13817 5321 13829 5324
rect 13863 5321 13875 5355
rect 13817 5315 13875 5321
rect 14090 5312 14096 5364
rect 14148 5312 14154 5364
rect 14826 5312 14832 5364
rect 14884 5352 14890 5364
rect 14884 5324 15056 5352
rect 14884 5312 14890 5324
rect 14108 5284 14136 5312
rect 13648 5256 14136 5284
rect 15028 5284 15056 5324
rect 15470 5312 15476 5364
rect 15528 5352 15534 5364
rect 15749 5355 15807 5361
rect 15749 5352 15761 5355
rect 15528 5324 15761 5352
rect 15528 5312 15534 5324
rect 15749 5321 15761 5324
rect 15795 5321 15807 5355
rect 15749 5315 15807 5321
rect 15028 5256 17448 5284
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 7377 5219 7435 5225
rect 7377 5185 7389 5219
rect 7423 5185 7435 5219
rect 7377 5179 7435 5185
rect 7650 5176 7656 5228
rect 7708 5216 7714 5228
rect 8294 5216 8300 5228
rect 7708 5188 8300 5216
rect 7708 5176 7714 5188
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 8481 5219 8539 5225
rect 8481 5185 8493 5219
rect 8527 5216 8539 5219
rect 8662 5216 8668 5228
rect 8527 5188 8668 5216
rect 8527 5185 8539 5188
rect 8481 5179 8539 5185
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 9306 5176 9312 5228
rect 9364 5216 9370 5228
rect 9401 5219 9459 5225
rect 9401 5216 9413 5219
rect 9364 5188 9413 5216
rect 9364 5176 9370 5188
rect 9401 5185 9413 5188
rect 9447 5216 9459 5219
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 9447 5188 10425 5216
rect 9447 5185 9459 5188
rect 9401 5179 9459 5185
rect 10413 5185 10425 5188
rect 10459 5216 10471 5219
rect 11425 5219 11483 5225
rect 11425 5216 11437 5219
rect 10459 5188 11437 5216
rect 10459 5185 10471 5188
rect 10413 5179 10471 5185
rect 11425 5185 11437 5188
rect 11471 5185 11483 5219
rect 12434 5216 12440 5228
rect 12395 5188 12440 5216
rect 11425 5179 11483 5185
rect 12434 5176 12440 5188
rect 12492 5176 12498 5228
rect 13446 5176 13452 5228
rect 13504 5216 13510 5228
rect 14093 5219 14151 5225
rect 14093 5216 14105 5219
rect 13504 5188 14105 5216
rect 13504 5176 13510 5188
rect 14093 5185 14105 5188
rect 14139 5185 14151 5219
rect 14093 5179 14151 5185
rect 15930 5176 15936 5228
rect 15988 5216 15994 5228
rect 16301 5219 16359 5225
rect 16301 5216 16313 5219
rect 15988 5188 16313 5216
rect 15988 5176 15994 5188
rect 16301 5185 16313 5188
rect 16347 5185 16359 5219
rect 16301 5179 16359 5185
rect 5491 5120 5948 5148
rect 5997 5151 6055 5157
rect 5491 5117 5503 5120
rect 5445 5111 5503 5117
rect 5997 5117 6009 5151
rect 6043 5148 6055 5151
rect 6270 5148 6276 5160
rect 6043 5120 6276 5148
rect 6043 5117 6055 5120
rect 5997 5111 6055 5117
rect 6270 5108 6276 5120
rect 6328 5108 6334 5160
rect 7116 5148 7144 5176
rect 7116 5120 9444 5148
rect 4522 5080 4528 5092
rect 3344 5052 4528 5080
rect 4522 5040 4528 5052
rect 4580 5040 4586 5092
rect 7193 5083 7251 5089
rect 7193 5080 7205 5083
rect 5000 5052 7205 5080
rect 2774 4972 2780 5024
rect 2832 5012 2838 5024
rect 3234 5012 3240 5024
rect 2832 4984 2877 5012
rect 3195 4984 3240 5012
rect 2832 4972 2838 4984
rect 3234 4972 3240 4984
rect 3292 4972 3298 5024
rect 4338 5012 4344 5024
rect 4299 4984 4344 5012
rect 4338 4972 4344 4984
rect 4396 4972 4402 5024
rect 4430 4972 4436 5024
rect 4488 5012 4494 5024
rect 5000 5021 5028 5052
rect 7193 5049 7205 5052
rect 7239 5049 7251 5083
rect 9309 5083 9367 5089
rect 9309 5080 9321 5083
rect 7193 5043 7251 5049
rect 7852 5052 9321 5080
rect 4985 5015 5043 5021
rect 4488 4984 4533 5012
rect 4488 4972 4494 4984
rect 4985 4981 4997 5015
rect 5031 4981 5043 5015
rect 4985 4975 5043 4981
rect 5166 4972 5172 5024
rect 5224 5012 5230 5024
rect 7852 5021 7880 5052
rect 9309 5049 9321 5052
rect 9355 5049 9367 5083
rect 9416 5080 9444 5120
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 11241 5151 11299 5157
rect 11241 5148 11253 5151
rect 9732 5120 11253 5148
rect 9732 5108 9738 5120
rect 11241 5117 11253 5120
rect 11287 5117 11299 5151
rect 11241 5111 11299 5117
rect 11514 5108 11520 5160
rect 11572 5148 11578 5160
rect 13630 5148 13636 5160
rect 11572 5120 13636 5148
rect 11572 5108 11578 5120
rect 13630 5108 13636 5120
rect 13688 5108 13694 5160
rect 13814 5108 13820 5160
rect 13872 5148 13878 5160
rect 14826 5148 14832 5160
rect 13872 5120 14832 5148
rect 13872 5108 13878 5120
rect 14826 5108 14832 5120
rect 14884 5108 14890 5160
rect 17420 5157 17448 5256
rect 17405 5151 17463 5157
rect 17405 5117 17417 5151
rect 17451 5117 17463 5151
rect 17405 5111 17463 5117
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5148 18107 5151
rect 18322 5148 18328 5160
rect 18095 5120 18328 5148
rect 18095 5117 18107 5120
rect 18049 5111 18107 5117
rect 18322 5108 18328 5120
rect 18380 5108 18386 5160
rect 11146 5080 11152 5092
rect 9416 5052 11152 5080
rect 9309 5043 9367 5049
rect 11146 5040 11152 5052
rect 11204 5080 11210 5092
rect 14366 5089 14372 5092
rect 11333 5083 11391 5089
rect 11333 5080 11345 5083
rect 11204 5052 11345 5080
rect 11204 5040 11210 5052
rect 11333 5049 11345 5052
rect 11379 5049 11391 5083
rect 11333 5043 11391 5049
rect 12704 5083 12762 5089
rect 12704 5049 12716 5083
rect 12750 5049 12762 5083
rect 12704 5043 12762 5049
rect 14360 5043 14372 5089
rect 14424 5080 14430 5092
rect 16114 5080 16120 5092
rect 14424 5052 14460 5080
rect 16027 5052 16120 5080
rect 6825 5015 6883 5021
rect 6825 5012 6837 5015
rect 5224 4984 6837 5012
rect 5224 4972 5230 4984
rect 6825 4981 6837 4984
rect 6871 4981 6883 5015
rect 6825 4975 6883 4981
rect 7837 5015 7895 5021
rect 7837 4981 7849 5015
rect 7883 4981 7895 5015
rect 8202 5012 8208 5024
rect 8163 4984 8208 5012
rect 7837 4975 7895 4981
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 9214 5012 9220 5024
rect 9175 4984 9220 5012
rect 9214 4972 9220 4984
rect 9272 4972 9278 5024
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 10134 5012 10140 5024
rect 9732 4984 10140 5012
rect 9732 4972 9738 4984
rect 10134 4972 10140 4984
rect 10192 5012 10198 5024
rect 10229 5015 10287 5021
rect 10229 5012 10241 5015
rect 10192 4984 10241 5012
rect 10192 4972 10198 4984
rect 10229 4981 10241 4984
rect 10275 4981 10287 5015
rect 10229 4975 10287 4981
rect 10321 5015 10379 5021
rect 10321 4981 10333 5015
rect 10367 5012 10379 5015
rect 10410 5012 10416 5024
rect 10367 4984 10416 5012
rect 10367 4981 10379 4984
rect 10321 4975 10379 4981
rect 10410 4972 10416 4984
rect 10468 4972 10474 5024
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 11885 5015 11943 5021
rect 11885 5012 11897 5015
rect 11848 4984 11897 5012
rect 11848 4972 11854 4984
rect 11885 4981 11897 4984
rect 11931 4981 11943 5015
rect 12719 5012 12747 5043
rect 14366 5040 14372 5043
rect 14424 5040 14430 5052
rect 16114 5040 16120 5052
rect 16172 5080 16178 5092
rect 17770 5080 17776 5092
rect 16172 5052 17776 5080
rect 16172 5040 16178 5052
rect 17770 5040 17776 5052
rect 17828 5040 17834 5092
rect 13354 5012 13360 5024
rect 12719 4984 13360 5012
rect 11885 4975 11943 4981
rect 13354 4972 13360 4984
rect 13412 5012 13418 5024
rect 15102 5012 15108 5024
rect 13412 4984 15108 5012
rect 13412 4972 13418 4984
rect 15102 4972 15108 4984
rect 15160 5012 15166 5024
rect 15473 5015 15531 5021
rect 15473 5012 15485 5015
rect 15160 4984 15485 5012
rect 15160 4972 15166 4984
rect 15473 4981 15485 4984
rect 15519 4981 15531 5015
rect 16206 5012 16212 5024
rect 16167 4984 16212 5012
rect 15473 4975 15531 4981
rect 16206 4972 16212 4984
rect 16264 4972 16270 5024
rect 17586 5012 17592 5024
rect 17547 4984 17592 5012
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 18230 5012 18236 5024
rect 18191 4984 18236 5012
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 1104 4922 18860 4944
rect 1104 4870 6912 4922
rect 6964 4870 6976 4922
rect 7028 4870 7040 4922
rect 7092 4870 7104 4922
rect 7156 4870 12843 4922
rect 12895 4870 12907 4922
rect 12959 4870 12971 4922
rect 13023 4870 13035 4922
rect 13087 4870 18860 4922
rect 1104 4848 18860 4870
rect 1504 4780 3096 4808
rect 1504 4681 1532 4780
rect 2308 4743 2366 4749
rect 2308 4709 2320 4743
rect 2354 4740 2366 4743
rect 2406 4740 2412 4752
rect 2354 4712 2412 4740
rect 2354 4709 2366 4712
rect 2308 4703 2366 4709
rect 2406 4700 2412 4712
rect 2464 4740 2470 4752
rect 2774 4740 2780 4752
rect 2464 4712 2780 4740
rect 2464 4700 2470 4712
rect 2774 4700 2780 4712
rect 2832 4700 2838 4752
rect 1489 4675 1547 4681
rect 1489 4641 1501 4675
rect 1535 4641 1547 4675
rect 1489 4635 1547 4641
rect 2038 4604 2044 4616
rect 1999 4576 2044 4604
rect 2038 4564 2044 4576
rect 2096 4564 2102 4616
rect 3068 4536 3096 4780
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 4798 4808 4804 4820
rect 4120 4780 4804 4808
rect 4120 4768 4126 4780
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 6089 4811 6147 4817
rect 6089 4777 6101 4811
rect 6135 4808 6147 4811
rect 7282 4808 7288 4820
rect 6135 4780 7288 4808
rect 6135 4777 6147 4780
rect 6089 4771 6147 4777
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 8294 4768 8300 4820
rect 8352 4808 8358 4820
rect 8846 4808 8852 4820
rect 8352 4780 8852 4808
rect 8352 4768 8358 4780
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 9217 4811 9275 4817
rect 9217 4777 9229 4811
rect 9263 4808 9275 4811
rect 9306 4808 9312 4820
rect 9263 4780 9312 4808
rect 9263 4777 9275 4780
rect 9217 4771 9275 4777
rect 9306 4768 9312 4780
rect 9364 4768 9370 4820
rect 11790 4808 11796 4820
rect 11751 4780 11796 4808
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 11885 4811 11943 4817
rect 11885 4777 11897 4811
rect 11931 4808 11943 4811
rect 12342 4808 12348 4820
rect 11931 4780 12348 4808
rect 11931 4777 11943 4780
rect 11885 4771 11943 4777
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 13173 4811 13231 4817
rect 13173 4777 13185 4811
rect 13219 4808 13231 4811
rect 13725 4811 13783 4817
rect 13725 4808 13737 4811
rect 13219 4780 13737 4808
rect 13219 4777 13231 4780
rect 13173 4771 13231 4777
rect 13725 4777 13737 4780
rect 13771 4777 13783 4811
rect 13725 4771 13783 4777
rect 14093 4811 14151 4817
rect 14093 4777 14105 4811
rect 14139 4808 14151 4811
rect 14458 4808 14464 4820
rect 14139 4780 14464 4808
rect 14139 4777 14151 4780
rect 14093 4771 14151 4777
rect 14458 4768 14464 4780
rect 14516 4808 14522 4820
rect 14918 4808 14924 4820
rect 14516 4780 14924 4808
rect 14516 4768 14522 4780
rect 14918 4768 14924 4780
rect 14976 4768 14982 4820
rect 15289 4811 15347 4817
rect 15289 4777 15301 4811
rect 15335 4777 15347 4811
rect 15654 4808 15660 4820
rect 15615 4780 15660 4808
rect 15289 4771 15347 4777
rect 3142 4700 3148 4752
rect 3200 4740 3206 4752
rect 6362 4740 6368 4752
rect 3200 4712 6368 4740
rect 3200 4700 3206 4712
rect 6362 4700 6368 4712
rect 6420 4700 6426 4752
rect 6549 4743 6607 4749
rect 6549 4709 6561 4743
rect 6595 4740 6607 4743
rect 10318 4740 10324 4752
rect 6595 4712 9720 4740
rect 6595 4709 6607 4712
rect 6549 4703 6607 4709
rect 3786 4632 3792 4684
rect 3844 4672 3850 4684
rect 4062 4672 4068 4684
rect 3844 4644 4068 4672
rect 3844 4632 3850 4644
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 4338 4681 4344 4684
rect 4332 4672 4344 4681
rect 4251 4644 4344 4672
rect 4332 4635 4344 4644
rect 4396 4672 4402 4684
rect 4396 4644 5304 4672
rect 4338 4632 4344 4635
rect 4396 4632 4402 4644
rect 3326 4564 3332 4616
rect 3384 4604 3390 4616
rect 3602 4604 3608 4616
rect 3384 4576 3608 4604
rect 3384 4564 3390 4576
rect 3602 4564 3608 4576
rect 3660 4564 3666 4616
rect 5276 4604 5304 4644
rect 6178 4632 6184 4684
rect 6236 4672 6242 4684
rect 6236 4644 6281 4672
rect 6236 4632 6242 4644
rect 6638 4632 6644 4684
rect 6696 4672 6702 4684
rect 7101 4675 7159 4681
rect 7101 4672 7113 4675
rect 6696 4644 7113 4672
rect 6696 4632 6702 4644
rect 7101 4641 7113 4644
rect 7147 4641 7159 4675
rect 7101 4635 7159 4641
rect 7193 4675 7251 4681
rect 7193 4641 7205 4675
rect 7239 4672 7251 4675
rect 7466 4672 7472 4684
rect 7239 4644 7472 4672
rect 7239 4641 7251 4644
rect 7193 4635 7251 4641
rect 7466 4632 7472 4644
rect 7524 4672 7530 4684
rect 7650 4672 7656 4684
rect 7524 4644 7656 4672
rect 7524 4632 7530 4644
rect 7650 4632 7656 4644
rect 7708 4632 7714 4684
rect 8104 4675 8162 4681
rect 8104 4641 8116 4675
rect 8150 4672 8162 4675
rect 8662 4672 8668 4684
rect 8150 4644 8668 4672
rect 8150 4641 8162 4644
rect 8104 4635 8162 4641
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 6273 4607 6331 4613
rect 6273 4604 6285 4607
rect 5276 4576 6285 4604
rect 6273 4573 6285 4576
rect 6319 4573 6331 4607
rect 7285 4607 7343 4613
rect 7285 4604 7297 4607
rect 6273 4567 6331 4573
rect 6472 4576 7297 4604
rect 3068 4508 4108 4536
rect 1670 4468 1676 4480
rect 1631 4440 1676 4468
rect 1670 4428 1676 4440
rect 1728 4428 1734 4480
rect 3421 4471 3479 4477
rect 3421 4437 3433 4471
rect 3467 4468 3479 4471
rect 3694 4468 3700 4480
rect 3467 4440 3700 4468
rect 3467 4437 3479 4440
rect 3421 4431 3479 4437
rect 3694 4428 3700 4440
rect 3752 4428 3758 4480
rect 4080 4468 4108 4508
rect 5276 4508 6040 4536
rect 5276 4468 5304 4508
rect 5442 4468 5448 4480
rect 4080 4440 5304 4468
rect 5403 4440 5448 4468
rect 5442 4428 5448 4440
rect 5500 4428 5506 4480
rect 5718 4468 5724 4480
rect 5679 4440 5724 4468
rect 5718 4428 5724 4440
rect 5776 4428 5782 4480
rect 6012 4468 6040 4508
rect 6086 4496 6092 4548
rect 6144 4536 6150 4548
rect 6288 4536 6316 4567
rect 6472 4536 6500 4576
rect 7285 4573 7297 4576
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 7742 4564 7748 4616
rect 7800 4604 7806 4616
rect 7837 4607 7895 4613
rect 7837 4604 7849 4607
rect 7800 4576 7849 4604
rect 7800 4564 7806 4576
rect 7837 4573 7849 4576
rect 7883 4573 7895 4607
rect 9692 4604 9720 4712
rect 9784 4712 10324 4740
rect 9784 4681 9812 4712
rect 10318 4700 10324 4712
rect 10376 4700 10382 4752
rect 11054 4740 11060 4752
rect 10704 4712 11060 4740
rect 9769 4675 9827 4681
rect 9769 4641 9781 4675
rect 9815 4641 9827 4675
rect 9769 4635 9827 4641
rect 9858 4632 9864 4684
rect 9916 4632 9922 4684
rect 10036 4675 10094 4681
rect 10036 4641 10048 4675
rect 10082 4672 10094 4675
rect 10704 4672 10732 4712
rect 11054 4700 11060 4712
rect 11112 4740 11118 4752
rect 11330 4740 11336 4752
rect 11112 4712 11336 4740
rect 11112 4700 11118 4712
rect 11330 4700 11336 4712
rect 11388 4700 11394 4752
rect 13081 4743 13139 4749
rect 13081 4709 13093 4743
rect 13127 4740 13139 4743
rect 15304 4740 15332 4771
rect 15654 4768 15660 4780
rect 15712 4768 15718 4820
rect 16574 4740 16580 4752
rect 13127 4712 15332 4740
rect 15396 4712 16580 4740
rect 13127 4709 13139 4712
rect 13081 4703 13139 4709
rect 15396 4672 15424 4712
rect 16574 4700 16580 4712
rect 16632 4700 16638 4752
rect 17310 4672 17316 4684
rect 10082 4644 10732 4672
rect 10796 4644 15424 4672
rect 17271 4644 17316 4672
rect 10082 4641 10094 4644
rect 10036 4635 10094 4641
rect 9876 4604 9904 4632
rect 9692 4576 9904 4604
rect 7837 4567 7895 4573
rect 6144 4508 6500 4536
rect 6144 4496 6150 4508
rect 8846 4496 8852 4548
rect 8904 4536 8910 4548
rect 8904 4508 9812 4536
rect 8904 4496 8910 4508
rect 6549 4471 6607 4477
rect 6549 4468 6561 4471
rect 6012 4440 6561 4468
rect 6549 4437 6561 4440
rect 6595 4437 6607 4471
rect 6730 4468 6736 4480
rect 6691 4440 6736 4468
rect 6549 4431 6607 4437
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 6822 4428 6828 4480
rect 6880 4468 6886 4480
rect 9674 4468 9680 4480
rect 6880 4440 9680 4468
rect 6880 4428 6886 4440
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 9784 4468 9812 4508
rect 10796 4468 10824 4644
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 17865 4675 17923 4681
rect 17865 4641 17877 4675
rect 17911 4641 17923 4675
rect 17865 4635 17923 4641
rect 11330 4564 11336 4616
rect 11388 4604 11394 4616
rect 11977 4607 12035 4613
rect 11977 4604 11989 4607
rect 11388 4576 11989 4604
rect 11388 4564 11394 4576
rect 11977 4573 11989 4576
rect 12023 4573 12035 4607
rect 11977 4567 12035 4573
rect 12526 4564 12532 4616
rect 12584 4564 12590 4616
rect 13354 4604 13360 4616
rect 13315 4576 13360 4604
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 14182 4604 14188 4616
rect 14143 4576 14188 4604
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14366 4604 14372 4616
rect 14279 4576 14372 4604
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 15194 4564 15200 4616
rect 15252 4604 15258 4616
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 15252 4576 15761 4604
rect 15252 4564 15258 4576
rect 15749 4573 15761 4576
rect 15795 4573 15807 4607
rect 15930 4604 15936 4616
rect 15891 4576 15936 4604
rect 15749 4567 15807 4573
rect 15930 4564 15936 4576
rect 15988 4564 15994 4616
rect 17880 4604 17908 4635
rect 16040 4576 17908 4604
rect 11606 4496 11612 4548
rect 11664 4536 11670 4548
rect 12544 4536 12572 4564
rect 13170 4536 13176 4548
rect 11664 4508 13176 4536
rect 11664 4496 11670 4508
rect 13170 4496 13176 4508
rect 13228 4496 13234 4548
rect 14384 4536 14412 4564
rect 15010 4536 15016 4548
rect 14384 4508 15016 4536
rect 15010 4496 15016 4508
rect 15068 4536 15074 4548
rect 15948 4536 15976 4564
rect 15068 4508 15976 4536
rect 15068 4496 15074 4508
rect 11146 4468 11152 4480
rect 9784 4440 10824 4468
rect 11107 4440 11152 4468
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 11425 4471 11483 4477
rect 11425 4437 11437 4471
rect 11471 4468 11483 4471
rect 12526 4468 12532 4480
rect 11471 4440 12532 4468
rect 11471 4437 11483 4440
rect 11425 4431 11483 4437
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 12710 4468 12716 4480
rect 12671 4440 12716 4468
rect 12710 4428 12716 4440
rect 12768 4428 12774 4480
rect 12802 4428 12808 4480
rect 12860 4468 12866 4480
rect 16040 4468 16068 4576
rect 17494 4468 17500 4480
rect 12860 4440 16068 4468
rect 17455 4440 17500 4468
rect 12860 4428 12866 4440
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 17862 4428 17868 4480
rect 17920 4468 17926 4480
rect 18049 4471 18107 4477
rect 18049 4468 18061 4471
rect 17920 4440 18061 4468
rect 17920 4428 17926 4440
rect 18049 4437 18061 4440
rect 18095 4437 18107 4471
rect 18049 4431 18107 4437
rect 1104 4378 18860 4400
rect 1104 4326 3947 4378
rect 3999 4326 4011 4378
rect 4063 4326 4075 4378
rect 4127 4326 4139 4378
rect 4191 4326 9878 4378
rect 9930 4326 9942 4378
rect 9994 4326 10006 4378
rect 10058 4326 10070 4378
rect 10122 4326 15808 4378
rect 15860 4326 15872 4378
rect 15924 4326 15936 4378
rect 15988 4326 16000 4378
rect 16052 4326 18860 4378
rect 1104 4304 18860 4326
rect 2038 4224 2044 4276
rect 2096 4264 2102 4276
rect 3786 4264 3792 4276
rect 2096 4236 3792 4264
rect 2096 4224 2102 4236
rect 2406 4196 2412 4208
rect 2332 4168 2412 4196
rect 2332 4137 2360 4168
rect 2406 4156 2412 4168
rect 2464 4156 2470 4208
rect 2700 4137 2728 4236
rect 3786 4224 3792 4236
rect 3844 4224 3850 4276
rect 4065 4267 4123 4273
rect 4065 4233 4077 4267
rect 4111 4264 4123 4267
rect 4338 4264 4344 4276
rect 4111 4236 4344 4264
rect 4111 4233 4123 4236
rect 4065 4227 4123 4233
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 11606 4264 11612 4276
rect 4488 4236 11612 4264
rect 4488 4224 4494 4236
rect 11606 4224 11612 4236
rect 11664 4224 11670 4276
rect 13170 4224 13176 4276
rect 13228 4264 13234 4276
rect 15010 4264 15016 4276
rect 13228 4236 14872 4264
rect 14971 4236 15016 4264
rect 13228 4224 13234 4236
rect 7466 4156 7472 4208
rect 7524 4196 7530 4208
rect 8202 4196 8208 4208
rect 7524 4168 8208 4196
rect 7524 4156 7530 4168
rect 8202 4156 8208 4168
rect 8260 4156 8266 4208
rect 9306 4196 9312 4208
rect 9232 4168 9312 4196
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4097 2375 4131
rect 2317 4091 2375 4097
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4097 2743 4131
rect 5166 4128 5172 4140
rect 2685 4091 2743 4097
rect 4264 4100 5172 4128
rect 2041 4063 2099 4069
rect 2041 4029 2053 4063
rect 2087 4060 2099 4063
rect 4264 4060 4292 4100
rect 5166 4088 5172 4100
rect 5224 4088 5230 4140
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 5537 4131 5595 4137
rect 5537 4128 5549 4131
rect 5500 4100 5549 4128
rect 5500 4088 5506 4100
rect 5537 4097 5549 4100
rect 5583 4097 5595 4131
rect 5537 4091 5595 4097
rect 5736 4100 7512 4128
rect 2087 4032 4292 4060
rect 4341 4063 4399 4069
rect 2087 4029 2099 4032
rect 2041 4023 2099 4029
rect 4341 4029 4353 4063
rect 4387 4060 4399 4063
rect 4890 4060 4896 4072
rect 4387 4032 4896 4060
rect 4387 4029 4399 4032
rect 4341 4023 4399 4029
rect 4890 4020 4896 4032
rect 4948 4020 4954 4072
rect 5353 4063 5411 4069
rect 5353 4029 5365 4063
rect 5399 4060 5411 4063
rect 5626 4060 5632 4072
rect 5399 4032 5632 4060
rect 5399 4029 5411 4032
rect 5353 4023 5411 4029
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 2952 3995 3010 4001
rect 2952 3961 2964 3995
rect 2998 3992 3010 3995
rect 3694 3992 3700 4004
rect 2998 3964 3700 3992
rect 2998 3961 3010 3964
rect 2952 3955 3010 3961
rect 3694 3952 3700 3964
rect 3752 3952 3758 4004
rect 3786 3952 3792 4004
rect 3844 3992 3850 4004
rect 3844 3964 4568 3992
rect 3844 3952 3850 3964
rect 1673 3927 1731 3933
rect 1673 3893 1685 3927
rect 1719 3924 1731 3927
rect 1946 3924 1952 3936
rect 1719 3896 1952 3924
rect 1719 3893 1731 3896
rect 1673 3887 1731 3893
rect 1946 3884 1952 3896
rect 2004 3884 2010 3936
rect 2133 3927 2191 3933
rect 2133 3893 2145 3927
rect 2179 3924 2191 3927
rect 4246 3924 4252 3936
rect 2179 3896 4252 3924
rect 2179 3893 2191 3896
rect 2133 3887 2191 3893
rect 4246 3884 4252 3896
rect 4304 3884 4310 3936
rect 4540 3933 4568 3964
rect 5166 3952 5172 4004
rect 5224 3992 5230 4004
rect 5736 3992 5764 4100
rect 5994 4060 6000 4072
rect 5955 4032 6000 4060
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 6454 4020 6460 4072
rect 6512 4060 6518 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6512 4032 6837 4060
rect 6512 4020 6518 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 7484 4060 7512 4100
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 8113 4131 8171 4137
rect 8113 4128 8125 4131
rect 7616 4100 8125 4128
rect 7616 4088 7622 4100
rect 8113 4097 8125 4100
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4128 8355 4131
rect 8662 4128 8668 4140
rect 8343 4100 8668 4128
rect 8343 4097 8355 4100
rect 8297 4091 8355 4097
rect 8662 4088 8668 4100
rect 8720 4088 8726 4140
rect 9232 4137 9260 4168
rect 9306 4156 9312 4168
rect 9364 4156 9370 4208
rect 13630 4196 13636 4208
rect 13188 4168 13636 4196
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4097 9275 4131
rect 10226 4128 10232 4140
rect 10187 4100 10232 4128
rect 9217 4091 9275 4097
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 10318 4088 10324 4140
rect 10376 4128 10382 4140
rect 10689 4131 10747 4137
rect 10689 4128 10701 4131
rect 10376 4100 10701 4128
rect 10376 4088 10382 4100
rect 10689 4097 10701 4100
rect 10735 4097 10747 4131
rect 10689 4091 10747 4097
rect 12710 4088 12716 4140
rect 12768 4128 12774 4140
rect 13188 4137 13216 4168
rect 13630 4156 13636 4168
rect 13688 4156 13694 4208
rect 14844 4196 14872 4236
rect 15010 4224 15016 4236
rect 15068 4224 15074 4276
rect 16206 4264 16212 4276
rect 15580 4236 16212 4264
rect 15580 4196 15608 4236
rect 16206 4224 16212 4236
rect 16264 4224 16270 4276
rect 14844 4168 15608 4196
rect 15654 4156 15660 4208
rect 15712 4196 15718 4208
rect 15712 4168 17448 4196
rect 15712 4156 15718 4168
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12768 4100 13001 4128
rect 12768 4088 12774 4100
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 13173 4131 13231 4137
rect 13173 4097 13185 4131
rect 13219 4097 13231 4131
rect 13173 4091 13231 4097
rect 15194 4088 15200 4140
rect 15252 4128 15258 4140
rect 15562 4128 15568 4140
rect 15252 4100 15568 4128
rect 15252 4088 15258 4100
rect 15562 4088 15568 4100
rect 15620 4088 15626 4140
rect 7650 4060 7656 4072
rect 7484 4032 7656 4060
rect 6825 4023 6883 4029
rect 7650 4020 7656 4032
rect 7708 4020 7714 4072
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 8021 4063 8079 4069
rect 8021 4060 8033 4063
rect 7984 4032 8033 4060
rect 7984 4020 7990 4032
rect 8021 4029 8033 4032
rect 8067 4029 8079 4063
rect 8021 4023 8079 4029
rect 10137 4063 10195 4069
rect 10137 4029 10149 4063
rect 10183 4060 10195 4063
rect 10594 4060 10600 4072
rect 10183 4032 10600 4060
rect 10183 4029 10195 4032
rect 10137 4023 10195 4029
rect 10594 4020 10600 4032
rect 10652 4020 10658 4072
rect 13446 4020 13452 4072
rect 13504 4060 13510 4072
rect 13633 4063 13691 4069
rect 13633 4060 13645 4063
rect 13504 4032 13645 4060
rect 13504 4020 13510 4032
rect 13633 4029 13645 4032
rect 13679 4029 13691 4063
rect 16298 4060 16304 4072
rect 13633 4023 13691 4029
rect 13740 4032 16304 4060
rect 5224 3964 5764 3992
rect 5224 3952 5230 3964
rect 5810 3952 5816 4004
rect 5868 3992 5874 4004
rect 6273 3995 6331 4001
rect 6273 3992 6285 3995
rect 5868 3964 6285 3992
rect 5868 3952 5874 3964
rect 6273 3961 6285 3964
rect 6319 3961 6331 3995
rect 6273 3955 6331 3961
rect 6546 3952 6552 4004
rect 6604 3992 6610 4004
rect 7101 3995 7159 4001
rect 7101 3992 7113 3995
rect 6604 3964 7113 3992
rect 6604 3952 6610 3964
rect 7101 3961 7113 3964
rect 7147 3961 7159 3995
rect 9033 3995 9091 4001
rect 9033 3992 9045 3995
rect 7101 3955 7159 3961
rect 7668 3964 9045 3992
rect 4525 3927 4583 3933
rect 4525 3893 4537 3927
rect 4571 3893 4583 3927
rect 4525 3887 4583 3893
rect 4890 3884 4896 3936
rect 4948 3924 4954 3936
rect 4985 3927 5043 3933
rect 4985 3924 4997 3927
rect 4948 3896 4997 3924
rect 4948 3884 4954 3896
rect 4985 3893 4997 3896
rect 5031 3893 5043 3927
rect 4985 3887 5043 3893
rect 5445 3927 5503 3933
rect 5445 3893 5457 3927
rect 5491 3924 5503 3927
rect 6730 3924 6736 3936
rect 5491 3896 6736 3924
rect 5491 3893 5503 3896
rect 5445 3887 5503 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 7668 3933 7696 3964
rect 9033 3961 9045 3964
rect 9079 3961 9091 3995
rect 9033 3955 9091 3961
rect 10045 3995 10103 4001
rect 10045 3961 10057 3995
rect 10091 3992 10103 3995
rect 10956 3995 11014 4001
rect 10091 3964 10916 3992
rect 10091 3961 10103 3964
rect 10045 3955 10103 3961
rect 7653 3927 7711 3933
rect 7653 3893 7665 3927
rect 7699 3893 7711 3927
rect 7653 3887 7711 3893
rect 8570 3884 8576 3936
rect 8628 3924 8634 3936
rect 8665 3927 8723 3933
rect 8665 3924 8677 3927
rect 8628 3896 8677 3924
rect 8628 3884 8634 3896
rect 8665 3893 8677 3896
rect 8711 3893 8723 3927
rect 8665 3887 8723 3893
rect 8754 3884 8760 3936
rect 8812 3924 8818 3936
rect 9125 3927 9183 3933
rect 9125 3924 9137 3927
rect 8812 3896 9137 3924
rect 8812 3884 8818 3896
rect 9125 3893 9137 3896
rect 9171 3893 9183 3927
rect 9125 3887 9183 3893
rect 9490 3884 9496 3936
rect 9548 3924 9554 3936
rect 9677 3927 9735 3933
rect 9677 3924 9689 3927
rect 9548 3896 9689 3924
rect 9548 3884 9554 3896
rect 9677 3893 9689 3896
rect 9723 3893 9735 3927
rect 10888 3924 10916 3964
rect 10956 3961 10968 3995
rect 11002 3992 11014 3995
rect 11146 3992 11152 4004
rect 11002 3964 11152 3992
rect 11002 3961 11014 3964
rect 10956 3955 11014 3961
rect 11146 3952 11152 3964
rect 11204 3952 11210 4004
rect 13740 3992 13768 4032
rect 16298 4020 16304 4032
rect 16356 4020 16362 4072
rect 17420 4069 17448 4168
rect 17405 4063 17463 4069
rect 17405 4029 17417 4063
rect 17451 4029 17463 4063
rect 17405 4023 17463 4029
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 13906 4001 13912 4004
rect 13900 3992 13912 4001
rect 11256 3964 13768 3992
rect 13867 3964 13912 3992
rect 11256 3924 11284 3964
rect 13900 3955 13912 3964
rect 13906 3952 13912 3955
rect 13964 3952 13970 4004
rect 14826 3952 14832 4004
rect 14884 3992 14890 4004
rect 18064 3992 18092 4023
rect 14884 3964 18092 3992
rect 14884 3952 14890 3964
rect 12066 3924 12072 3936
rect 10888 3896 11284 3924
rect 12027 3896 12072 3924
rect 9677 3887 9735 3893
rect 12066 3884 12072 3896
rect 12124 3884 12130 3936
rect 12529 3927 12587 3933
rect 12529 3893 12541 3927
rect 12575 3924 12587 3927
rect 12710 3924 12716 3936
rect 12575 3896 12716 3924
rect 12575 3893 12587 3896
rect 12529 3887 12587 3893
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 12897 3927 12955 3933
rect 12897 3893 12909 3927
rect 12943 3924 12955 3927
rect 14550 3924 14556 3936
rect 12943 3896 14556 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 16666 3884 16672 3936
rect 16724 3924 16730 3936
rect 17402 3924 17408 3936
rect 16724 3896 17408 3924
rect 16724 3884 16730 3896
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 17586 3924 17592 3936
rect 17547 3896 17592 3924
rect 17586 3884 17592 3896
rect 17644 3884 17650 3936
rect 18233 3927 18291 3933
rect 18233 3893 18245 3927
rect 18279 3924 18291 3927
rect 18322 3924 18328 3936
rect 18279 3896 18328 3924
rect 18279 3893 18291 3896
rect 18233 3887 18291 3893
rect 18322 3884 18328 3896
rect 18380 3884 18386 3936
rect 1104 3834 18860 3856
rect 1104 3782 6912 3834
rect 6964 3782 6976 3834
rect 7028 3782 7040 3834
rect 7092 3782 7104 3834
rect 7156 3782 12843 3834
rect 12895 3782 12907 3834
rect 12959 3782 12971 3834
rect 13023 3782 13035 3834
rect 13087 3782 18860 3834
rect 1104 3760 18860 3782
rect 2501 3723 2559 3729
rect 2501 3689 2513 3723
rect 2547 3720 2559 3723
rect 2774 3720 2780 3732
rect 2547 3692 2780 3720
rect 2547 3689 2559 3692
rect 2501 3683 2559 3689
rect 2774 3680 2780 3692
rect 2832 3680 2838 3732
rect 2961 3723 3019 3729
rect 2961 3689 2973 3723
rect 3007 3720 3019 3723
rect 4893 3723 4951 3729
rect 4893 3720 4905 3723
rect 3007 3692 4905 3720
rect 3007 3689 3019 3692
rect 2961 3683 3019 3689
rect 4893 3689 4905 3692
rect 4939 3689 4951 3723
rect 4893 3683 4951 3689
rect 4982 3680 4988 3732
rect 5040 3720 5046 3732
rect 8386 3720 8392 3732
rect 5040 3692 8392 3720
rect 5040 3680 5046 3692
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 10318 3680 10324 3732
rect 10376 3720 10382 3732
rect 13909 3723 13967 3729
rect 10376 3692 11652 3720
rect 10376 3680 10382 3692
rect 5166 3652 5172 3664
rect 2332 3624 5172 3652
rect 1578 3584 1584 3596
rect 1539 3556 1584 3584
rect 1578 3544 1584 3556
rect 1636 3544 1642 3596
rect 2332 3593 2360 3624
rect 5166 3612 5172 3624
rect 5224 3612 5230 3664
rect 5261 3655 5319 3661
rect 5261 3621 5273 3655
rect 5307 3652 5319 3655
rect 5442 3652 5448 3664
rect 5307 3624 5448 3652
rect 5307 3621 5319 3624
rect 5261 3615 5319 3621
rect 5442 3612 5448 3624
rect 5500 3652 5506 3664
rect 5690 3655 5748 3661
rect 5690 3652 5702 3655
rect 5500 3624 5702 3652
rect 5500 3612 5506 3624
rect 5690 3621 5702 3624
rect 5736 3621 5748 3655
rect 5690 3615 5748 3621
rect 10045 3655 10103 3661
rect 10045 3621 10057 3655
rect 10091 3652 10103 3655
rect 10410 3652 10416 3664
rect 10091 3624 10416 3652
rect 10091 3621 10103 3624
rect 10045 3615 10103 3621
rect 10410 3612 10416 3624
rect 10468 3612 10474 3664
rect 10502 3612 10508 3664
rect 10560 3652 10566 3664
rect 11517 3655 11575 3661
rect 11517 3652 11529 3655
rect 10560 3624 11529 3652
rect 10560 3612 10566 3624
rect 11517 3621 11529 3624
rect 11563 3621 11575 3655
rect 11624 3652 11652 3692
rect 13909 3689 13921 3723
rect 13955 3720 13967 3723
rect 14182 3720 14188 3732
rect 13955 3692 14188 3720
rect 13955 3689 13967 3692
rect 13909 3683 13967 3689
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 14369 3723 14427 3729
rect 14369 3689 14381 3723
rect 14415 3720 14427 3723
rect 17126 3720 17132 3732
rect 14415 3692 17132 3720
rect 14415 3689 14427 3692
rect 14369 3683 14427 3689
rect 17126 3680 17132 3692
rect 17184 3720 17190 3732
rect 17184 3692 17908 3720
rect 17184 3680 17190 3692
rect 12066 3652 12072 3664
rect 11624 3624 12072 3652
rect 11517 3615 11575 3621
rect 12066 3612 12072 3624
rect 12124 3652 12130 3664
rect 12498 3655 12556 3661
rect 12498 3652 12510 3655
rect 12124 3624 12510 3652
rect 12124 3612 12130 3624
rect 12498 3621 12510 3624
rect 12544 3621 12556 3655
rect 12498 3615 12556 3621
rect 12710 3612 12716 3664
rect 12768 3652 12774 3664
rect 12768 3624 15332 3652
rect 12768 3612 12774 3624
rect 2317 3587 2375 3593
rect 2317 3553 2329 3587
rect 2363 3553 2375 3587
rect 3326 3584 3332 3596
rect 3287 3556 3332 3584
rect 2317 3547 2375 3553
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 4801 3587 4859 3593
rect 4801 3553 4813 3587
rect 4847 3584 4859 3587
rect 5534 3584 5540 3596
rect 4847 3556 5540 3584
rect 4847 3553 4859 3556
rect 4801 3547 4859 3553
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 7357 3587 7415 3593
rect 7357 3584 7369 3587
rect 6840 3556 7369 3584
rect 1210 3476 1216 3528
rect 1268 3516 1274 3528
rect 1765 3519 1823 3525
rect 1765 3516 1777 3519
rect 1268 3488 1777 3516
rect 1268 3476 1274 3488
rect 1765 3485 1777 3488
rect 1811 3485 1823 3519
rect 1765 3479 1823 3485
rect 3142 3476 3148 3528
rect 3200 3516 3206 3528
rect 3421 3519 3479 3525
rect 3421 3516 3433 3519
rect 3200 3488 3433 3516
rect 3200 3476 3206 3488
rect 3421 3485 3433 3488
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 4338 3516 4344 3528
rect 3651 3488 4344 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 5077 3519 5135 3525
rect 5077 3485 5089 3519
rect 5123 3516 5135 3519
rect 5261 3519 5319 3525
rect 5261 3516 5273 3519
rect 5123 3488 5273 3516
rect 5123 3485 5135 3488
rect 5077 3479 5135 3485
rect 5261 3485 5273 3488
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 5445 3519 5503 3525
rect 5445 3485 5457 3519
rect 5491 3485 5503 3519
rect 5445 3479 5503 3485
rect 4798 3408 4804 3460
rect 4856 3448 4862 3460
rect 5460 3448 5488 3479
rect 4856 3420 5488 3448
rect 4856 3408 4862 3420
rect 4433 3383 4491 3389
rect 4433 3349 4445 3383
rect 4479 3380 4491 3383
rect 4982 3380 4988 3392
rect 4479 3352 4988 3380
rect 4479 3349 4491 3352
rect 4433 3343 4491 3349
rect 4982 3340 4988 3352
rect 5040 3340 5046 3392
rect 5166 3340 5172 3392
rect 5224 3380 5230 3392
rect 6840 3389 6868 3556
rect 7357 3553 7369 3556
rect 7403 3553 7415 3587
rect 7357 3547 7415 3553
rect 8757 3587 8815 3593
rect 8757 3553 8769 3587
rect 8803 3584 8815 3587
rect 9122 3584 9128 3596
rect 8803 3556 9128 3584
rect 8803 3553 8815 3556
rect 8757 3547 8815 3553
rect 9122 3544 9128 3556
rect 9180 3544 9186 3596
rect 10137 3587 10195 3593
rect 10137 3553 10149 3587
rect 10183 3584 10195 3587
rect 10778 3584 10784 3596
rect 10183 3556 10784 3584
rect 10183 3553 10195 3556
rect 10137 3547 10195 3553
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3584 11115 3587
rect 11701 3587 11759 3593
rect 11701 3584 11713 3587
rect 11103 3556 11713 3584
rect 11103 3553 11115 3556
rect 11057 3547 11115 3553
rect 11701 3553 11713 3556
rect 11747 3584 11759 3587
rect 11882 3584 11888 3596
rect 11747 3556 11888 3584
rect 11747 3553 11759 3556
rect 11701 3547 11759 3553
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 12253 3587 12311 3593
rect 12253 3553 12265 3587
rect 12299 3584 12311 3587
rect 12342 3584 12348 3596
rect 12299 3556 12348 3584
rect 12299 3553 12311 3556
rect 12253 3547 12311 3553
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 14090 3544 14096 3596
rect 14148 3584 14154 3596
rect 15304 3593 15332 3624
rect 14277 3587 14335 3593
rect 14277 3584 14289 3587
rect 14148 3556 14289 3584
rect 14148 3544 14154 3556
rect 14277 3553 14289 3556
rect 14323 3553 14335 3587
rect 15289 3587 15347 3593
rect 14277 3547 14335 3553
rect 14384 3556 14596 3584
rect 7101 3519 7159 3525
rect 7101 3485 7113 3519
rect 7147 3485 7159 3519
rect 7101 3479 7159 3485
rect 6825 3383 6883 3389
rect 6825 3380 6837 3383
rect 5224 3352 6837 3380
rect 5224 3340 5230 3352
rect 6825 3349 6837 3352
rect 6871 3349 6883 3383
rect 7116 3380 7144 3479
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8536 3488 8953 3516
rect 8536 3476 8542 3488
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 10226 3516 10232 3528
rect 10187 3488 10232 3516
rect 8941 3479 8999 3485
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10410 3476 10416 3528
rect 10468 3516 10474 3528
rect 10870 3516 10876 3528
rect 10468 3488 10876 3516
rect 10468 3476 10474 3488
rect 10870 3476 10876 3488
rect 10928 3476 10934 3528
rect 11149 3519 11207 3525
rect 11149 3485 11161 3519
rect 11195 3485 11207 3519
rect 11149 3479 11207 3485
rect 9766 3408 9772 3460
rect 9824 3448 9830 3460
rect 11164 3448 11192 3479
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 11333 3519 11391 3525
rect 11333 3516 11345 3519
rect 11296 3488 11345 3516
rect 11296 3476 11302 3488
rect 11333 3485 11345 3488
rect 11379 3485 11391 3519
rect 11333 3479 11391 3485
rect 11517 3519 11575 3525
rect 11517 3485 11529 3519
rect 11563 3516 11575 3519
rect 12161 3519 12219 3525
rect 12161 3516 12173 3519
rect 11563 3488 12173 3516
rect 11563 3485 11575 3488
rect 11517 3479 11575 3485
rect 12161 3485 12173 3488
rect 12207 3485 12219 3519
rect 12161 3479 12219 3485
rect 13262 3476 13268 3528
rect 13320 3516 13326 3528
rect 14384 3516 14412 3556
rect 13320 3488 14412 3516
rect 14461 3519 14519 3525
rect 13320 3476 13326 3488
rect 14461 3485 14473 3519
rect 14507 3485 14519 3519
rect 14568 3516 14596 3556
rect 15289 3553 15301 3587
rect 15335 3553 15347 3587
rect 15562 3584 15568 3596
rect 15289 3547 15347 3553
rect 15396 3556 15568 3584
rect 15396 3516 15424 3556
rect 15562 3544 15568 3556
rect 15620 3544 15626 3596
rect 16574 3544 16580 3596
rect 16632 3584 16638 3596
rect 17880 3593 17908 3692
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 16632 3556 17325 3584
rect 16632 3544 16638 3556
rect 17313 3553 17325 3556
rect 17359 3553 17371 3587
rect 17313 3547 17371 3553
rect 17865 3587 17923 3593
rect 17865 3553 17877 3587
rect 17911 3553 17923 3587
rect 17865 3547 17923 3553
rect 14568 3488 15424 3516
rect 15473 3519 15531 3525
rect 14461 3479 14519 3485
rect 15473 3485 15485 3519
rect 15519 3485 15531 3519
rect 15473 3479 15531 3485
rect 12250 3448 12256 3460
rect 9824 3420 10824 3448
rect 11164 3420 12256 3448
rect 9824 3408 9830 3420
rect 7742 3380 7748 3392
rect 7116 3352 7748 3380
rect 6825 3343 6883 3349
rect 7742 3340 7748 3352
rect 7800 3340 7806 3392
rect 8481 3383 8539 3389
rect 8481 3349 8493 3383
rect 8527 3380 8539 3383
rect 8662 3380 8668 3392
rect 8527 3352 8668 3380
rect 8527 3349 8539 3352
rect 8481 3343 8539 3349
rect 8662 3340 8668 3352
rect 8720 3340 8726 3392
rect 9582 3340 9588 3392
rect 9640 3380 9646 3392
rect 9677 3383 9735 3389
rect 9677 3380 9689 3383
rect 9640 3352 9689 3380
rect 9640 3340 9646 3352
rect 9677 3349 9689 3352
rect 9723 3349 9735 3383
rect 9677 3343 9735 3349
rect 10594 3340 10600 3392
rect 10652 3380 10658 3392
rect 10689 3383 10747 3389
rect 10689 3380 10701 3383
rect 10652 3352 10701 3380
rect 10652 3340 10658 3352
rect 10689 3349 10701 3352
rect 10735 3349 10747 3383
rect 10796 3380 10824 3420
rect 12250 3408 12256 3420
rect 12308 3408 12314 3460
rect 13633 3451 13691 3457
rect 13633 3417 13645 3451
rect 13679 3448 13691 3451
rect 13906 3448 13912 3460
rect 13679 3420 13912 3448
rect 13679 3417 13691 3420
rect 13633 3411 13691 3417
rect 13906 3408 13912 3420
rect 13964 3448 13970 3460
rect 14476 3448 14504 3479
rect 13964 3420 14504 3448
rect 13964 3408 13970 3420
rect 11790 3380 11796 3392
rect 10796 3352 11796 3380
rect 10689 3343 10747 3349
rect 11790 3340 11796 3352
rect 11848 3340 11854 3392
rect 11885 3383 11943 3389
rect 11885 3349 11897 3383
rect 11931 3380 11943 3383
rect 12066 3380 12072 3392
rect 11931 3352 12072 3380
rect 11931 3349 11943 3352
rect 11885 3343 11943 3349
rect 12066 3340 12072 3352
rect 12124 3340 12130 3392
rect 12161 3383 12219 3389
rect 12161 3349 12173 3383
rect 12207 3380 12219 3383
rect 15488 3380 15516 3479
rect 17494 3380 17500 3392
rect 12207 3352 15516 3380
rect 17455 3352 17500 3380
rect 12207 3349 12219 3352
rect 12161 3343 12219 3349
rect 17494 3340 17500 3352
rect 17552 3340 17558 3392
rect 18046 3380 18052 3392
rect 18007 3352 18052 3380
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 1104 3290 18860 3312
rect 1104 3238 3947 3290
rect 3999 3238 4011 3290
rect 4063 3238 4075 3290
rect 4127 3238 4139 3290
rect 4191 3238 9878 3290
rect 9930 3238 9942 3290
rect 9994 3238 10006 3290
rect 10058 3238 10070 3290
rect 10122 3238 15808 3290
rect 15860 3238 15872 3290
rect 15924 3238 15936 3290
rect 15988 3238 16000 3290
rect 16052 3238 18860 3290
rect 1104 3216 18860 3238
rect 3142 3176 3148 3188
rect 3103 3148 3148 3176
rect 3142 3136 3148 3148
rect 3200 3136 3206 3188
rect 5534 3176 5540 3188
rect 5495 3148 5540 3176
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 8113 3179 8171 3185
rect 8113 3145 8125 3179
rect 8159 3176 8171 3179
rect 8754 3176 8760 3188
rect 8159 3148 8760 3176
rect 8159 3145 8171 3148
rect 8113 3139 8171 3145
rect 8754 3136 8760 3148
rect 8812 3136 8818 3188
rect 9122 3176 9128 3188
rect 9083 3148 9128 3176
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 10137 3179 10195 3185
rect 10137 3145 10149 3179
rect 10183 3176 10195 3179
rect 11698 3176 11704 3188
rect 10183 3148 11704 3176
rect 10183 3145 10195 3148
rect 10137 3139 10195 3145
rect 11698 3136 11704 3148
rect 11756 3136 11762 3188
rect 11790 3136 11796 3188
rect 11848 3176 11854 3188
rect 15381 3179 15439 3185
rect 15381 3176 15393 3179
rect 11848 3148 15393 3176
rect 11848 3136 11854 3148
rect 15381 3145 15393 3148
rect 15427 3145 15439 3179
rect 15381 3139 15439 3145
rect 15470 3136 15476 3188
rect 15528 3176 15534 3188
rect 16390 3176 16396 3188
rect 15528 3148 16396 3176
rect 15528 3136 15534 3148
rect 16390 3136 16396 3148
rect 16448 3176 16454 3188
rect 16448 3148 18092 3176
rect 16448 3136 16454 3148
rect 4525 3111 4583 3117
rect 4525 3077 4537 3111
rect 4571 3108 4583 3111
rect 5442 3108 5448 3120
rect 4571 3080 5448 3108
rect 4571 3077 4583 3080
rect 4525 3071 4583 3077
rect 5442 3068 5448 3080
rect 5500 3068 5506 3120
rect 5902 3068 5908 3120
rect 5960 3108 5966 3120
rect 9030 3108 9036 3120
rect 5960 3080 9036 3108
rect 5960 3068 5966 3080
rect 9030 3068 9036 3080
rect 9088 3068 9094 3120
rect 9398 3068 9404 3120
rect 9456 3108 9462 3120
rect 9456 3080 9720 3108
rect 9456 3068 9462 3080
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 2774 3040 2780 3052
rect 1903 3012 2780 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 3694 3040 3700 3052
rect 3655 3012 3700 3040
rect 3694 3000 3700 3012
rect 3752 3000 3758 3052
rect 4982 3040 4988 3052
rect 4943 3012 4988 3040
rect 4982 3000 4988 3012
rect 5040 3000 5046 3052
rect 5166 3040 5172 3052
rect 5127 3012 5172 3040
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 6086 3040 6092 3052
rect 6047 3012 6092 3040
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 8662 3040 8668 3052
rect 8623 3012 8668 3040
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 9582 3040 9588 3052
rect 9543 3012 9588 3040
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 9692 3049 9720 3080
rect 11146 3068 11152 3120
rect 11204 3108 11210 3120
rect 11204 3080 11836 3108
rect 11204 3068 11210 3080
rect 9677 3043 9735 3049
rect 9677 3009 9689 3043
rect 9723 3009 9735 3043
rect 10594 3040 10600 3052
rect 10555 3012 10600 3040
rect 9677 3003 9735 3009
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 10781 3043 10839 3049
rect 10781 3009 10793 3043
rect 10827 3040 10839 3043
rect 11054 3040 11060 3052
rect 10827 3012 11060 3040
rect 10827 3009 10839 3012
rect 10781 3003 10839 3009
rect 11054 3000 11060 3012
rect 11112 3000 11118 3052
rect 11606 3040 11612 3052
rect 11567 3012 11612 3040
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3009 11759 3043
rect 11808 3040 11836 3080
rect 11882 3068 11888 3120
rect 11940 3108 11946 3120
rect 12437 3111 12495 3117
rect 12437 3108 12449 3111
rect 11940 3080 12449 3108
rect 11940 3068 11946 3080
rect 12437 3077 12449 3080
rect 12483 3077 12495 3111
rect 12437 3071 12495 3077
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 11808 3012 13001 3040
rect 11701 3003 11759 3009
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 1581 2975 1639 2981
rect 1581 2941 1593 2975
rect 1627 2941 1639 2975
rect 2314 2972 2320 2984
rect 2275 2944 2320 2972
rect 1581 2935 1639 2941
rect 1596 2836 1624 2935
rect 2314 2932 2320 2944
rect 2372 2932 2378 2984
rect 2866 2932 2872 2984
rect 2924 2972 2930 2984
rect 3513 2975 3571 2981
rect 3513 2972 3525 2975
rect 2924 2944 3525 2972
rect 2924 2932 2930 2944
rect 3513 2941 3525 2944
rect 3559 2941 3571 2975
rect 3513 2935 3571 2941
rect 3602 2932 3608 2984
rect 3660 2972 3666 2984
rect 4890 2972 4896 2984
rect 3660 2944 3705 2972
rect 4851 2944 4896 2972
rect 3660 2932 3666 2944
rect 4890 2932 4896 2944
rect 4948 2932 4954 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 5736 2944 6837 2972
rect 2130 2864 2136 2916
rect 2188 2904 2194 2916
rect 2593 2907 2651 2913
rect 2593 2904 2605 2907
rect 2188 2876 2605 2904
rect 2188 2864 2194 2876
rect 2593 2873 2605 2876
rect 2639 2873 2651 2907
rect 2593 2867 2651 2873
rect 5736 2836 5764 2944
rect 6825 2941 6837 2944
rect 6871 2972 6883 2975
rect 9490 2972 9496 2984
rect 6871 2944 7788 2972
rect 9451 2944 9496 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 7653 2907 7711 2913
rect 7653 2873 7665 2907
rect 7699 2873 7711 2907
rect 7760 2904 7788 2944
rect 9490 2932 9496 2944
rect 9548 2932 9554 2984
rect 10505 2975 10563 2981
rect 10505 2941 10517 2975
rect 10551 2972 10563 2975
rect 10686 2972 10692 2984
rect 10551 2944 10692 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 10686 2932 10692 2944
rect 10744 2932 10750 2984
rect 11072 2972 11100 3000
rect 11716 2972 11744 3003
rect 13906 3000 13912 3052
rect 13964 3040 13970 3052
rect 14921 3043 14979 3049
rect 14921 3040 14933 3043
rect 13964 3012 14933 3040
rect 13964 3000 13970 3012
rect 14921 3009 14933 3012
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 15381 3043 15439 3049
rect 15381 3009 15393 3043
rect 15427 3040 15439 3043
rect 15657 3043 15715 3049
rect 15657 3040 15669 3043
rect 15427 3012 15669 3040
rect 15427 3009 15439 3012
rect 15381 3003 15439 3009
rect 15657 3009 15669 3012
rect 15703 3009 15715 3043
rect 17678 3040 17684 3052
rect 15657 3003 15715 3009
rect 16868 3012 17684 3040
rect 11072 2944 11744 2972
rect 14001 2975 14059 2981
rect 14001 2941 14013 2975
rect 14047 2972 14059 2975
rect 14642 2972 14648 2984
rect 14047 2944 14648 2972
rect 14047 2941 14059 2944
rect 14001 2935 14059 2941
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 15562 2981 15568 2984
rect 14737 2975 14795 2981
rect 14737 2941 14749 2975
rect 14783 2972 14795 2975
rect 15504 2975 15568 2981
rect 14783 2944 14964 2972
rect 14783 2941 14795 2944
rect 14737 2935 14795 2941
rect 11238 2904 11244 2916
rect 7760 2876 11244 2904
rect 7653 2867 7711 2873
rect 5902 2836 5908 2848
rect 1596 2808 5764 2836
rect 5863 2808 5908 2836
rect 5902 2796 5908 2808
rect 5960 2796 5966 2848
rect 5994 2796 6000 2848
rect 6052 2836 6058 2848
rect 7668 2836 7696 2867
rect 11238 2864 11244 2876
rect 11296 2864 11302 2916
rect 11514 2904 11520 2916
rect 11475 2876 11520 2904
rect 11514 2864 11520 2876
rect 11572 2864 11578 2916
rect 12526 2864 12532 2916
rect 12584 2904 12590 2916
rect 12805 2907 12863 2913
rect 12805 2904 12817 2907
rect 12584 2876 12817 2904
rect 12584 2864 12590 2876
rect 12805 2873 12817 2876
rect 12851 2873 12863 2907
rect 12805 2867 12863 2873
rect 14277 2907 14335 2913
rect 14277 2873 14289 2907
rect 14323 2904 14335 2907
rect 14826 2904 14832 2916
rect 14323 2876 14832 2904
rect 14323 2873 14335 2876
rect 14277 2867 14335 2873
rect 14826 2864 14832 2876
rect 14884 2864 14890 2916
rect 14936 2904 14964 2944
rect 15504 2941 15516 2975
rect 15550 2941 15568 2975
rect 15504 2935 15568 2941
rect 15562 2932 15568 2935
rect 15620 2932 15626 2984
rect 16209 2975 16267 2981
rect 16209 2941 16221 2975
rect 16255 2972 16267 2975
rect 16666 2972 16672 2984
rect 16255 2944 16672 2972
rect 16255 2941 16267 2944
rect 16209 2935 16267 2941
rect 16666 2932 16672 2944
rect 16724 2932 16730 2984
rect 16868 2981 16896 3012
rect 17678 3000 17684 3012
rect 17736 3000 17742 3052
rect 16853 2975 16911 2981
rect 16853 2941 16865 2975
rect 16899 2941 16911 2975
rect 16853 2935 16911 2941
rect 17034 2932 17040 2984
rect 17092 2972 17098 2984
rect 18064 2981 18092 3148
rect 17405 2975 17463 2981
rect 17405 2972 17417 2975
rect 17092 2944 17417 2972
rect 17092 2932 17098 2944
rect 17405 2941 17417 2944
rect 17451 2941 17463 2975
rect 17405 2935 17463 2941
rect 18049 2975 18107 2981
rect 18049 2941 18061 2975
rect 18095 2941 18107 2975
rect 18049 2935 18107 2941
rect 15194 2904 15200 2916
rect 14936 2876 15200 2904
rect 15194 2864 15200 2876
rect 15252 2864 15258 2916
rect 8110 2836 8116 2848
rect 6052 2808 6097 2836
rect 7668 2808 8116 2836
rect 6052 2796 6058 2808
rect 8110 2796 8116 2808
rect 8168 2796 8174 2848
rect 8386 2796 8392 2848
rect 8444 2836 8450 2848
rect 8481 2839 8539 2845
rect 8481 2836 8493 2839
rect 8444 2808 8493 2836
rect 8444 2796 8450 2808
rect 8481 2805 8493 2808
rect 8527 2805 8539 2839
rect 8481 2799 8539 2805
rect 8570 2796 8576 2848
rect 8628 2836 8634 2848
rect 8628 2808 8673 2836
rect 8628 2796 8634 2808
rect 8754 2796 8760 2848
rect 8812 2836 8818 2848
rect 10870 2836 10876 2848
rect 8812 2808 10876 2836
rect 8812 2796 8818 2808
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 11149 2839 11207 2845
rect 11149 2805 11161 2839
rect 11195 2836 11207 2839
rect 12897 2839 12955 2845
rect 12897 2836 12909 2839
rect 11195 2808 12909 2836
rect 11195 2805 11207 2808
rect 11149 2799 11207 2805
rect 12897 2805 12909 2808
rect 12943 2805 12955 2839
rect 16390 2836 16396 2848
rect 16351 2808 16396 2836
rect 12897 2799 12955 2805
rect 16390 2796 16396 2808
rect 16448 2796 16454 2848
rect 17034 2836 17040 2848
rect 16995 2808 17040 2836
rect 17034 2796 17040 2808
rect 17092 2796 17098 2848
rect 17589 2839 17647 2845
rect 17589 2805 17601 2839
rect 17635 2836 17647 2839
rect 17678 2836 17684 2848
rect 17635 2808 17684 2836
rect 17635 2805 17647 2808
rect 17589 2799 17647 2805
rect 17678 2796 17684 2808
rect 17736 2796 17742 2848
rect 18230 2836 18236 2848
rect 18191 2808 18236 2836
rect 18230 2796 18236 2808
rect 18288 2796 18294 2848
rect 1104 2746 18860 2768
rect 1104 2694 6912 2746
rect 6964 2694 6976 2746
rect 7028 2694 7040 2746
rect 7092 2694 7104 2746
rect 7156 2694 12843 2746
rect 12895 2694 12907 2746
rect 12959 2694 12971 2746
rect 13023 2694 13035 2746
rect 13087 2694 18860 2746
rect 1104 2672 18860 2694
rect 1854 2632 1860 2644
rect 1815 2604 1860 2632
rect 1854 2592 1860 2604
rect 1912 2592 1918 2644
rect 2682 2592 2688 2644
rect 2740 2632 2746 2644
rect 3329 2635 3387 2641
rect 3329 2632 3341 2635
rect 2740 2604 3341 2632
rect 2740 2592 2746 2604
rect 3329 2601 3341 2604
rect 3375 2601 3387 2635
rect 3329 2595 3387 2601
rect 3421 2635 3479 2641
rect 3421 2601 3433 2635
rect 3467 2632 3479 2635
rect 3510 2632 3516 2644
rect 3467 2604 3516 2632
rect 3467 2601 3479 2604
rect 3421 2595 3479 2601
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 4893 2635 4951 2641
rect 4893 2601 4905 2635
rect 4939 2632 4951 2635
rect 5166 2632 5172 2644
rect 4939 2604 5172 2632
rect 4939 2601 4951 2604
rect 4893 2595 4951 2601
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 5261 2635 5319 2641
rect 5261 2601 5273 2635
rect 5307 2632 5319 2635
rect 6365 2635 6423 2641
rect 6365 2632 6377 2635
rect 5307 2604 6377 2632
rect 5307 2601 5319 2604
rect 5261 2595 5319 2601
rect 6365 2601 6377 2604
rect 6411 2601 6423 2635
rect 6365 2595 6423 2601
rect 9033 2635 9091 2641
rect 9033 2601 9045 2635
rect 9079 2632 9091 2635
rect 9766 2632 9772 2644
rect 9079 2604 9772 2632
rect 9079 2601 9091 2604
rect 9033 2595 9091 2601
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 10229 2635 10287 2641
rect 10229 2601 10241 2635
rect 10275 2601 10287 2635
rect 10229 2595 10287 2601
rect 10689 2635 10747 2641
rect 10689 2601 10701 2635
rect 10735 2632 10747 2635
rect 10962 2632 10968 2644
rect 10735 2604 10968 2632
rect 10735 2601 10747 2604
rect 10689 2595 10747 2601
rect 4246 2564 4252 2576
rect 1688 2536 4252 2564
rect 1688 2505 1716 2536
rect 4246 2524 4252 2536
rect 4304 2524 4310 2576
rect 4801 2567 4859 2573
rect 4801 2533 4813 2567
rect 4847 2564 4859 2567
rect 6086 2564 6092 2576
rect 4847 2536 6092 2564
rect 4847 2533 4859 2536
rect 4801 2527 4859 2533
rect 6086 2524 6092 2536
rect 6144 2524 6150 2576
rect 7466 2564 7472 2576
rect 6196 2536 7472 2564
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2465 1731 2499
rect 1673 2459 1731 2465
rect 1946 2456 1952 2508
rect 2004 2496 2010 2508
rect 2225 2499 2283 2505
rect 2225 2496 2237 2499
rect 2004 2468 2237 2496
rect 2004 2456 2010 2468
rect 2225 2465 2237 2468
rect 2271 2465 2283 2499
rect 2225 2459 2283 2465
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 5261 2499 5319 2505
rect 5261 2496 5273 2499
rect 4120 2468 5273 2496
rect 4120 2456 4126 2468
rect 5261 2465 5273 2468
rect 5307 2465 5319 2499
rect 5442 2496 5448 2508
rect 5403 2468 5448 2496
rect 5261 2459 5319 2465
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 6196 2505 6224 2536
rect 7466 2524 7472 2536
rect 7524 2524 7530 2576
rect 10244 2564 10272 2595
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 11698 2632 11704 2644
rect 11659 2604 11704 2632
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 11609 2567 11667 2573
rect 11609 2564 11621 2567
rect 10244 2536 11621 2564
rect 11609 2533 11621 2536
rect 11655 2533 11667 2567
rect 11609 2527 11667 2533
rect 11882 2524 11888 2576
rect 11940 2564 11946 2576
rect 12897 2567 12955 2573
rect 12897 2564 12909 2567
rect 11940 2536 12909 2564
rect 11940 2524 11946 2536
rect 12897 2533 12909 2536
rect 12943 2533 12955 2567
rect 15286 2564 15292 2576
rect 12897 2527 12955 2533
rect 13372 2536 15292 2564
rect 6181 2499 6239 2505
rect 6181 2465 6193 2499
rect 6227 2465 6239 2499
rect 6181 2459 6239 2465
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7374 2496 7380 2508
rect 6963 2468 7380 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7374 2456 7380 2468
rect 7432 2456 7438 2508
rect 7745 2499 7803 2505
rect 7745 2465 7757 2499
rect 7791 2496 7803 2499
rect 7834 2496 7840 2508
rect 7791 2468 7840 2496
rect 7791 2465 7803 2468
rect 7745 2459 7803 2465
rect 7834 2456 7840 2468
rect 7892 2456 7898 2508
rect 10597 2499 10655 2505
rect 10597 2465 10609 2499
rect 10643 2496 10655 2499
rect 10778 2496 10784 2508
rect 10643 2468 10784 2496
rect 10643 2465 10655 2468
rect 10597 2459 10655 2465
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 11422 2456 11428 2508
rect 11480 2496 11486 2508
rect 13372 2505 13400 2536
rect 15286 2524 15292 2536
rect 15344 2524 15350 2576
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 11480 2468 12633 2496
rect 11480 2456 11486 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 13357 2499 13415 2505
rect 13357 2465 13369 2499
rect 13403 2465 13415 2499
rect 13357 2459 13415 2465
rect 14093 2499 14151 2505
rect 14093 2465 14105 2499
rect 14139 2496 14151 2499
rect 14182 2496 14188 2508
rect 14139 2468 14188 2496
rect 14139 2465 14151 2468
rect 14093 2459 14151 2465
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 17405 2499 17463 2505
rect 17405 2496 17417 2499
rect 14516 2468 17417 2496
rect 14516 2456 14522 2468
rect 17405 2465 17417 2468
rect 17451 2465 17463 2499
rect 17405 2459 17463 2465
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2428 2559 2431
rect 3050 2428 3056 2440
rect 2547 2400 3056 2428
rect 2547 2397 2559 2400
rect 2501 2391 2559 2397
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 3694 2428 3700 2440
rect 3651 2400 3700 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 3694 2388 3700 2400
rect 3752 2428 3758 2440
rect 4985 2431 5043 2437
rect 4985 2428 4997 2431
rect 3752 2400 4997 2428
rect 3752 2388 3758 2400
rect 4985 2397 4997 2400
rect 5031 2397 5043 2431
rect 5626 2428 5632 2440
rect 5587 2400 5632 2428
rect 4985 2391 5043 2397
rect 5626 2388 5632 2400
rect 5684 2388 5690 2440
rect 7101 2431 7159 2437
rect 7101 2397 7113 2431
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 2961 2363 3019 2369
rect 2961 2329 2973 2363
rect 3007 2360 3019 2363
rect 3326 2360 3332 2372
rect 3007 2332 3332 2360
rect 3007 2329 3019 2332
rect 2961 2323 3019 2329
rect 3326 2320 3332 2332
rect 3384 2320 3390 2372
rect 4890 2320 4896 2372
rect 4948 2360 4954 2372
rect 7116 2360 7144 2391
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 7616 2400 7941 2428
rect 7616 2388 7622 2400
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 10318 2428 10324 2440
rect 9355 2400 10324 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 4948 2332 7144 2360
rect 9140 2360 9168 2391
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 10873 2431 10931 2437
rect 10873 2397 10885 2431
rect 10919 2428 10931 2431
rect 11054 2428 11060 2440
rect 10919 2400 11060 2428
rect 10919 2397 10931 2400
rect 10873 2391 10931 2397
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 11793 2431 11851 2437
rect 11793 2428 11805 2431
rect 11204 2400 11805 2428
rect 11204 2388 11210 2400
rect 11793 2397 11805 2400
rect 11839 2397 11851 2431
rect 11793 2391 11851 2397
rect 13078 2388 13084 2440
rect 13136 2428 13142 2440
rect 13541 2431 13599 2437
rect 13541 2428 13553 2431
rect 13136 2400 13553 2428
rect 13136 2388 13142 2400
rect 13541 2397 13553 2400
rect 13587 2397 13599 2431
rect 13541 2391 13599 2397
rect 14277 2431 14335 2437
rect 14277 2397 14289 2431
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 11241 2363 11299 2369
rect 11241 2360 11253 2363
rect 9140 2332 11253 2360
rect 4948 2320 4954 2332
rect 11241 2329 11253 2332
rect 11287 2329 11299 2363
rect 11241 2323 11299 2329
rect 12158 2320 12164 2372
rect 12216 2360 12222 2372
rect 14292 2360 14320 2391
rect 12216 2332 14320 2360
rect 12216 2320 12222 2332
rect 4433 2295 4491 2301
rect 4433 2261 4445 2295
rect 4479 2292 4491 2295
rect 5994 2292 6000 2304
rect 4479 2264 6000 2292
rect 4479 2261 4491 2264
rect 4433 2255 4491 2261
rect 5994 2252 6000 2264
rect 6052 2252 6058 2304
rect 8665 2295 8723 2301
rect 8665 2261 8677 2295
rect 8711 2292 8723 2295
rect 11422 2292 11428 2304
rect 8711 2264 11428 2292
rect 8711 2261 8723 2264
rect 8665 2255 8723 2261
rect 11422 2252 11428 2264
rect 11480 2252 11486 2304
rect 17586 2292 17592 2304
rect 17547 2264 17592 2292
rect 17586 2252 17592 2264
rect 17644 2252 17650 2304
rect 1104 2202 18860 2224
rect 1104 2150 3947 2202
rect 3999 2150 4011 2202
rect 4063 2150 4075 2202
rect 4127 2150 4139 2202
rect 4191 2150 9878 2202
rect 9930 2150 9942 2202
rect 9994 2150 10006 2202
rect 10058 2150 10070 2202
rect 10122 2150 15808 2202
rect 15860 2150 15872 2202
rect 15924 2150 15936 2202
rect 15988 2150 16000 2202
rect 16052 2150 18860 2202
rect 1104 2128 18860 2150
rect 3694 2048 3700 2100
rect 3752 2088 3758 2100
rect 5074 2088 5080 2100
rect 3752 2060 5080 2088
rect 3752 2048 3758 2060
rect 5074 2048 5080 2060
rect 5132 2048 5138 2100
rect 9398 2048 9404 2100
rect 9456 2088 9462 2100
rect 11882 2088 11888 2100
rect 9456 2060 11888 2088
rect 9456 2048 9462 2060
rect 11882 2048 11888 2060
rect 11940 2048 11946 2100
rect 11238 1504 11244 1556
rect 11296 1544 11302 1556
rect 19426 1544 19432 1556
rect 11296 1516 19432 1544
rect 11296 1504 11302 1516
rect 19426 1504 19432 1516
rect 19484 1504 19490 1556
rect 3970 1368 3976 1420
rect 4028 1408 4034 1420
rect 5626 1408 5632 1420
rect 4028 1380 5632 1408
rect 4028 1368 4034 1380
rect 5626 1368 5632 1380
rect 5684 1368 5690 1420
rect 3326 1300 3332 1352
rect 3384 1340 3390 1352
rect 12066 1340 12072 1352
rect 3384 1312 12072 1340
rect 3384 1300 3390 1312
rect 12066 1300 12072 1312
rect 12124 1300 12130 1352
rect 382 960 388 1012
rect 440 1000 446 1012
rect 8754 1000 8760 1012
rect 440 972 8760 1000
rect 440 960 446 972
rect 8754 960 8760 972
rect 8812 960 8818 1012
<< via1 >>
rect 4068 15172 4120 15224
rect 9496 15172 9548 15224
rect 6912 14662 6964 14714
rect 6976 14662 7028 14714
rect 7040 14662 7092 14714
rect 7104 14662 7156 14714
rect 12843 14662 12895 14714
rect 12907 14662 12959 14714
rect 12971 14662 13023 14714
rect 13035 14662 13087 14714
rect 3424 14560 3476 14612
rect 11152 14560 11204 14612
rect 5356 14492 5408 14544
rect 14280 14492 14332 14544
rect 4528 14467 4580 14476
rect 4528 14433 4537 14467
rect 4537 14433 4571 14467
rect 4571 14433 4580 14467
rect 4528 14424 4580 14433
rect 10048 14424 10100 14476
rect 10416 14424 10468 14476
rect 13912 14424 13964 14476
rect 14372 14424 14424 14476
rect 18788 14492 18840 14544
rect 17408 14467 17460 14476
rect 17408 14433 17417 14467
rect 17417 14433 17451 14467
rect 17451 14433 17460 14467
rect 17408 14424 17460 14433
rect 3056 14356 3108 14408
rect 4712 14399 4764 14408
rect 4712 14365 4721 14399
rect 4721 14365 4755 14399
rect 4755 14365 4764 14399
rect 4712 14356 4764 14365
rect 10508 14356 10560 14408
rect 11060 14356 11112 14408
rect 15384 14356 15436 14408
rect 17500 14399 17552 14408
rect 17500 14365 17509 14399
rect 17509 14365 17543 14399
rect 17543 14365 17552 14399
rect 17500 14356 17552 14365
rect 17684 14399 17736 14408
rect 17684 14365 17693 14399
rect 17693 14365 17727 14399
rect 17727 14365 17736 14399
rect 17684 14356 17736 14365
rect 3332 14288 3384 14340
rect 18052 14288 18104 14340
rect 9680 14220 9732 14272
rect 10784 14220 10836 14272
rect 15660 14220 15712 14272
rect 17040 14263 17092 14272
rect 17040 14229 17049 14263
rect 17049 14229 17083 14263
rect 17083 14229 17092 14263
rect 17040 14220 17092 14229
rect 3947 14118 3999 14170
rect 4011 14118 4063 14170
rect 4075 14118 4127 14170
rect 4139 14118 4191 14170
rect 9878 14118 9930 14170
rect 9942 14118 9994 14170
rect 10006 14118 10058 14170
rect 10070 14118 10122 14170
rect 15808 14118 15860 14170
rect 15872 14118 15924 14170
rect 15936 14118 15988 14170
rect 16000 14118 16052 14170
rect 4528 14016 4580 14068
rect 10692 14016 10744 14068
rect 2964 13948 3016 14000
rect 3608 13948 3660 14000
rect 2688 13880 2740 13932
rect 4804 13880 4856 13932
rect 5356 13923 5408 13932
rect 5356 13889 5365 13923
rect 5365 13889 5399 13923
rect 5399 13889 5408 13923
rect 5356 13880 5408 13889
rect 5448 13923 5500 13932
rect 5448 13889 5457 13923
rect 5457 13889 5491 13923
rect 5491 13889 5500 13923
rect 7472 13923 7524 13932
rect 5448 13880 5500 13889
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 2780 13812 2832 13864
rect 6644 13812 6696 13864
rect 8116 13812 8168 13864
rect 10600 13948 10652 14000
rect 10508 13880 10560 13932
rect 13452 14016 13504 14068
rect 16212 14016 16264 14068
rect 14740 13948 14792 14000
rect 14924 13948 14976 14000
rect 11060 13880 11112 13932
rect 12164 13880 12216 13932
rect 13912 13880 13964 13932
rect 14188 13923 14240 13932
rect 14188 13889 14197 13923
rect 14197 13889 14231 13923
rect 14231 13889 14240 13923
rect 14188 13880 14240 13889
rect 17132 13948 17184 14000
rect 17684 13948 17736 14000
rect 18512 13948 18564 14000
rect 16580 13880 16632 13932
rect 17592 13880 17644 13932
rect 9588 13812 9640 13864
rect 9680 13812 9732 13864
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 13268 13812 13320 13864
rect 1952 13676 2004 13728
rect 4344 13719 4396 13728
rect 4344 13685 4353 13719
rect 4353 13685 4387 13719
rect 4387 13685 4396 13719
rect 5540 13744 5592 13796
rect 4344 13676 4396 13685
rect 5264 13719 5316 13728
rect 5264 13685 5273 13719
rect 5273 13685 5307 13719
rect 5307 13685 5316 13719
rect 5264 13676 5316 13685
rect 6368 13676 6420 13728
rect 10140 13744 10192 13796
rect 10324 13744 10376 13796
rect 10508 13676 10560 13728
rect 10692 13676 10744 13728
rect 11244 13744 11296 13796
rect 15200 13855 15252 13864
rect 15200 13821 15209 13855
rect 15209 13821 15243 13855
rect 15243 13821 15252 13855
rect 15200 13812 15252 13821
rect 15660 13812 15712 13864
rect 17224 13855 17276 13864
rect 13268 13676 13320 13728
rect 13912 13719 13964 13728
rect 13912 13685 13921 13719
rect 13921 13685 13955 13719
rect 13955 13685 13964 13719
rect 13912 13676 13964 13685
rect 14832 13719 14884 13728
rect 14832 13685 14841 13719
rect 14841 13685 14875 13719
rect 14875 13685 14884 13719
rect 14832 13676 14884 13685
rect 15292 13744 15344 13796
rect 17224 13821 17233 13855
rect 17233 13821 17267 13855
rect 17267 13821 17276 13855
rect 17224 13812 17276 13821
rect 18052 13855 18104 13864
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 6912 13574 6964 13626
rect 6976 13574 7028 13626
rect 7040 13574 7092 13626
rect 7104 13574 7156 13626
rect 12843 13574 12895 13626
rect 12907 13574 12959 13626
rect 12971 13574 13023 13626
rect 13035 13574 13087 13626
rect 2872 13515 2924 13524
rect 2872 13481 2881 13515
rect 2881 13481 2915 13515
rect 2915 13481 2924 13515
rect 2872 13472 2924 13481
rect 4068 13472 4120 13524
rect 4344 13472 4396 13524
rect 6368 13515 6420 13524
rect 6368 13481 6377 13515
rect 6377 13481 6411 13515
rect 6411 13481 6420 13515
rect 6368 13472 6420 13481
rect 7472 13472 7524 13524
rect 9956 13472 10008 13524
rect 11152 13472 11204 13524
rect 11520 13472 11572 13524
rect 13268 13515 13320 13524
rect 13268 13481 13277 13515
rect 13277 13481 13311 13515
rect 13311 13481 13320 13515
rect 13268 13472 13320 13481
rect 13912 13472 13964 13524
rect 15292 13515 15344 13524
rect 15292 13481 15301 13515
rect 15301 13481 15335 13515
rect 15335 13481 15344 13515
rect 15292 13472 15344 13481
rect 17960 13515 18012 13524
rect 17960 13481 17969 13515
rect 17969 13481 18003 13515
rect 18003 13481 18012 13515
rect 17960 13472 18012 13481
rect 1768 13336 1820 13388
rect 1124 13268 1176 13320
rect 3148 13336 3200 13388
rect 3792 13336 3844 13388
rect 2688 13268 2740 13320
rect 2044 13200 2096 13252
rect 5356 13336 5408 13388
rect 6276 13379 6328 13388
rect 6276 13345 6285 13379
rect 6285 13345 6319 13379
rect 6319 13345 6328 13379
rect 6276 13336 6328 13345
rect 7748 13404 7800 13456
rect 12440 13404 12492 13456
rect 8300 13336 8352 13388
rect 10692 13336 10744 13388
rect 13912 13379 13964 13388
rect 5448 13311 5500 13320
rect 5448 13277 5457 13311
rect 5457 13277 5491 13311
rect 5491 13277 5500 13311
rect 6552 13311 6604 13320
rect 5448 13268 5500 13277
rect 6552 13277 6561 13311
rect 6561 13277 6595 13311
rect 6595 13277 6604 13311
rect 6552 13268 6604 13277
rect 6920 13311 6972 13320
rect 6920 13277 6929 13311
rect 6929 13277 6963 13311
rect 6963 13277 6972 13311
rect 6920 13268 6972 13277
rect 9036 13311 9088 13320
rect 9036 13277 9045 13311
rect 9045 13277 9079 13311
rect 9079 13277 9088 13311
rect 9036 13268 9088 13277
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 11152 13311 11204 13320
rect 11152 13277 11161 13311
rect 11161 13277 11195 13311
rect 11195 13277 11204 13311
rect 11152 13268 11204 13277
rect 11336 13311 11388 13320
rect 11336 13277 11345 13311
rect 11345 13277 11379 13311
rect 11379 13277 11388 13311
rect 11336 13268 11388 13277
rect 11888 13311 11940 13320
rect 11888 13277 11897 13311
rect 11897 13277 11931 13311
rect 11931 13277 11940 13311
rect 11888 13268 11940 13277
rect 2228 13132 2280 13184
rect 4344 13132 4396 13184
rect 9772 13200 9824 13252
rect 9864 13200 9916 13252
rect 9956 13200 10008 13252
rect 11704 13200 11756 13252
rect 13912 13345 13921 13379
rect 13921 13345 13955 13379
rect 13955 13345 13964 13379
rect 13912 13336 13964 13345
rect 15568 13336 15620 13388
rect 14004 13311 14056 13320
rect 14004 13277 14013 13311
rect 14013 13277 14047 13311
rect 14047 13277 14056 13311
rect 14004 13268 14056 13277
rect 14096 13311 14148 13320
rect 14096 13277 14105 13311
rect 14105 13277 14139 13311
rect 14139 13277 14148 13311
rect 16948 13336 17000 13388
rect 17868 13379 17920 13388
rect 17868 13345 17877 13379
rect 17877 13345 17911 13379
rect 17911 13345 17920 13379
rect 17868 13336 17920 13345
rect 14096 13268 14148 13277
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 16856 13311 16908 13320
rect 16856 13277 16865 13311
rect 16865 13277 16899 13311
rect 16899 13277 16908 13311
rect 16856 13268 16908 13277
rect 14188 13200 14240 13252
rect 15660 13200 15712 13252
rect 17684 13200 17736 13252
rect 9680 13175 9732 13184
rect 9680 13141 9689 13175
rect 9689 13141 9723 13175
rect 9723 13141 9732 13175
rect 9680 13132 9732 13141
rect 12624 13132 12676 13184
rect 15476 13132 15528 13184
rect 17316 13132 17368 13184
rect 3947 13030 3999 13082
rect 4011 13030 4063 13082
rect 4075 13030 4127 13082
rect 4139 13030 4191 13082
rect 9878 13030 9930 13082
rect 9942 13030 9994 13082
rect 10006 13030 10058 13082
rect 10070 13030 10122 13082
rect 15808 13030 15860 13082
rect 15872 13030 15924 13082
rect 15936 13030 15988 13082
rect 16000 13030 16052 13082
rect 1768 12971 1820 12980
rect 1768 12937 1777 12971
rect 1777 12937 1811 12971
rect 1811 12937 1820 12971
rect 1768 12928 1820 12937
rect 4252 12928 4304 12980
rect 4712 12928 4764 12980
rect 4804 12928 4856 12980
rect 6552 12928 6604 12980
rect 9128 12928 9180 12980
rect 2044 12792 2096 12844
rect 7932 12792 7984 12844
rect 4436 12724 4488 12776
rect 5080 12767 5132 12776
rect 5080 12733 5114 12767
rect 5114 12733 5132 12767
rect 5080 12724 5132 12733
rect 5448 12724 5500 12776
rect 2320 12656 2372 12708
rect 3608 12656 3660 12708
rect 4712 12656 4764 12708
rect 2136 12631 2188 12640
rect 2136 12597 2145 12631
rect 2145 12597 2179 12631
rect 2179 12597 2188 12631
rect 2136 12588 2188 12597
rect 3976 12588 4028 12640
rect 6736 12656 6788 12708
rect 7472 12724 7524 12776
rect 6920 12656 6972 12708
rect 7656 12724 7708 12776
rect 11244 12928 11296 12980
rect 11336 12928 11388 12980
rect 15568 12928 15620 12980
rect 16948 12971 17000 12980
rect 16948 12937 16957 12971
rect 16957 12937 16991 12971
rect 16991 12937 17000 12971
rect 16948 12928 17000 12937
rect 14188 12860 14240 12912
rect 16488 12835 16540 12844
rect 16488 12801 16497 12835
rect 16497 12801 16531 12835
rect 16531 12801 16540 12835
rect 16488 12792 16540 12801
rect 17776 12792 17828 12844
rect 11428 12724 11480 12776
rect 11888 12724 11940 12776
rect 9220 12656 9272 12708
rect 10324 12656 10376 12708
rect 11244 12656 11296 12708
rect 13820 12724 13872 12776
rect 15292 12724 15344 12776
rect 17316 12767 17368 12776
rect 17316 12733 17325 12767
rect 17325 12733 17359 12767
rect 17359 12733 17368 12767
rect 17316 12724 17368 12733
rect 14096 12656 14148 12708
rect 14464 12656 14516 12708
rect 16304 12699 16356 12708
rect 16304 12665 16313 12699
rect 16313 12665 16347 12699
rect 16347 12665 16356 12699
rect 16304 12656 16356 12665
rect 5356 12588 5408 12640
rect 7932 12588 7984 12640
rect 8116 12588 8168 12640
rect 11612 12588 11664 12640
rect 16396 12631 16448 12640
rect 16396 12597 16405 12631
rect 16405 12597 16439 12631
rect 16439 12597 16448 12631
rect 16396 12588 16448 12597
rect 16580 12588 16632 12640
rect 6912 12486 6964 12538
rect 6976 12486 7028 12538
rect 7040 12486 7092 12538
rect 7104 12486 7156 12538
rect 12843 12486 12895 12538
rect 12907 12486 12959 12538
rect 12971 12486 13023 12538
rect 13035 12486 13087 12538
rect 3056 12384 3108 12436
rect 4344 12316 4396 12368
rect 5172 12316 5224 12368
rect 8300 12384 8352 12436
rect 9036 12384 9088 12436
rect 11152 12384 11204 12436
rect 11336 12384 11388 12436
rect 11612 12384 11664 12436
rect 13268 12384 13320 12436
rect 14004 12384 14056 12436
rect 15660 12427 15712 12436
rect 15660 12393 15669 12427
rect 15669 12393 15703 12427
rect 15703 12393 15712 12427
rect 15660 12384 15712 12393
rect 17040 12384 17092 12436
rect 6736 12316 6788 12368
rect 8484 12316 8536 12368
rect 1952 12155 2004 12164
rect 1952 12121 1961 12155
rect 1961 12121 1995 12155
rect 1995 12121 2004 12155
rect 1952 12112 2004 12121
rect 4896 12291 4948 12300
rect 4896 12257 4905 12291
rect 4905 12257 4939 12291
rect 4939 12257 4948 12291
rect 4896 12248 4948 12257
rect 6368 12248 6420 12300
rect 8852 12248 8904 12300
rect 9404 12248 9456 12300
rect 2412 12223 2464 12232
rect 2412 12189 2421 12223
rect 2421 12189 2455 12223
rect 2455 12189 2464 12223
rect 2412 12180 2464 12189
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 3608 12223 3660 12232
rect 2596 12180 2648 12189
rect 3608 12189 3617 12223
rect 3617 12189 3651 12223
rect 3651 12189 3660 12223
rect 3608 12180 3660 12189
rect 4160 12180 4212 12232
rect 5080 12223 5132 12232
rect 5080 12189 5089 12223
rect 5089 12189 5123 12223
rect 5123 12189 5132 12223
rect 5080 12180 5132 12189
rect 5540 12180 5592 12232
rect 7012 12223 7064 12232
rect 3516 12112 3568 12164
rect 4620 12112 4672 12164
rect 7012 12189 7021 12223
rect 7021 12189 7055 12223
rect 7055 12189 7064 12223
rect 7012 12180 7064 12189
rect 7380 12180 7432 12232
rect 7564 12180 7616 12232
rect 8116 12180 8168 12232
rect 9036 12223 9088 12232
rect 6920 12112 6972 12164
rect 7472 12112 7524 12164
rect 9036 12189 9045 12223
rect 9045 12189 9079 12223
rect 9079 12189 9088 12223
rect 9036 12180 9088 12189
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 11704 12316 11756 12368
rect 14096 12316 14148 12368
rect 14832 12316 14884 12368
rect 17132 12316 17184 12368
rect 9220 12180 9272 12189
rect 9312 12112 9364 12164
rect 10324 12112 10376 12164
rect 11980 12248 12032 12300
rect 12348 12291 12400 12300
rect 12348 12257 12357 12291
rect 12357 12257 12391 12291
rect 12391 12257 12400 12291
rect 12348 12248 12400 12257
rect 15108 12248 15160 12300
rect 15292 12248 15344 12300
rect 11244 12180 11296 12232
rect 11612 12180 11664 12232
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 13728 12180 13780 12232
rect 13820 12180 13872 12232
rect 14372 12223 14424 12232
rect 14372 12189 14381 12223
rect 14381 12189 14415 12223
rect 14415 12189 14424 12223
rect 14372 12180 14424 12189
rect 14464 12180 14516 12232
rect 16304 12112 16356 12164
rect 2872 12044 2924 12096
rect 3792 12044 3844 12096
rect 7288 12044 7340 12096
rect 8208 12044 8260 12096
rect 8300 12044 8352 12096
rect 10876 12044 10928 12096
rect 11152 12044 11204 12096
rect 14188 12044 14240 12096
rect 16488 12180 16540 12232
rect 3947 11942 3999 11994
rect 4011 11942 4063 11994
rect 4075 11942 4127 11994
rect 4139 11942 4191 11994
rect 9878 11942 9930 11994
rect 9942 11942 9994 11994
rect 10006 11942 10058 11994
rect 10070 11942 10122 11994
rect 15808 11942 15860 11994
rect 15872 11942 15924 11994
rect 15936 11942 15988 11994
rect 16000 11942 16052 11994
rect 2412 11840 2464 11892
rect 3792 11840 3844 11892
rect 2780 11772 2832 11824
rect 6276 11840 6328 11892
rect 8944 11883 8996 11892
rect 8944 11849 8953 11883
rect 8953 11849 8987 11883
rect 8987 11849 8996 11883
rect 8944 11840 8996 11849
rect 9036 11840 9088 11892
rect 11796 11840 11848 11892
rect 12348 11840 12400 11892
rect 13912 11840 13964 11892
rect 14004 11840 14056 11892
rect 14924 11840 14976 11892
rect 16396 11840 16448 11892
rect 7472 11772 7524 11824
rect 8576 11772 8628 11824
rect 10692 11815 10744 11824
rect 2044 11704 2096 11756
rect 2596 11704 2648 11756
rect 5264 11747 5316 11756
rect 2872 11568 2924 11620
rect 3516 11568 3568 11620
rect 2780 11500 2832 11552
rect 3424 11500 3476 11552
rect 5264 11713 5273 11747
rect 5273 11713 5307 11747
rect 5307 11713 5316 11747
rect 5264 11704 5316 11713
rect 6920 11704 6972 11756
rect 8852 11704 8904 11756
rect 10324 11747 10376 11756
rect 10324 11713 10333 11747
rect 10333 11713 10367 11747
rect 10367 11713 10376 11747
rect 10324 11704 10376 11713
rect 10692 11781 10701 11815
rect 10701 11781 10735 11815
rect 10735 11781 10744 11815
rect 10692 11772 10744 11781
rect 15016 11772 15068 11824
rect 17132 11772 17184 11824
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 11336 11747 11388 11756
rect 11336 11713 11345 11747
rect 11345 11713 11379 11747
rect 11379 11713 11388 11747
rect 11336 11704 11388 11713
rect 12072 11704 12124 11756
rect 14464 11747 14516 11756
rect 4252 11636 4304 11688
rect 4712 11636 4764 11688
rect 7012 11636 7064 11688
rect 7656 11636 7708 11688
rect 9128 11636 9180 11688
rect 3792 11568 3844 11620
rect 3976 11568 4028 11620
rect 10692 11636 10744 11688
rect 13728 11636 13780 11688
rect 4436 11500 4488 11552
rect 4988 11543 5040 11552
rect 4988 11509 4997 11543
rect 4997 11509 5031 11543
rect 5031 11509 5040 11543
rect 4988 11500 5040 11509
rect 6092 11543 6144 11552
rect 6092 11509 6101 11543
rect 6101 11509 6135 11543
rect 6135 11509 6144 11543
rect 6092 11500 6144 11509
rect 6368 11500 6420 11552
rect 9588 11500 9640 11552
rect 13912 11568 13964 11620
rect 14464 11713 14473 11747
rect 14473 11713 14507 11747
rect 14507 11713 14516 11747
rect 14464 11704 14516 11713
rect 15292 11747 15344 11756
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 16488 11704 16540 11756
rect 17408 11704 17460 11756
rect 16856 11636 16908 11688
rect 18144 11568 18196 11620
rect 10048 11543 10100 11552
rect 10048 11509 10057 11543
rect 10057 11509 10091 11543
rect 10091 11509 10100 11543
rect 10048 11500 10100 11509
rect 11704 11500 11756 11552
rect 13268 11500 13320 11552
rect 13636 11500 13688 11552
rect 14280 11543 14332 11552
rect 14280 11509 14289 11543
rect 14289 11509 14323 11543
rect 14323 11509 14332 11543
rect 14280 11500 14332 11509
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 6912 11398 6964 11450
rect 6976 11398 7028 11450
rect 7040 11398 7092 11450
rect 7104 11398 7156 11450
rect 12843 11398 12895 11450
rect 12907 11398 12959 11450
rect 12971 11398 13023 11450
rect 13035 11398 13087 11450
rect 2412 11296 2464 11348
rect 2688 11296 2740 11348
rect 2320 11228 2372 11280
rect 2596 11271 2648 11280
rect 2596 11237 2630 11271
rect 2630 11237 2648 11271
rect 2596 11228 2648 11237
rect 9312 11296 9364 11348
rect 9588 11296 9640 11348
rect 7012 11228 7064 11280
rect 3792 11160 3844 11212
rect 4988 11160 5040 11212
rect 6644 11160 6696 11212
rect 2044 11092 2096 11144
rect 3516 11092 3568 11144
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 5724 11092 5776 11144
rect 9128 11228 9180 11280
rect 10324 11296 10376 11348
rect 11244 11296 11296 11348
rect 12072 11296 12124 11348
rect 10692 11228 10744 11280
rect 8944 11160 8996 11212
rect 9588 11160 9640 11212
rect 11980 11228 12032 11280
rect 12624 11296 12676 11348
rect 13728 11296 13780 11348
rect 13912 11339 13964 11348
rect 13912 11305 13921 11339
rect 13921 11305 13955 11339
rect 13955 11305 13964 11339
rect 13912 11296 13964 11305
rect 15016 11296 15068 11348
rect 16856 11296 16908 11348
rect 13820 11228 13872 11280
rect 17776 11228 17828 11280
rect 1400 11024 1452 11076
rect 3332 11024 3384 11076
rect 3976 11024 4028 11076
rect 5816 11024 5868 11076
rect 6460 11067 6512 11076
rect 2596 10956 2648 11008
rect 6460 11033 6469 11067
rect 6469 11033 6503 11067
rect 6503 11033 6512 11067
rect 6460 11024 6512 11033
rect 7656 10956 7708 11008
rect 11704 11160 11756 11212
rect 14004 11160 14056 11212
rect 14280 11203 14332 11212
rect 14280 11169 14289 11203
rect 14289 11169 14323 11203
rect 14323 11169 14332 11203
rect 14280 11160 14332 11169
rect 14832 11160 14884 11212
rect 15292 11203 15344 11212
rect 15292 11169 15301 11203
rect 15301 11169 15335 11203
rect 15335 11169 15344 11203
rect 15292 11160 15344 11169
rect 16396 11160 16448 11212
rect 16672 11160 16724 11212
rect 17132 11160 17184 11212
rect 12256 11135 12308 11144
rect 12256 11101 12265 11135
rect 12265 11101 12299 11135
rect 12299 11101 12308 11135
rect 12256 11092 12308 11101
rect 13912 11092 13964 11144
rect 10324 10956 10376 11008
rect 10692 10956 10744 11008
rect 11428 10999 11480 11008
rect 11428 10965 11437 10999
rect 11437 10965 11471 10999
rect 11471 10965 11480 10999
rect 13360 11024 13412 11076
rect 15200 11092 15252 11144
rect 16948 11067 17000 11076
rect 16948 11033 16957 11067
rect 16957 11033 16991 11067
rect 16991 11033 17000 11067
rect 16948 11024 17000 11033
rect 17316 11024 17368 11076
rect 17684 11092 17736 11144
rect 11428 10956 11480 10965
rect 13176 10956 13228 11008
rect 17040 10956 17092 11008
rect 3947 10854 3999 10906
rect 4011 10854 4063 10906
rect 4075 10854 4127 10906
rect 4139 10854 4191 10906
rect 9878 10854 9930 10906
rect 9942 10854 9994 10906
rect 10006 10854 10058 10906
rect 10070 10854 10122 10906
rect 15808 10854 15860 10906
rect 15872 10854 15924 10906
rect 15936 10854 15988 10906
rect 16000 10854 16052 10906
rect 2780 10752 2832 10804
rect 5172 10752 5224 10804
rect 7012 10752 7064 10804
rect 8024 10752 8076 10804
rect 9128 10795 9180 10804
rect 4160 10684 4212 10736
rect 6000 10684 6052 10736
rect 3516 10616 3568 10668
rect 3792 10616 3844 10668
rect 5908 10616 5960 10668
rect 6276 10659 6328 10668
rect 6276 10625 6285 10659
rect 6285 10625 6319 10659
rect 6319 10625 6328 10659
rect 6276 10616 6328 10625
rect 7656 10616 7708 10668
rect 9128 10761 9137 10795
rect 9137 10761 9171 10795
rect 9171 10761 9180 10795
rect 9128 10752 9180 10761
rect 9496 10752 9548 10804
rect 8944 10684 8996 10736
rect 2412 10548 2464 10600
rect 7564 10548 7616 10600
rect 7840 10548 7892 10600
rect 2044 10480 2096 10532
rect 3424 10480 3476 10532
rect 2504 10412 2556 10464
rect 3240 10455 3292 10464
rect 3240 10421 3249 10455
rect 3249 10421 3283 10455
rect 3283 10421 3292 10455
rect 3240 10412 3292 10421
rect 4068 10455 4120 10464
rect 4068 10421 4077 10455
rect 4077 10421 4111 10455
rect 4111 10421 4120 10455
rect 4068 10412 4120 10421
rect 4712 10412 4764 10464
rect 5080 10455 5132 10464
rect 5080 10421 5089 10455
rect 5089 10421 5123 10455
rect 5123 10421 5132 10455
rect 5080 10412 5132 10421
rect 5172 10455 5224 10464
rect 5172 10421 5181 10455
rect 5181 10421 5215 10455
rect 5215 10421 5224 10455
rect 5172 10412 5224 10421
rect 5448 10412 5500 10464
rect 8024 10523 8076 10532
rect 6736 10412 6788 10464
rect 8024 10489 8058 10523
rect 8058 10489 8076 10523
rect 8024 10480 8076 10489
rect 8576 10412 8628 10464
rect 9680 10616 9732 10668
rect 10692 10659 10744 10668
rect 10692 10625 10701 10659
rect 10701 10625 10735 10659
rect 10735 10625 10744 10659
rect 10692 10616 10744 10625
rect 9772 10591 9824 10600
rect 9772 10557 9781 10591
rect 9781 10557 9815 10591
rect 9815 10557 9824 10591
rect 9772 10548 9824 10557
rect 16212 10752 16264 10804
rect 12072 10727 12124 10736
rect 12072 10693 12081 10727
rect 12081 10693 12115 10727
rect 12115 10693 12124 10727
rect 12072 10684 12124 10693
rect 16580 10752 16632 10804
rect 16672 10752 16724 10804
rect 17500 10752 17552 10804
rect 13084 10659 13136 10668
rect 13084 10625 13093 10659
rect 13093 10625 13127 10659
rect 13127 10625 13136 10659
rect 13084 10616 13136 10625
rect 14464 10616 14516 10668
rect 14648 10616 14700 10668
rect 13728 10591 13780 10600
rect 13728 10557 13762 10591
rect 13762 10557 13780 10591
rect 11704 10480 11756 10532
rect 12256 10480 12308 10532
rect 13728 10548 13780 10557
rect 14924 10548 14976 10600
rect 16120 10548 16172 10600
rect 16304 10591 16356 10600
rect 16304 10557 16313 10591
rect 16313 10557 16347 10591
rect 16347 10557 16356 10591
rect 16304 10548 16356 10557
rect 17868 10616 17920 10668
rect 17684 10548 17736 10600
rect 13820 10480 13872 10532
rect 12532 10412 12584 10464
rect 12716 10412 12768 10464
rect 13176 10412 13228 10464
rect 18052 10480 18104 10532
rect 14832 10455 14884 10464
rect 14832 10421 14841 10455
rect 14841 10421 14875 10455
rect 14875 10421 14884 10455
rect 14832 10412 14884 10421
rect 17592 10412 17644 10464
rect 17776 10412 17828 10464
rect 6912 10310 6964 10362
rect 6976 10310 7028 10362
rect 7040 10310 7092 10362
rect 7104 10310 7156 10362
rect 12843 10310 12895 10362
rect 12907 10310 12959 10362
rect 12971 10310 13023 10362
rect 13035 10310 13087 10362
rect 2228 10251 2280 10260
rect 2228 10217 2237 10251
rect 2237 10217 2271 10251
rect 2271 10217 2280 10251
rect 2228 10208 2280 10217
rect 2872 10208 2924 10260
rect 4436 10208 4488 10260
rect 5172 10208 5224 10260
rect 8116 10208 8168 10260
rect 8208 10208 8260 10260
rect 9128 10208 9180 10260
rect 9588 10208 9640 10260
rect 11980 10251 12032 10260
rect 2136 10140 2188 10192
rect 3976 10140 4028 10192
rect 5540 10140 5592 10192
rect 2964 10072 3016 10124
rect 3148 10072 3200 10124
rect 3424 10115 3476 10124
rect 3424 10081 3433 10115
rect 3433 10081 3467 10115
rect 3467 10081 3476 10115
rect 3424 10072 3476 10081
rect 2504 10047 2556 10056
rect 2504 10013 2513 10047
rect 2513 10013 2547 10047
rect 2547 10013 2556 10047
rect 2504 10004 2556 10013
rect 3516 10047 3568 10056
rect 3516 10013 3525 10047
rect 3525 10013 3559 10047
rect 3559 10013 3568 10047
rect 3516 10004 3568 10013
rect 5816 10072 5868 10124
rect 7656 10140 7708 10192
rect 7472 10072 7524 10124
rect 5356 10047 5408 10056
rect 4160 9936 4212 9988
rect 4896 9936 4948 9988
rect 1584 9868 1636 9920
rect 4252 9911 4304 9920
rect 4252 9877 4261 9911
rect 4261 9877 4295 9911
rect 4295 9877 4304 9911
rect 4252 9868 4304 9877
rect 5356 10013 5365 10047
rect 5365 10013 5399 10047
rect 5399 10013 5408 10047
rect 5356 10004 5408 10013
rect 8944 10140 8996 10192
rect 11980 10217 11989 10251
rect 11989 10217 12023 10251
rect 12023 10217 12032 10251
rect 11980 10208 12032 10217
rect 12256 10251 12308 10260
rect 12256 10217 12265 10251
rect 12265 10217 12299 10251
rect 12299 10217 12308 10251
rect 12256 10208 12308 10217
rect 13268 10251 13320 10260
rect 13268 10217 13277 10251
rect 13277 10217 13311 10251
rect 13311 10217 13320 10251
rect 13268 10208 13320 10217
rect 13452 10208 13504 10260
rect 14280 10251 14332 10260
rect 14280 10217 14289 10251
rect 14289 10217 14323 10251
rect 14323 10217 14332 10251
rect 14280 10208 14332 10217
rect 16212 10208 16264 10260
rect 16672 10208 16724 10260
rect 17684 10208 17736 10260
rect 10324 10140 10376 10192
rect 10692 10140 10744 10192
rect 11152 10140 11204 10192
rect 13544 10140 13596 10192
rect 5172 9936 5224 9988
rect 8024 9936 8076 9988
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8668 10047 8720 10056
rect 8208 10004 8260 10013
rect 8668 10013 8677 10047
rect 8677 10013 8711 10047
rect 8711 10013 8720 10047
rect 8668 10004 8720 10013
rect 12164 10115 12216 10124
rect 12164 10081 12173 10115
rect 12173 10081 12207 10115
rect 12207 10081 12216 10115
rect 12164 10072 12216 10081
rect 12624 10115 12676 10124
rect 12624 10081 12633 10115
rect 12633 10081 12667 10115
rect 12667 10081 12676 10115
rect 16120 10140 16172 10192
rect 16488 10140 16540 10192
rect 16580 10140 16632 10192
rect 17960 10140 18012 10192
rect 12624 10072 12676 10081
rect 9496 10004 9548 10056
rect 8760 9936 8812 9988
rect 12624 9936 12676 9988
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 13912 10047 13964 10056
rect 12808 10004 12860 10013
rect 13912 10013 13921 10047
rect 13921 10013 13955 10047
rect 13955 10013 13964 10047
rect 13912 10004 13964 10013
rect 14832 10004 14884 10056
rect 16304 10072 16356 10124
rect 17500 10072 17552 10124
rect 13820 9936 13872 9988
rect 14188 9936 14240 9988
rect 8300 9868 8352 9920
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 11980 9868 12032 9920
rect 15292 9911 15344 9920
rect 15292 9877 15301 9911
rect 15301 9877 15335 9911
rect 15335 9877 15344 9911
rect 15292 9868 15344 9877
rect 17960 9868 18012 9920
rect 3947 9766 3999 9818
rect 4011 9766 4063 9818
rect 4075 9766 4127 9818
rect 4139 9766 4191 9818
rect 9878 9766 9930 9818
rect 9942 9766 9994 9818
rect 10006 9766 10058 9818
rect 10070 9766 10122 9818
rect 15808 9766 15860 9818
rect 15872 9766 15924 9818
rect 15936 9766 15988 9818
rect 16000 9766 16052 9818
rect 2044 9503 2096 9512
rect 2044 9469 2053 9503
rect 2053 9469 2087 9503
rect 2087 9469 2096 9503
rect 2044 9460 2096 9469
rect 3056 9460 3108 9512
rect 8300 9664 8352 9716
rect 8392 9664 8444 9716
rect 11428 9664 11480 9716
rect 11704 9664 11756 9716
rect 5080 9596 5132 9648
rect 5724 9639 5776 9648
rect 5724 9605 5733 9639
rect 5733 9605 5767 9639
rect 5767 9605 5776 9639
rect 5724 9596 5776 9605
rect 5172 9528 5224 9580
rect 6276 9528 6328 9580
rect 8024 9596 8076 9648
rect 9312 9639 9364 9648
rect 7288 9571 7340 9580
rect 7288 9537 7297 9571
rect 7297 9537 7331 9571
rect 7331 9537 7340 9571
rect 7288 9528 7340 9537
rect 7472 9571 7524 9580
rect 7472 9537 7481 9571
rect 7481 9537 7515 9571
rect 7515 9537 7524 9571
rect 8208 9571 8260 9580
rect 7472 9528 7524 9537
rect 8208 9537 8217 9571
rect 8217 9537 8251 9571
rect 8251 9537 8260 9571
rect 8208 9528 8260 9537
rect 9312 9605 9321 9639
rect 9321 9605 9355 9639
rect 9355 9605 9364 9639
rect 9312 9596 9364 9605
rect 9496 9528 9548 9580
rect 10232 9596 10284 9648
rect 14188 9664 14240 9716
rect 16304 9664 16356 9716
rect 5448 9460 5500 9512
rect 5724 9460 5776 9512
rect 7564 9460 7616 9512
rect 8392 9460 8444 9512
rect 8668 9460 8720 9512
rect 8944 9503 8996 9512
rect 8944 9469 8953 9503
rect 8953 9469 8987 9503
rect 8987 9469 8996 9503
rect 8944 9460 8996 9469
rect 9128 9460 9180 9512
rect 13912 9596 13964 9648
rect 10692 9571 10744 9580
rect 10692 9537 10701 9571
rect 10701 9537 10735 9571
rect 10735 9537 10744 9571
rect 10692 9528 10744 9537
rect 11704 9528 11756 9580
rect 2504 9392 2556 9444
rect 4344 9392 4396 9444
rect 5264 9392 5316 9444
rect 3056 9324 3108 9376
rect 3516 9324 3568 9376
rect 4804 9324 4856 9376
rect 5632 9324 5684 9376
rect 7288 9324 7340 9376
rect 7932 9392 7984 9444
rect 8024 9324 8076 9376
rect 8392 9324 8444 9376
rect 9864 9392 9916 9444
rect 10416 9392 10468 9444
rect 9496 9324 9548 9376
rect 10876 9324 10928 9376
rect 12348 9460 12400 9512
rect 17684 9528 17736 9580
rect 11888 9392 11940 9444
rect 12256 9392 12308 9444
rect 12716 9435 12768 9444
rect 12716 9401 12750 9435
rect 12750 9401 12768 9435
rect 12716 9392 12768 9401
rect 14832 9460 14884 9512
rect 15016 9460 15068 9512
rect 15660 9392 15712 9444
rect 16120 9392 16172 9444
rect 18144 9392 18196 9444
rect 11336 9367 11388 9376
rect 11336 9333 11345 9367
rect 11345 9333 11379 9367
rect 11379 9333 11388 9367
rect 11336 9324 11388 9333
rect 12440 9324 12492 9376
rect 14832 9324 14884 9376
rect 16672 9324 16724 9376
rect 16856 9367 16908 9376
rect 16856 9333 16865 9367
rect 16865 9333 16899 9367
rect 16899 9333 16908 9367
rect 16856 9324 16908 9333
rect 6912 9222 6964 9274
rect 6976 9222 7028 9274
rect 7040 9222 7092 9274
rect 7104 9222 7156 9274
rect 12843 9222 12895 9274
rect 12907 9222 12959 9274
rect 12971 9222 13023 9274
rect 13035 9222 13087 9274
rect 2504 9052 2556 9104
rect 4068 9052 4120 9104
rect 4712 9052 4764 9104
rect 5264 9052 5316 9104
rect 5908 9052 5960 9104
rect 7472 9120 7524 9172
rect 8208 9120 8260 9172
rect 2320 9027 2372 9036
rect 2320 8993 2329 9027
rect 2329 8993 2363 9027
rect 2363 8993 2372 9027
rect 2320 8984 2372 8993
rect 2780 8984 2832 9036
rect 7564 9052 7616 9104
rect 8024 9052 8076 9104
rect 3424 8959 3476 8968
rect 1952 8823 2004 8832
rect 1952 8789 1961 8823
rect 1961 8789 1995 8823
rect 1995 8789 2004 8823
rect 1952 8780 2004 8789
rect 2412 8848 2464 8900
rect 3424 8925 3433 8959
rect 3433 8925 3467 8959
rect 3467 8925 3476 8959
rect 3424 8916 3476 8925
rect 3516 8959 3568 8968
rect 3516 8925 3525 8959
rect 3525 8925 3559 8959
rect 3559 8925 3568 8959
rect 3516 8916 3568 8925
rect 8484 8984 8536 9036
rect 9588 8984 9640 9036
rect 10048 8984 10100 9036
rect 11152 9052 11204 9104
rect 10692 8984 10744 9036
rect 10876 9027 10928 9036
rect 10876 8993 10885 9027
rect 10885 8993 10919 9027
rect 10919 8993 10928 9027
rect 10876 8984 10928 8993
rect 11336 9120 11388 9172
rect 11888 9120 11940 9172
rect 12532 9052 12584 9104
rect 15292 9120 15344 9172
rect 16304 9120 16356 9172
rect 17500 9163 17552 9172
rect 17500 9129 17509 9163
rect 17509 9129 17543 9163
rect 17543 9129 17552 9163
rect 17500 9120 17552 9129
rect 10324 8959 10376 8968
rect 2596 8848 2648 8900
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 10416 8916 10468 8968
rect 11152 8959 11204 8968
rect 11152 8925 11161 8959
rect 11161 8925 11195 8959
rect 11195 8925 11204 8959
rect 11152 8916 11204 8925
rect 12072 8916 12124 8968
rect 12348 8916 12400 8968
rect 15016 9052 15068 9104
rect 14004 8984 14056 9036
rect 14188 8984 14240 9036
rect 16120 9027 16172 9036
rect 16120 8993 16129 9027
rect 16129 8993 16163 9027
rect 16163 8993 16172 9027
rect 16120 8984 16172 8993
rect 17132 8984 17184 9036
rect 13360 8959 13412 8968
rect 2872 8780 2924 8832
rect 3516 8780 3568 8832
rect 7380 8848 7432 8900
rect 9864 8848 9916 8900
rect 10508 8891 10560 8900
rect 10508 8857 10517 8891
rect 10517 8857 10551 8891
rect 10551 8857 10560 8891
rect 10508 8848 10560 8857
rect 11612 8848 11664 8900
rect 12716 8848 12768 8900
rect 13360 8925 13369 8959
rect 13369 8925 13403 8959
rect 13403 8925 13412 8959
rect 13360 8916 13412 8925
rect 14832 8959 14884 8968
rect 14832 8925 14841 8959
rect 14841 8925 14875 8959
rect 14875 8925 14884 8959
rect 14832 8916 14884 8925
rect 15292 8959 15344 8968
rect 15292 8925 15301 8959
rect 15301 8925 15335 8959
rect 15335 8925 15344 8959
rect 15292 8916 15344 8925
rect 4436 8780 4488 8832
rect 4712 8780 4764 8832
rect 5632 8780 5684 8832
rect 9404 8780 9456 8832
rect 13912 8780 13964 8832
rect 14004 8780 14056 8832
rect 14924 8848 14976 8900
rect 15568 8848 15620 8900
rect 15200 8780 15252 8832
rect 16488 8780 16540 8832
rect 3947 8678 3999 8730
rect 4011 8678 4063 8730
rect 4075 8678 4127 8730
rect 4139 8678 4191 8730
rect 9878 8678 9930 8730
rect 9942 8678 9994 8730
rect 10006 8678 10058 8730
rect 10070 8678 10122 8730
rect 15808 8678 15860 8730
rect 15872 8678 15924 8730
rect 15936 8678 15988 8730
rect 16000 8678 16052 8730
rect 2044 8576 2096 8628
rect 2596 8576 2648 8628
rect 5908 8576 5960 8628
rect 2412 8508 2464 8560
rect 2504 8440 2556 8492
rect 3332 8508 3384 8560
rect 6644 8508 6696 8560
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 4712 8440 4764 8492
rect 3700 8304 3752 8356
rect 4436 8372 4488 8424
rect 10876 8576 10928 8628
rect 12440 8619 12492 8628
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 12440 8576 12492 8585
rect 9220 8508 9272 8560
rect 9588 8508 9640 8560
rect 10324 8508 10376 8560
rect 13268 8508 13320 8560
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 12716 8440 12768 8492
rect 14004 8483 14056 8492
rect 7656 8372 7708 8424
rect 11060 8372 11112 8424
rect 13452 8372 13504 8424
rect 5172 8347 5224 8356
rect 5172 8313 5206 8347
rect 5206 8313 5224 8347
rect 5172 8304 5224 8313
rect 8116 8304 8168 8356
rect 9496 8304 9548 8356
rect 11612 8347 11664 8356
rect 2964 8236 3016 8288
rect 3516 8236 3568 8288
rect 6736 8236 6788 8288
rect 7564 8236 7616 8288
rect 8760 8236 8812 8288
rect 11612 8313 11621 8347
rect 11621 8313 11655 8347
rect 11655 8313 11664 8347
rect 11612 8304 11664 8313
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14004 8440 14056 8449
rect 15568 8508 15620 8560
rect 14832 8440 14884 8492
rect 16120 8576 16172 8628
rect 16212 8576 16264 8628
rect 17132 8576 17184 8628
rect 17868 8508 17920 8560
rect 12256 8236 12308 8288
rect 13544 8236 13596 8288
rect 15108 8304 15160 8356
rect 17132 8372 17184 8424
rect 18052 8415 18104 8424
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 16488 8304 16540 8356
rect 14924 8279 14976 8288
rect 14924 8245 14933 8279
rect 14933 8245 14967 8279
rect 14967 8245 14976 8279
rect 14924 8236 14976 8245
rect 6912 8134 6964 8186
rect 6976 8134 7028 8186
rect 7040 8134 7092 8186
rect 7104 8134 7156 8186
rect 12843 8134 12895 8186
rect 12907 8134 12959 8186
rect 12971 8134 13023 8186
rect 13035 8134 13087 8186
rect 4620 8032 4672 8084
rect 5356 8032 5408 8084
rect 2964 7964 3016 8016
rect 3608 7964 3660 8016
rect 8576 8032 8628 8084
rect 8852 8032 8904 8084
rect 12716 8075 12768 8084
rect 7380 7964 7432 8016
rect 9680 7964 9732 8016
rect 10048 8007 10100 8016
rect 10048 7973 10057 8007
rect 10057 7973 10091 8007
rect 10091 7973 10100 8007
rect 10048 7964 10100 7973
rect 10416 7964 10468 8016
rect 10692 7964 10744 8016
rect 11704 7964 11756 8016
rect 2228 7939 2280 7948
rect 2228 7905 2237 7939
rect 2237 7905 2271 7939
rect 2271 7905 2280 7939
rect 2228 7896 2280 7905
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 2320 7760 2372 7812
rect 3240 7760 3292 7812
rect 6092 7896 6144 7948
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 6552 7828 6604 7837
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 9772 7896 9824 7948
rect 9864 7896 9916 7948
rect 10140 7939 10192 7948
rect 10140 7905 10149 7939
rect 10149 7905 10183 7939
rect 10183 7905 10192 7939
rect 10140 7896 10192 7905
rect 10324 7896 10376 7948
rect 12716 8041 12725 8075
rect 12725 8041 12759 8075
rect 12759 8041 12768 8075
rect 12716 8032 12768 8041
rect 13360 8075 13412 8084
rect 13360 8041 13369 8075
rect 13369 8041 13403 8075
rect 13403 8041 13412 8075
rect 13360 8032 13412 8041
rect 14372 8032 14424 8084
rect 16488 8032 16540 8084
rect 16856 8032 16908 8084
rect 17316 8075 17368 8084
rect 17316 8041 17325 8075
rect 17325 8041 17359 8075
rect 17359 8041 17368 8075
rect 17316 8032 17368 8041
rect 13912 7964 13964 8016
rect 13360 7896 13412 7948
rect 8208 7871 8260 7880
rect 7104 7760 7156 7812
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 8944 7828 8996 7880
rect 10692 7871 10744 7880
rect 10692 7837 10701 7871
rect 10701 7837 10735 7871
rect 10735 7837 10744 7871
rect 10692 7828 10744 7837
rect 13636 7896 13688 7948
rect 1860 7735 1912 7744
rect 1860 7701 1869 7735
rect 1869 7701 1903 7735
rect 1903 7701 1912 7735
rect 1860 7692 1912 7701
rect 3792 7692 3844 7744
rect 8024 7692 8076 7744
rect 8208 7692 8260 7744
rect 8300 7692 8352 7744
rect 14832 7871 14884 7880
rect 13176 7760 13228 7812
rect 14832 7837 14841 7871
rect 14841 7837 14875 7871
rect 14875 7837 14884 7871
rect 14832 7828 14884 7837
rect 13636 7760 13688 7812
rect 17132 7828 17184 7880
rect 17500 7871 17552 7880
rect 17500 7837 17509 7871
rect 17509 7837 17543 7871
rect 17543 7837 17552 7871
rect 17500 7828 17552 7837
rect 18144 7803 18196 7812
rect 18144 7769 18153 7803
rect 18153 7769 18187 7803
rect 18187 7769 18196 7803
rect 18144 7760 18196 7769
rect 13820 7692 13872 7744
rect 15660 7692 15712 7744
rect 3947 7590 3999 7642
rect 4011 7590 4063 7642
rect 4075 7590 4127 7642
rect 4139 7590 4191 7642
rect 9878 7590 9930 7642
rect 9942 7590 9994 7642
rect 10006 7590 10058 7642
rect 10070 7590 10122 7642
rect 15808 7590 15860 7642
rect 15872 7590 15924 7642
rect 15936 7590 15988 7642
rect 16000 7590 16052 7642
rect 2228 7488 2280 7540
rect 5172 7488 5224 7540
rect 7104 7531 7156 7540
rect 7104 7497 7113 7531
rect 7113 7497 7147 7531
rect 7147 7497 7156 7531
rect 7104 7488 7156 7497
rect 11704 7531 11756 7540
rect 6184 7420 6236 7472
rect 11704 7497 11713 7531
rect 11713 7497 11747 7531
rect 11747 7497 11756 7531
rect 11704 7488 11756 7497
rect 12164 7488 12216 7540
rect 12348 7488 12400 7540
rect 16396 7488 16448 7540
rect 16764 7488 16816 7540
rect 13452 7463 13504 7472
rect 13452 7429 13461 7463
rect 13461 7429 13495 7463
rect 13495 7429 13504 7463
rect 13452 7420 13504 7429
rect 18236 7463 18288 7472
rect 2688 7352 2740 7404
rect 3148 7352 3200 7404
rect 4712 7352 4764 7404
rect 4804 7352 4856 7404
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 10324 7395 10376 7404
rect 10324 7361 10333 7395
rect 10333 7361 10367 7395
rect 10367 7361 10376 7395
rect 10324 7352 10376 7361
rect 11336 7352 11388 7404
rect 11796 7352 11848 7404
rect 13176 7352 13228 7404
rect 2412 7284 2464 7336
rect 3700 7284 3752 7336
rect 2320 7216 2372 7268
rect 6644 7284 6696 7336
rect 7196 7284 7248 7336
rect 7748 7284 7800 7336
rect 8484 7327 8536 7336
rect 8484 7293 8493 7327
rect 8493 7293 8527 7327
rect 8527 7293 8536 7327
rect 8484 7284 8536 7293
rect 8760 7327 8812 7336
rect 8760 7293 8794 7327
rect 8794 7293 8812 7327
rect 8760 7284 8812 7293
rect 10232 7284 10284 7336
rect 10876 7284 10928 7336
rect 12256 7284 12308 7336
rect 18236 7429 18245 7463
rect 18245 7429 18279 7463
rect 18279 7429 18288 7463
rect 18236 7420 18288 7429
rect 2964 7191 3016 7200
rect 2964 7157 2973 7191
rect 2973 7157 3007 7191
rect 3007 7157 3016 7191
rect 2964 7148 3016 7157
rect 4712 7191 4764 7200
rect 4712 7157 4721 7191
rect 4721 7157 4755 7191
rect 4755 7157 4764 7191
rect 4712 7148 4764 7157
rect 5724 7216 5776 7268
rect 8944 7216 8996 7268
rect 9680 7216 9732 7268
rect 14832 7352 14884 7404
rect 15660 7352 15712 7404
rect 16488 7352 16540 7404
rect 16672 7352 16724 7404
rect 17592 7352 17644 7404
rect 15292 7284 15344 7336
rect 16948 7327 17000 7336
rect 16948 7293 16957 7327
rect 16957 7293 16991 7327
rect 16991 7293 17000 7327
rect 16948 7284 17000 7293
rect 17960 7284 18012 7336
rect 13820 7259 13872 7268
rect 6184 7148 6236 7200
rect 7564 7148 7616 7200
rect 7748 7148 7800 7200
rect 9404 7148 9456 7200
rect 10508 7148 10560 7200
rect 13820 7225 13829 7259
rect 13829 7225 13863 7259
rect 13863 7225 13872 7259
rect 13820 7216 13872 7225
rect 14096 7148 14148 7200
rect 14648 7148 14700 7200
rect 15660 7148 15712 7200
rect 6912 7046 6964 7098
rect 6976 7046 7028 7098
rect 7040 7046 7092 7098
rect 7104 7046 7156 7098
rect 12843 7046 12895 7098
rect 12907 7046 12959 7098
rect 12971 7046 13023 7098
rect 13035 7046 13087 7098
rect 2320 6944 2372 6996
rect 4804 6944 4856 6996
rect 6552 6944 6604 6996
rect 8024 6944 8076 6996
rect 8944 6944 8996 6996
rect 9588 6944 9640 6996
rect 10140 6944 10192 6996
rect 13176 6944 13228 6996
rect 15660 6987 15712 6996
rect 15660 6953 15669 6987
rect 15669 6953 15703 6987
rect 15703 6953 15712 6987
rect 15660 6944 15712 6953
rect 3976 6876 4028 6928
rect 4620 6876 4672 6928
rect 2320 6851 2372 6860
rect 2320 6817 2329 6851
rect 2329 6817 2363 6851
rect 2363 6817 2372 6851
rect 2320 6808 2372 6817
rect 2964 6808 3016 6860
rect 5264 6808 5316 6860
rect 8852 6876 8904 6928
rect 7104 6808 7156 6860
rect 7472 6808 7524 6860
rect 7656 6851 7708 6860
rect 7656 6817 7690 6851
rect 7690 6817 7708 6851
rect 7656 6808 7708 6817
rect 8208 6808 8260 6860
rect 10324 6876 10376 6928
rect 10692 6876 10744 6928
rect 11704 6808 11756 6860
rect 11888 6851 11940 6860
rect 11888 6817 11897 6851
rect 11897 6817 11931 6851
rect 11931 6817 11940 6851
rect 11888 6808 11940 6817
rect 12072 6808 12124 6860
rect 12900 6851 12952 6860
rect 6552 6740 6604 6792
rect 5080 6672 5132 6724
rect 1400 6604 1452 6656
rect 4344 6604 4396 6656
rect 9680 6740 9732 6792
rect 11612 6672 11664 6724
rect 12256 6740 12308 6792
rect 8576 6604 8628 6656
rect 12256 6604 12308 6656
rect 12900 6817 12909 6851
rect 12909 6817 12943 6851
rect 12943 6817 12952 6851
rect 12900 6808 12952 6817
rect 13452 6808 13504 6860
rect 13820 6851 13872 6860
rect 13820 6817 13854 6851
rect 13854 6817 13872 6851
rect 13820 6808 13872 6817
rect 14096 6808 14148 6860
rect 12992 6783 13044 6792
rect 12992 6749 13001 6783
rect 13001 6749 13035 6783
rect 13035 6749 13044 6783
rect 12992 6740 13044 6749
rect 13084 6740 13136 6792
rect 15568 6808 15620 6860
rect 16212 6740 16264 6792
rect 16580 6740 16632 6792
rect 18052 6715 18104 6724
rect 18052 6681 18061 6715
rect 18061 6681 18095 6715
rect 18095 6681 18104 6715
rect 18052 6672 18104 6681
rect 15292 6647 15344 6656
rect 15292 6613 15301 6647
rect 15301 6613 15335 6647
rect 15335 6613 15344 6647
rect 15292 6604 15344 6613
rect 16304 6647 16356 6656
rect 16304 6613 16313 6647
rect 16313 6613 16347 6647
rect 16347 6613 16356 6647
rect 16304 6604 16356 6613
rect 3947 6502 3999 6554
rect 4011 6502 4063 6554
rect 4075 6502 4127 6554
rect 4139 6502 4191 6554
rect 9878 6502 9930 6554
rect 9942 6502 9994 6554
rect 10006 6502 10058 6554
rect 10070 6502 10122 6554
rect 15808 6502 15860 6554
rect 15872 6502 15924 6554
rect 15936 6502 15988 6554
rect 16000 6502 16052 6554
rect 2688 6400 2740 6452
rect 4528 6400 4580 6452
rect 7104 6400 7156 6452
rect 8208 6443 8260 6452
rect 4068 6332 4120 6384
rect 4436 6332 4488 6384
rect 1952 6264 2004 6316
rect 2964 6264 3016 6316
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 4344 6264 4396 6273
rect 5264 6307 5316 6316
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 8208 6409 8217 6443
rect 8217 6409 8251 6443
rect 8251 6409 8260 6443
rect 8208 6400 8260 6409
rect 8300 6400 8352 6452
rect 10324 6400 10376 6452
rect 11888 6400 11940 6452
rect 11244 6332 11296 6384
rect 11796 6332 11848 6384
rect 12716 6400 12768 6452
rect 12900 6400 12952 6452
rect 13728 6400 13780 6452
rect 15660 6400 15712 6452
rect 18236 6443 18288 6452
rect 18236 6409 18245 6443
rect 18245 6409 18279 6443
rect 18279 6409 18288 6443
rect 18236 6400 18288 6409
rect 12624 6332 12676 6384
rect 12992 6332 13044 6384
rect 15936 6332 15988 6384
rect 17960 6332 18012 6384
rect 1860 6196 1912 6248
rect 4988 6196 5040 6248
rect 5448 6196 5500 6248
rect 7472 6196 7524 6248
rect 8484 6196 8536 6248
rect 11336 6264 11388 6316
rect 11704 6264 11756 6316
rect 13084 6264 13136 6316
rect 13544 6264 13596 6316
rect 13820 6264 13872 6316
rect 15108 6307 15160 6316
rect 10968 6239 11020 6248
rect 10968 6205 10977 6239
rect 10977 6205 11011 6239
rect 11011 6205 11020 6239
rect 10968 6196 11020 6205
rect 2964 6128 3016 6180
rect 3608 6128 3660 6180
rect 5908 6128 5960 6180
rect 6736 6128 6788 6180
rect 9404 6171 9456 6180
rect 2320 6060 2372 6112
rect 3700 6103 3752 6112
rect 3700 6069 3709 6103
rect 3709 6069 3743 6103
rect 3743 6069 3752 6103
rect 3700 6060 3752 6069
rect 4896 6060 4948 6112
rect 5264 6060 5316 6112
rect 6092 6103 6144 6112
rect 6092 6069 6101 6103
rect 6101 6069 6135 6103
rect 6135 6069 6144 6103
rect 6092 6060 6144 6069
rect 7288 6060 7340 6112
rect 9404 6137 9438 6171
rect 9438 6137 9456 6171
rect 9404 6128 9456 6137
rect 12624 6196 12676 6248
rect 13728 6196 13780 6248
rect 13912 6239 13964 6248
rect 13912 6205 13921 6239
rect 13921 6205 13955 6239
rect 13955 6205 13964 6239
rect 13912 6196 13964 6205
rect 15108 6273 15117 6307
rect 15117 6273 15151 6307
rect 15151 6273 15160 6307
rect 15108 6264 15160 6273
rect 17040 6196 17092 6248
rect 17776 6196 17828 6248
rect 11520 6128 11572 6180
rect 17316 6128 17368 6180
rect 11612 6060 11664 6112
rect 12716 6060 12768 6112
rect 13360 6060 13412 6112
rect 13820 6060 13872 6112
rect 13912 6060 13964 6112
rect 14188 6060 14240 6112
rect 14556 6103 14608 6112
rect 14556 6069 14565 6103
rect 14565 6069 14599 6103
rect 14599 6069 14608 6103
rect 14556 6060 14608 6069
rect 14924 6103 14976 6112
rect 14924 6069 14933 6103
rect 14933 6069 14967 6103
rect 14967 6069 14976 6103
rect 14924 6060 14976 6069
rect 15476 6060 15528 6112
rect 15936 6103 15988 6112
rect 15936 6069 15945 6103
rect 15945 6069 15979 6103
rect 15979 6069 15988 6103
rect 15936 6060 15988 6069
rect 16396 6060 16448 6112
rect 17592 6103 17644 6112
rect 17592 6069 17601 6103
rect 17601 6069 17635 6103
rect 17635 6069 17644 6103
rect 17592 6060 17644 6069
rect 6912 5958 6964 6010
rect 6976 5958 7028 6010
rect 7040 5958 7092 6010
rect 7104 5958 7156 6010
rect 12843 5958 12895 6010
rect 12907 5958 12959 6010
rect 12971 5958 13023 6010
rect 13035 5958 13087 6010
rect 6092 5856 6144 5908
rect 6736 5856 6788 5908
rect 8024 5856 8076 5908
rect 10968 5856 11020 5908
rect 4344 5788 4396 5840
rect 2688 5720 2740 5772
rect 3240 5763 3292 5772
rect 3240 5729 3249 5763
rect 3249 5729 3283 5763
rect 3283 5729 3292 5763
rect 3240 5720 3292 5729
rect 4160 5720 4212 5772
rect 1492 5652 1544 5704
rect 4068 5652 4120 5704
rect 5172 5788 5224 5840
rect 4712 5720 4764 5772
rect 5448 5763 5500 5772
rect 5448 5729 5457 5763
rect 5457 5729 5491 5763
rect 5491 5729 5500 5763
rect 5448 5720 5500 5729
rect 7104 5763 7156 5772
rect 7104 5729 7113 5763
rect 7113 5729 7147 5763
rect 7147 5729 7156 5763
rect 7104 5720 7156 5729
rect 9312 5720 9364 5772
rect 10324 5788 10376 5840
rect 11244 5720 11296 5772
rect 12164 5788 12216 5840
rect 13728 5720 13780 5772
rect 14924 5856 14976 5908
rect 18052 5899 18104 5908
rect 18052 5865 18061 5899
rect 18061 5865 18095 5899
rect 18095 5865 18104 5899
rect 18052 5856 18104 5865
rect 14096 5788 14148 5840
rect 14648 5831 14700 5840
rect 14648 5797 14657 5831
rect 14657 5797 14691 5831
rect 14691 5797 14700 5831
rect 14648 5788 14700 5797
rect 17316 5763 17368 5772
rect 17316 5729 17325 5763
rect 17325 5729 17359 5763
rect 17359 5729 17368 5763
rect 17316 5720 17368 5729
rect 4344 5584 4396 5636
rect 4988 5652 5040 5704
rect 5356 5652 5408 5704
rect 3148 5516 3200 5568
rect 3424 5559 3476 5568
rect 3424 5525 3433 5559
rect 3433 5525 3467 5559
rect 3467 5525 3476 5559
rect 3424 5516 3476 5525
rect 3792 5516 3844 5568
rect 4804 5516 4856 5568
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 15016 5652 15068 5704
rect 13544 5627 13596 5636
rect 13544 5593 13553 5627
rect 13553 5593 13587 5627
rect 13587 5593 13596 5627
rect 13544 5584 13596 5593
rect 13636 5584 13688 5636
rect 7472 5516 7524 5568
rect 7748 5516 7800 5568
rect 11336 5559 11388 5568
rect 11336 5525 11345 5559
rect 11345 5525 11379 5559
rect 11379 5525 11388 5559
rect 11336 5516 11388 5525
rect 12164 5516 12216 5568
rect 12440 5516 12492 5568
rect 13452 5516 13504 5568
rect 17500 5559 17552 5568
rect 17500 5525 17509 5559
rect 17509 5525 17543 5559
rect 17543 5525 17552 5559
rect 17500 5516 17552 5525
rect 3947 5414 3999 5466
rect 4011 5414 4063 5466
rect 4075 5414 4127 5466
rect 4139 5414 4191 5466
rect 9878 5414 9930 5466
rect 9942 5414 9994 5466
rect 10006 5414 10058 5466
rect 10070 5414 10122 5466
rect 15808 5414 15860 5466
rect 15872 5414 15924 5466
rect 15936 5414 15988 5466
rect 16000 5414 16052 5466
rect 3700 5312 3752 5364
rect 4988 5312 5040 5364
rect 5080 5312 5132 5364
rect 6368 5312 6420 5364
rect 8852 5355 8904 5364
rect 4344 5176 4396 5228
rect 1492 5108 1544 5160
rect 2044 5108 2096 5160
rect 5356 5151 5408 5160
rect 3148 5040 3200 5092
rect 5356 5117 5365 5151
rect 5365 5117 5399 5151
rect 5399 5117 5408 5151
rect 5356 5108 5408 5117
rect 7104 5176 7156 5228
rect 8852 5321 8861 5355
rect 8861 5321 8895 5355
rect 8895 5321 8904 5355
rect 8852 5312 8904 5321
rect 7472 5244 7524 5296
rect 9588 5312 9640 5364
rect 9772 5312 9824 5364
rect 10508 5312 10560 5364
rect 11152 5312 11204 5364
rect 9220 5244 9272 5296
rect 12256 5244 12308 5296
rect 13728 5312 13780 5364
rect 14096 5312 14148 5364
rect 14832 5312 14884 5364
rect 15476 5312 15528 5364
rect 7656 5176 7708 5228
rect 8300 5219 8352 5228
rect 8300 5185 8309 5219
rect 8309 5185 8343 5219
rect 8343 5185 8352 5219
rect 8300 5176 8352 5185
rect 8668 5176 8720 5228
rect 9312 5176 9364 5228
rect 12440 5219 12492 5228
rect 12440 5185 12449 5219
rect 12449 5185 12483 5219
rect 12483 5185 12492 5219
rect 12440 5176 12492 5185
rect 13452 5176 13504 5228
rect 15936 5176 15988 5228
rect 6276 5108 6328 5160
rect 4528 5040 4580 5092
rect 2780 5015 2832 5024
rect 2780 4981 2789 5015
rect 2789 4981 2823 5015
rect 2823 4981 2832 5015
rect 3240 5015 3292 5024
rect 2780 4972 2832 4981
rect 3240 4981 3249 5015
rect 3249 4981 3283 5015
rect 3283 4981 3292 5015
rect 3240 4972 3292 4981
rect 4344 5015 4396 5024
rect 4344 4981 4353 5015
rect 4353 4981 4387 5015
rect 4387 4981 4396 5015
rect 4344 4972 4396 4981
rect 4436 5015 4488 5024
rect 4436 4981 4445 5015
rect 4445 4981 4479 5015
rect 4479 4981 4488 5015
rect 4436 4972 4488 4981
rect 5172 4972 5224 5024
rect 9680 5108 9732 5160
rect 11520 5108 11572 5160
rect 13636 5108 13688 5160
rect 13820 5108 13872 5160
rect 14832 5108 14884 5160
rect 18328 5108 18380 5160
rect 11152 5040 11204 5092
rect 14372 5083 14424 5092
rect 14372 5049 14406 5083
rect 14406 5049 14424 5083
rect 16120 5083 16172 5092
rect 8208 5015 8260 5024
rect 8208 4981 8217 5015
rect 8217 4981 8251 5015
rect 8251 4981 8260 5015
rect 8208 4972 8260 4981
rect 9220 5015 9272 5024
rect 9220 4981 9229 5015
rect 9229 4981 9263 5015
rect 9263 4981 9272 5015
rect 9220 4972 9272 4981
rect 9680 4972 9732 5024
rect 10140 4972 10192 5024
rect 10416 4972 10468 5024
rect 11796 4972 11848 5024
rect 14372 5040 14424 5049
rect 16120 5049 16129 5083
rect 16129 5049 16163 5083
rect 16163 5049 16172 5083
rect 16120 5040 16172 5049
rect 17776 5040 17828 5092
rect 13360 4972 13412 5024
rect 15108 4972 15160 5024
rect 16212 5015 16264 5024
rect 16212 4981 16221 5015
rect 16221 4981 16255 5015
rect 16255 4981 16264 5015
rect 16212 4972 16264 4981
rect 17592 5015 17644 5024
rect 17592 4981 17601 5015
rect 17601 4981 17635 5015
rect 17635 4981 17644 5015
rect 17592 4972 17644 4981
rect 18236 5015 18288 5024
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 6912 4870 6964 4922
rect 6976 4870 7028 4922
rect 7040 4870 7092 4922
rect 7104 4870 7156 4922
rect 12843 4870 12895 4922
rect 12907 4870 12959 4922
rect 12971 4870 13023 4922
rect 13035 4870 13087 4922
rect 2412 4700 2464 4752
rect 2780 4700 2832 4752
rect 2044 4607 2096 4616
rect 2044 4573 2053 4607
rect 2053 4573 2087 4607
rect 2087 4573 2096 4607
rect 2044 4564 2096 4573
rect 4068 4768 4120 4820
rect 4804 4768 4856 4820
rect 7288 4768 7340 4820
rect 8300 4768 8352 4820
rect 8852 4768 8904 4820
rect 9312 4768 9364 4820
rect 11796 4811 11848 4820
rect 11796 4777 11805 4811
rect 11805 4777 11839 4811
rect 11839 4777 11848 4811
rect 11796 4768 11848 4777
rect 12348 4768 12400 4820
rect 14464 4768 14516 4820
rect 14924 4768 14976 4820
rect 15660 4811 15712 4820
rect 3148 4700 3200 4752
rect 6368 4700 6420 4752
rect 3792 4632 3844 4684
rect 4068 4675 4120 4684
rect 4068 4641 4077 4675
rect 4077 4641 4111 4675
rect 4111 4641 4120 4675
rect 4068 4632 4120 4641
rect 4344 4675 4396 4684
rect 4344 4641 4378 4675
rect 4378 4641 4396 4675
rect 4344 4632 4396 4641
rect 3332 4564 3384 4616
rect 3608 4564 3660 4616
rect 6184 4675 6236 4684
rect 6184 4641 6193 4675
rect 6193 4641 6227 4675
rect 6227 4641 6236 4675
rect 6184 4632 6236 4641
rect 6644 4632 6696 4684
rect 7472 4632 7524 4684
rect 7656 4632 7708 4684
rect 8668 4632 8720 4684
rect 1676 4471 1728 4480
rect 1676 4437 1685 4471
rect 1685 4437 1719 4471
rect 1719 4437 1728 4471
rect 1676 4428 1728 4437
rect 3700 4428 3752 4480
rect 5448 4471 5500 4480
rect 5448 4437 5457 4471
rect 5457 4437 5491 4471
rect 5491 4437 5500 4471
rect 5448 4428 5500 4437
rect 5724 4471 5776 4480
rect 5724 4437 5733 4471
rect 5733 4437 5767 4471
rect 5767 4437 5776 4471
rect 5724 4428 5776 4437
rect 6092 4496 6144 4548
rect 7748 4564 7800 4616
rect 10324 4700 10376 4752
rect 9864 4632 9916 4684
rect 11060 4700 11112 4752
rect 11336 4700 11388 4752
rect 15660 4777 15669 4811
rect 15669 4777 15703 4811
rect 15703 4777 15712 4811
rect 15660 4768 15712 4777
rect 16580 4700 16632 4752
rect 17316 4675 17368 4684
rect 8852 4496 8904 4548
rect 6736 4471 6788 4480
rect 6736 4437 6745 4471
rect 6745 4437 6779 4471
rect 6779 4437 6788 4471
rect 6736 4428 6788 4437
rect 6828 4428 6880 4480
rect 9680 4428 9732 4480
rect 17316 4641 17325 4675
rect 17325 4641 17359 4675
rect 17359 4641 17368 4675
rect 17316 4632 17368 4641
rect 11336 4564 11388 4616
rect 12532 4564 12584 4616
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 14188 4607 14240 4616
rect 14188 4573 14197 4607
rect 14197 4573 14231 4607
rect 14231 4573 14240 4607
rect 14188 4564 14240 4573
rect 14372 4607 14424 4616
rect 14372 4573 14381 4607
rect 14381 4573 14415 4607
rect 14415 4573 14424 4607
rect 14372 4564 14424 4573
rect 15200 4564 15252 4616
rect 15936 4607 15988 4616
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 15936 4564 15988 4573
rect 11612 4496 11664 4548
rect 13176 4496 13228 4548
rect 15016 4496 15068 4548
rect 11152 4471 11204 4480
rect 11152 4437 11161 4471
rect 11161 4437 11195 4471
rect 11195 4437 11204 4471
rect 11152 4428 11204 4437
rect 12532 4428 12584 4480
rect 12716 4471 12768 4480
rect 12716 4437 12725 4471
rect 12725 4437 12759 4471
rect 12759 4437 12768 4471
rect 12716 4428 12768 4437
rect 12808 4428 12860 4480
rect 17500 4471 17552 4480
rect 17500 4437 17509 4471
rect 17509 4437 17543 4471
rect 17543 4437 17552 4471
rect 17500 4428 17552 4437
rect 17868 4428 17920 4480
rect 3947 4326 3999 4378
rect 4011 4326 4063 4378
rect 4075 4326 4127 4378
rect 4139 4326 4191 4378
rect 9878 4326 9930 4378
rect 9942 4326 9994 4378
rect 10006 4326 10058 4378
rect 10070 4326 10122 4378
rect 15808 4326 15860 4378
rect 15872 4326 15924 4378
rect 15936 4326 15988 4378
rect 16000 4326 16052 4378
rect 2044 4224 2096 4276
rect 2412 4156 2464 4208
rect 3792 4224 3844 4276
rect 4344 4224 4396 4276
rect 4436 4224 4488 4276
rect 11612 4224 11664 4276
rect 13176 4224 13228 4276
rect 15016 4267 15068 4276
rect 7472 4156 7524 4208
rect 8208 4156 8260 4208
rect 5172 4088 5224 4140
rect 5448 4088 5500 4140
rect 4896 4020 4948 4072
rect 5632 4020 5684 4072
rect 3700 3952 3752 4004
rect 3792 3952 3844 4004
rect 1952 3884 2004 3936
rect 4252 3884 4304 3936
rect 5172 3952 5224 4004
rect 6000 4063 6052 4072
rect 6000 4029 6009 4063
rect 6009 4029 6043 4063
rect 6043 4029 6052 4063
rect 6000 4020 6052 4029
rect 6460 4020 6512 4072
rect 7564 4088 7616 4140
rect 8668 4088 8720 4140
rect 9312 4156 9364 4208
rect 10232 4131 10284 4140
rect 10232 4097 10241 4131
rect 10241 4097 10275 4131
rect 10275 4097 10284 4131
rect 10232 4088 10284 4097
rect 10324 4088 10376 4140
rect 12716 4088 12768 4140
rect 13636 4156 13688 4208
rect 15016 4233 15025 4267
rect 15025 4233 15059 4267
rect 15059 4233 15068 4267
rect 15016 4224 15068 4233
rect 16212 4224 16264 4276
rect 15660 4156 15712 4208
rect 15200 4088 15252 4140
rect 15568 4088 15620 4140
rect 7656 4020 7708 4072
rect 7932 4020 7984 4072
rect 10600 4020 10652 4072
rect 13452 4020 13504 4072
rect 5816 3952 5868 4004
rect 6552 3952 6604 4004
rect 4896 3884 4948 3936
rect 6736 3884 6788 3936
rect 8576 3884 8628 3936
rect 8760 3884 8812 3936
rect 9496 3884 9548 3936
rect 11152 3952 11204 4004
rect 16304 4020 16356 4072
rect 13912 3995 13964 4004
rect 13912 3961 13946 3995
rect 13946 3961 13964 3995
rect 13912 3952 13964 3961
rect 14832 3952 14884 4004
rect 12072 3927 12124 3936
rect 12072 3893 12081 3927
rect 12081 3893 12115 3927
rect 12115 3893 12124 3927
rect 12072 3884 12124 3893
rect 12716 3884 12768 3936
rect 14556 3884 14608 3936
rect 16672 3884 16724 3936
rect 17408 3884 17460 3936
rect 17592 3927 17644 3936
rect 17592 3893 17601 3927
rect 17601 3893 17635 3927
rect 17635 3893 17644 3927
rect 17592 3884 17644 3893
rect 18328 3884 18380 3936
rect 6912 3782 6964 3834
rect 6976 3782 7028 3834
rect 7040 3782 7092 3834
rect 7104 3782 7156 3834
rect 12843 3782 12895 3834
rect 12907 3782 12959 3834
rect 12971 3782 13023 3834
rect 13035 3782 13087 3834
rect 2780 3680 2832 3732
rect 4988 3680 5040 3732
rect 8392 3680 8444 3732
rect 10324 3680 10376 3732
rect 1584 3587 1636 3596
rect 1584 3553 1593 3587
rect 1593 3553 1627 3587
rect 1627 3553 1636 3587
rect 1584 3544 1636 3553
rect 5172 3612 5224 3664
rect 5448 3612 5500 3664
rect 10416 3612 10468 3664
rect 10508 3612 10560 3664
rect 14188 3680 14240 3732
rect 17132 3680 17184 3732
rect 12072 3612 12124 3664
rect 12716 3612 12768 3664
rect 3332 3587 3384 3596
rect 3332 3553 3341 3587
rect 3341 3553 3375 3587
rect 3375 3553 3384 3587
rect 3332 3544 3384 3553
rect 5540 3544 5592 3596
rect 1216 3476 1268 3528
rect 3148 3476 3200 3528
rect 4344 3476 4396 3528
rect 4804 3408 4856 3460
rect 4988 3340 5040 3392
rect 5172 3340 5224 3392
rect 9128 3544 9180 3596
rect 10784 3544 10836 3596
rect 11888 3544 11940 3596
rect 12348 3544 12400 3596
rect 14096 3544 14148 3596
rect 8484 3476 8536 3528
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 10416 3476 10468 3528
rect 10876 3476 10928 3528
rect 9772 3408 9824 3460
rect 11244 3476 11296 3528
rect 13268 3476 13320 3528
rect 15568 3544 15620 3596
rect 16580 3544 16632 3596
rect 7748 3340 7800 3392
rect 8668 3340 8720 3392
rect 9588 3340 9640 3392
rect 10600 3340 10652 3392
rect 12256 3408 12308 3460
rect 13912 3408 13964 3460
rect 11796 3340 11848 3392
rect 12072 3340 12124 3392
rect 17500 3383 17552 3392
rect 17500 3349 17509 3383
rect 17509 3349 17543 3383
rect 17543 3349 17552 3383
rect 17500 3340 17552 3349
rect 18052 3383 18104 3392
rect 18052 3349 18061 3383
rect 18061 3349 18095 3383
rect 18095 3349 18104 3383
rect 18052 3340 18104 3349
rect 3947 3238 3999 3290
rect 4011 3238 4063 3290
rect 4075 3238 4127 3290
rect 4139 3238 4191 3290
rect 9878 3238 9930 3290
rect 9942 3238 9994 3290
rect 10006 3238 10058 3290
rect 10070 3238 10122 3290
rect 15808 3238 15860 3290
rect 15872 3238 15924 3290
rect 15936 3238 15988 3290
rect 16000 3238 16052 3290
rect 3148 3179 3200 3188
rect 3148 3145 3157 3179
rect 3157 3145 3191 3179
rect 3191 3145 3200 3179
rect 3148 3136 3200 3145
rect 5540 3179 5592 3188
rect 5540 3145 5549 3179
rect 5549 3145 5583 3179
rect 5583 3145 5592 3179
rect 5540 3136 5592 3145
rect 8760 3136 8812 3188
rect 9128 3179 9180 3188
rect 9128 3145 9137 3179
rect 9137 3145 9171 3179
rect 9171 3145 9180 3179
rect 9128 3136 9180 3145
rect 11704 3136 11756 3188
rect 11796 3136 11848 3188
rect 15476 3136 15528 3188
rect 16396 3136 16448 3188
rect 5448 3068 5500 3120
rect 5908 3068 5960 3120
rect 9036 3068 9088 3120
rect 9404 3068 9456 3120
rect 2780 3000 2832 3052
rect 3700 3043 3752 3052
rect 3700 3009 3709 3043
rect 3709 3009 3743 3043
rect 3743 3009 3752 3043
rect 3700 3000 3752 3009
rect 4988 3043 5040 3052
rect 4988 3009 4997 3043
rect 4997 3009 5031 3043
rect 5031 3009 5040 3043
rect 4988 3000 5040 3009
rect 5172 3043 5224 3052
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 6092 3043 6144 3052
rect 6092 3009 6101 3043
rect 6101 3009 6135 3043
rect 6135 3009 6144 3043
rect 6092 3000 6144 3009
rect 8668 3043 8720 3052
rect 8668 3009 8677 3043
rect 8677 3009 8711 3043
rect 8711 3009 8720 3043
rect 8668 3000 8720 3009
rect 9588 3043 9640 3052
rect 9588 3009 9597 3043
rect 9597 3009 9631 3043
rect 9631 3009 9640 3043
rect 9588 3000 9640 3009
rect 11152 3068 11204 3120
rect 10600 3043 10652 3052
rect 10600 3009 10609 3043
rect 10609 3009 10643 3043
rect 10643 3009 10652 3043
rect 10600 3000 10652 3009
rect 11060 3000 11112 3052
rect 11612 3043 11664 3052
rect 11612 3009 11621 3043
rect 11621 3009 11655 3043
rect 11655 3009 11664 3043
rect 11612 3000 11664 3009
rect 11888 3068 11940 3120
rect 2320 2975 2372 2984
rect 2320 2941 2329 2975
rect 2329 2941 2363 2975
rect 2363 2941 2372 2975
rect 2320 2932 2372 2941
rect 2872 2932 2924 2984
rect 3608 2975 3660 2984
rect 3608 2941 3617 2975
rect 3617 2941 3651 2975
rect 3651 2941 3660 2975
rect 4896 2975 4948 2984
rect 3608 2932 3660 2941
rect 4896 2941 4905 2975
rect 4905 2941 4939 2975
rect 4939 2941 4948 2975
rect 4896 2932 4948 2941
rect 2136 2864 2188 2916
rect 9496 2975 9548 2984
rect 9496 2941 9505 2975
rect 9505 2941 9539 2975
rect 9539 2941 9548 2975
rect 9496 2932 9548 2941
rect 10692 2932 10744 2984
rect 13912 3000 13964 3052
rect 14648 2932 14700 2984
rect 5908 2839 5960 2848
rect 5908 2805 5917 2839
rect 5917 2805 5951 2839
rect 5951 2805 5960 2839
rect 5908 2796 5960 2805
rect 6000 2839 6052 2848
rect 6000 2805 6009 2839
rect 6009 2805 6043 2839
rect 6043 2805 6052 2839
rect 11244 2864 11296 2916
rect 11520 2907 11572 2916
rect 11520 2873 11529 2907
rect 11529 2873 11563 2907
rect 11563 2873 11572 2907
rect 11520 2864 11572 2873
rect 12532 2864 12584 2916
rect 14832 2864 14884 2916
rect 15568 2932 15620 2984
rect 16672 2932 16724 2984
rect 17684 3000 17736 3052
rect 17040 2932 17092 2984
rect 15200 2864 15252 2916
rect 6000 2796 6052 2805
rect 8116 2796 8168 2848
rect 8392 2796 8444 2848
rect 8576 2839 8628 2848
rect 8576 2805 8585 2839
rect 8585 2805 8619 2839
rect 8619 2805 8628 2839
rect 8576 2796 8628 2805
rect 8760 2796 8812 2848
rect 10876 2796 10928 2848
rect 16396 2839 16448 2848
rect 16396 2805 16405 2839
rect 16405 2805 16439 2839
rect 16439 2805 16448 2839
rect 16396 2796 16448 2805
rect 17040 2839 17092 2848
rect 17040 2805 17049 2839
rect 17049 2805 17083 2839
rect 17083 2805 17092 2839
rect 17040 2796 17092 2805
rect 17684 2796 17736 2848
rect 18236 2839 18288 2848
rect 18236 2805 18245 2839
rect 18245 2805 18279 2839
rect 18279 2805 18288 2839
rect 18236 2796 18288 2805
rect 6912 2694 6964 2746
rect 6976 2694 7028 2746
rect 7040 2694 7092 2746
rect 7104 2694 7156 2746
rect 12843 2694 12895 2746
rect 12907 2694 12959 2746
rect 12971 2694 13023 2746
rect 13035 2694 13087 2746
rect 1860 2635 1912 2644
rect 1860 2601 1869 2635
rect 1869 2601 1903 2635
rect 1903 2601 1912 2635
rect 1860 2592 1912 2601
rect 2688 2592 2740 2644
rect 3516 2592 3568 2644
rect 5172 2592 5224 2644
rect 9772 2592 9824 2644
rect 4252 2524 4304 2576
rect 6092 2524 6144 2576
rect 1952 2456 2004 2508
rect 4068 2456 4120 2508
rect 5448 2499 5500 2508
rect 5448 2465 5457 2499
rect 5457 2465 5491 2499
rect 5491 2465 5500 2499
rect 5448 2456 5500 2465
rect 7472 2524 7524 2576
rect 10968 2592 11020 2644
rect 11704 2635 11756 2644
rect 11704 2601 11713 2635
rect 11713 2601 11747 2635
rect 11747 2601 11756 2635
rect 11704 2592 11756 2601
rect 11888 2524 11940 2576
rect 7380 2456 7432 2508
rect 7840 2456 7892 2508
rect 10784 2456 10836 2508
rect 11428 2456 11480 2508
rect 15292 2524 15344 2576
rect 14188 2456 14240 2508
rect 14464 2456 14516 2508
rect 3056 2388 3108 2440
rect 3700 2388 3752 2440
rect 5632 2431 5684 2440
rect 5632 2397 5641 2431
rect 5641 2397 5675 2431
rect 5675 2397 5684 2431
rect 5632 2388 5684 2397
rect 3332 2320 3384 2372
rect 4896 2320 4948 2372
rect 7564 2388 7616 2440
rect 10324 2388 10376 2440
rect 11060 2388 11112 2440
rect 11152 2388 11204 2440
rect 13084 2388 13136 2440
rect 12164 2320 12216 2372
rect 6000 2252 6052 2304
rect 11428 2252 11480 2304
rect 17592 2295 17644 2304
rect 17592 2261 17601 2295
rect 17601 2261 17635 2295
rect 17635 2261 17644 2295
rect 17592 2252 17644 2261
rect 3947 2150 3999 2202
rect 4011 2150 4063 2202
rect 4075 2150 4127 2202
rect 4139 2150 4191 2202
rect 9878 2150 9930 2202
rect 9942 2150 9994 2202
rect 10006 2150 10058 2202
rect 10070 2150 10122 2202
rect 15808 2150 15860 2202
rect 15872 2150 15924 2202
rect 15936 2150 15988 2202
rect 16000 2150 16052 2202
rect 3700 2048 3752 2100
rect 5080 2048 5132 2100
rect 9404 2048 9456 2100
rect 11888 2048 11940 2100
rect 11244 1504 11296 1556
rect 19432 1504 19484 1556
rect 3976 1368 4028 1420
rect 5632 1368 5684 1420
rect 3332 1300 3384 1352
rect 12072 1300 12124 1352
rect 388 960 440 1012
rect 8760 960 8812 1012
<< metal2 >>
rect 1122 16520 1178 17000
rect 3330 16520 3386 17000
rect 4066 16688 4122 16697
rect 4066 16623 4122 16632
rect 1136 13326 1164 16520
rect 2870 15872 2926 15881
rect 2870 15807 2926 15816
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1124 13320 1176 13326
rect 1124 13262 1176 13268
rect 1780 12986 1808 13330
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1964 12170 1992 13670
rect 2700 13326 2728 13874
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2044 13252 2096 13258
rect 2044 13194 2096 13200
rect 2056 12850 2084 13194
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1952 12164 2004 12170
rect 1952 12106 2004 12112
rect 2056 11762 2084 12786
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 1400 11076 1452 11082
rect 1400 11018 1452 11024
rect 1412 7585 1440 11018
rect 2056 10538 2084 11086
rect 2044 10532 2096 10538
rect 2044 10474 2096 10480
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1398 7576 1454 7585
rect 1398 7511 1454 7520
rect 1400 6656 1452 6662
rect 1400 6598 1452 6604
rect 1412 4729 1440 6598
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1504 5166 1532 5646
rect 1492 5160 1544 5166
rect 1492 5102 1544 5108
rect 1398 4720 1454 4729
rect 1398 4655 1454 4664
rect 1596 3602 1624 9862
rect 2056 9518 2084 10474
rect 2148 10198 2176 12582
rect 2240 10266 2268 13126
rect 2318 12744 2374 12753
rect 2318 12679 2320 12688
rect 2372 12679 2374 12688
rect 2320 12650 2372 12656
rect 2332 11286 2360 12650
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2424 11898 2452 12174
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2608 11762 2636 12174
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2320 11280 2372 11286
rect 2320 11222 2372 11228
rect 2424 10606 2452 11290
rect 2608 11286 2636 11698
rect 2700 11354 2728 13262
rect 2792 11830 2820 13806
rect 2884 13530 2912 15807
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 2964 14000 3016 14006
rect 2964 13942 3016 13948
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2870 13424 2926 13433
rect 2870 13359 2926 13368
rect 2884 12102 2912 13359
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2780 11824 2832 11830
rect 2780 11766 2832 11772
rect 2872 11620 2924 11626
rect 2872 11562 2924 11568
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2596 11280 2648 11286
rect 2596 11222 2648 11228
rect 2608 11014 2636 11222
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2792 10810 2820 11494
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2136 10192 2188 10198
rect 2136 10134 2188 10140
rect 2516 10062 2544 10406
rect 2884 10266 2912 11562
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2976 10130 3004 13942
rect 3068 12442 3096 14350
rect 3344 14346 3372 16520
rect 3790 15464 3846 15473
rect 3790 15399 3846 15408
rect 3698 15056 3754 15065
rect 3698 14991 3754 15000
rect 3514 14648 3570 14657
rect 3424 14612 3476 14618
rect 3514 14583 3570 14592
rect 3424 14554 3476 14560
rect 3332 14340 3384 14346
rect 3332 14282 3384 14288
rect 3436 13841 3464 14554
rect 3422 13832 3478 13841
rect 3422 13767 3478 13776
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 3160 10554 3188 13330
rect 3528 12170 3556 14583
rect 3606 14240 3662 14249
rect 3606 14175 3662 14184
rect 3620 14006 3648 14175
rect 3608 14000 3660 14006
rect 3608 13942 3660 13948
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 3620 12238 3648 12650
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 3516 11620 3568 11626
rect 3516 11562 3568 11568
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 3068 10526 3188 10554
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1872 6254 1900 7686
rect 1964 6322 1992 8774
rect 2056 8634 2084 9454
rect 2516 9450 2544 9998
rect 2778 9752 2834 9761
rect 2778 9687 2834 9696
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 2792 9160 2820 9687
rect 3068 9518 3096 10526
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2792 9132 3004 9160
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 2240 7546 2268 7890
rect 2332 7818 2360 8978
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2424 8566 2452 8842
rect 2412 8560 2464 8566
rect 2412 8502 2464 8508
rect 2424 7886 2452 8502
rect 2516 8498 2544 9046
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2596 8900 2648 8906
rect 2596 8842 2648 8848
rect 2608 8634 2636 8842
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2424 7342 2452 7822
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2332 7002 2360 7210
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2332 6866 2360 6938
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2700 6458 2728 7346
rect 2792 7313 2820 8978
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2778 7304 2834 7313
rect 2778 7239 2834 7248
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 2056 4622 2084 5102
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 1676 4480 1728 4486
rect 1676 4422 1728 4428
rect 1688 4321 1716 4422
rect 1674 4312 1730 4321
rect 2056 4282 2084 4558
rect 1674 4247 1730 4256
rect 2044 4276 2096 4282
rect 2044 4218 2096 4224
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1216 3528 1268 3534
rect 1216 3470 1268 3476
rect 1858 3496 1914 3505
rect 388 1012 440 1018
rect 388 954 440 960
rect 400 480 428 954
rect 1228 480 1256 3470
rect 1858 3431 1914 3440
rect 1872 2650 1900 3431
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 1964 2514 1992 3878
rect 2332 2990 2360 6054
rect 2792 5828 2820 7239
rect 2884 5953 2912 8774
rect 2976 8294 3004 9132
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2962 8120 3018 8129
rect 2962 8055 3018 8064
rect 2976 8022 3004 8055
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2976 6866 3004 7142
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2976 6322 3004 6802
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2870 5944 2926 5953
rect 2870 5879 2926 5888
rect 2792 5800 2912 5828
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2412 4752 2464 4758
rect 2412 4694 2464 4700
rect 2424 4214 2452 4694
rect 2412 4208 2464 4214
rect 2412 4150 2464 4156
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 2136 2916 2188 2922
rect 2136 2858 2188 2864
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 2148 480 2176 2858
rect 2700 2650 2728 5714
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2792 4758 2820 4966
rect 2780 4752 2832 4758
rect 2780 4694 2832 4700
rect 2778 3904 2834 3913
rect 2778 3839 2834 3848
rect 2792 3738 2820 3839
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 386 0 442 480
rect 1214 0 1270 480
rect 2134 0 2190 480
rect 2792 241 2820 2994
rect 2884 2990 2912 5800
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 2976 1873 3004 6122
rect 3068 5137 3096 9318
rect 3160 7410 3188 10066
rect 3252 7993 3280 10406
rect 3344 9761 3372 11018
rect 3436 10985 3464 11494
rect 3528 11150 3556 11562
rect 3606 11384 3662 11393
rect 3606 11319 3662 11328
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3422 10976 3478 10985
rect 3422 10911 3478 10920
rect 3436 10538 3464 10911
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3422 10160 3478 10169
rect 3422 10095 3424 10104
rect 3476 10095 3478 10104
rect 3424 10066 3476 10072
rect 3528 10062 3556 10610
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3330 9752 3386 9761
rect 3330 9687 3386 9696
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3528 8974 3556 9318
rect 3424 8968 3476 8974
rect 3422 8936 3424 8945
rect 3516 8968 3568 8974
rect 3476 8936 3478 8945
rect 3516 8910 3568 8916
rect 3422 8871 3478 8880
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 3238 7984 3294 7993
rect 3238 7919 3294 7928
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3252 5778 3280 7754
rect 3344 6361 3372 8502
rect 3330 6352 3386 6361
rect 3330 6287 3386 6296
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3436 5658 3464 8871
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3528 8498 3556 8774
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3344 5630 3464 5658
rect 3528 8004 3556 8230
rect 3620 8129 3648 11319
rect 3712 10282 3740 14991
rect 3804 13394 3832 15399
rect 4080 15230 4108 16623
rect 5538 16520 5594 17000
rect 7746 16520 7802 17000
rect 9954 16520 10010 17000
rect 12162 16520 12218 17000
rect 14370 16520 14426 17000
rect 16578 16520 16634 17000
rect 17958 16688 18014 16697
rect 17958 16623 18014 16632
rect 4068 15224 4120 15230
rect 4068 15166 4120 15172
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 4528 14476 4580 14482
rect 4528 14418 4580 14424
rect 3921 14172 4217 14192
rect 3977 14170 4001 14172
rect 4057 14170 4081 14172
rect 4137 14170 4161 14172
rect 3999 14118 4001 14170
rect 4063 14118 4075 14170
rect 4137 14118 4139 14170
rect 3977 14116 4001 14118
rect 4057 14116 4081 14118
rect 4137 14116 4161 14118
rect 3921 14096 4217 14116
rect 4540 14074 4568 14418
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4356 13530 4384 13670
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 4080 13297 4108 13466
rect 4066 13288 4122 13297
rect 4066 13223 4122 13232
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 3921 13084 4217 13104
rect 3977 13082 4001 13084
rect 4057 13082 4081 13084
rect 4137 13082 4161 13084
rect 3999 13030 4001 13082
rect 4063 13030 4075 13082
rect 4137 13030 4139 13082
rect 3977 13028 4001 13030
rect 4057 13028 4081 13030
rect 4137 13028 4161 13030
rect 3921 13008 4217 13028
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4066 12880 4122 12889
rect 4122 12838 4200 12866
rect 4066 12815 4122 12824
rect 3976 12640 4028 12646
rect 3974 12608 3976 12617
rect 4028 12608 4030 12617
rect 3974 12543 4030 12552
rect 4172 12238 4200 12838
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3804 11898 3832 12038
rect 3921 11996 4217 12016
rect 3977 11994 4001 11996
rect 4057 11994 4081 11996
rect 4137 11994 4161 11996
rect 3999 11942 4001 11994
rect 4063 11942 4075 11994
rect 4137 11942 4139 11994
rect 3977 11940 4001 11942
rect 4057 11940 4081 11942
rect 4137 11940 4161 11942
rect 3921 11920 4217 11940
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 4264 11694 4292 12922
rect 4356 12374 4384 13126
rect 4724 12986 4752 14350
rect 5368 13938 5396 14486
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 4816 12986 4844 13874
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4436 12776 4488 12782
rect 4816 12730 4844 12922
rect 4436 12718 4488 12724
rect 4344 12368 4396 12374
rect 4344 12310 4396 12316
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 3792 11620 3844 11626
rect 3792 11562 3844 11568
rect 3976 11620 4028 11626
rect 3976 11562 4028 11568
rect 3804 11218 3832 11562
rect 3792 11212 3844 11218
rect 3792 11154 3844 11160
rect 3804 10674 3832 11154
rect 3988 11082 4016 11562
rect 4448 11558 4476 12718
rect 4724 12714 4844 12730
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 4712 12708 4844 12714
rect 4764 12702 4844 12708
rect 4712 12650 4764 12656
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 4526 11792 4582 11801
rect 4526 11727 4582 11736
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4448 11234 4476 11494
rect 4264 11206 4476 11234
rect 4264 11150 4292 11206
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 3921 10908 4217 10928
rect 3977 10906 4001 10908
rect 4057 10906 4081 10908
rect 4137 10906 4161 10908
rect 3999 10854 4001 10906
rect 4063 10854 4075 10906
rect 4137 10854 4139 10906
rect 3977 10852 4001 10854
rect 4057 10852 4081 10854
rect 4137 10852 4161 10854
rect 3921 10832 4217 10852
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3974 10568 4030 10577
rect 3974 10503 4030 10512
rect 3712 10254 3832 10282
rect 3698 10160 3754 10169
rect 3698 10095 3754 10104
rect 3712 8480 3740 10095
rect 3804 9081 3832 10254
rect 3988 10198 4016 10503
rect 4068 10464 4120 10470
rect 4172 10452 4200 10678
rect 4120 10424 4200 10452
rect 4068 10406 4120 10412
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 4172 9994 4200 10424
rect 4448 10266 4476 11206
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 4160 9988 4212 9994
rect 4160 9930 4212 9936
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 3921 9820 4217 9840
rect 3977 9818 4001 9820
rect 4057 9818 4081 9820
rect 4137 9818 4161 9820
rect 3999 9766 4001 9818
rect 4063 9766 4075 9818
rect 4137 9766 4139 9818
rect 3977 9764 4001 9766
rect 4057 9764 4081 9766
rect 4137 9764 4161 9766
rect 3921 9744 4217 9764
rect 4066 9344 4122 9353
rect 4066 9279 4122 9288
rect 4080 9110 4108 9279
rect 4068 9104 4120 9110
rect 3790 9072 3846 9081
rect 4068 9046 4120 9052
rect 3790 9007 3846 9016
rect 3921 8732 4217 8752
rect 3977 8730 4001 8732
rect 4057 8730 4081 8732
rect 4137 8730 4161 8732
rect 3999 8678 4001 8730
rect 4063 8678 4075 8730
rect 4137 8678 4139 8730
rect 3977 8676 4001 8678
rect 4057 8676 4081 8678
rect 4137 8676 4161 8678
rect 3921 8656 4217 8676
rect 3712 8452 3832 8480
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3606 8120 3662 8129
rect 3606 8055 3662 8064
rect 3608 8016 3660 8022
rect 3528 7976 3608 8004
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3054 5128 3110 5137
rect 3160 5098 3188 5510
rect 3054 5063 3110 5072
rect 3148 5092 3200 5098
rect 3148 5034 3200 5040
rect 3160 4758 3188 5034
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 3160 3194 3188 3470
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3252 3097 3280 4966
rect 3344 4622 3372 5630
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 3238 3088 3294 3097
rect 3238 3023 3294 3032
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 2962 1864 3018 1873
rect 2962 1799 3018 1808
rect 3068 480 3096 2382
rect 3344 2378 3372 3538
rect 3332 2372 3384 2378
rect 3332 2314 3384 2320
rect 3436 1465 3464 5510
rect 3528 2650 3556 7976
rect 3608 7958 3660 7964
rect 3606 7712 3662 7721
rect 3606 7647 3662 7656
rect 3620 6186 3648 7647
rect 3712 7342 3740 8298
rect 3804 7993 3832 8452
rect 4066 8392 4122 8401
rect 4264 8378 4292 9862
rect 4344 9444 4396 9450
rect 4344 9386 4396 9392
rect 4122 8350 4292 8378
rect 4066 8327 4122 8336
rect 4356 8276 4384 9386
rect 4448 8838 4476 10202
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4448 8430 4476 8774
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 4264 8248 4384 8276
rect 3790 7984 3846 7993
rect 3790 7919 3846 7928
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3804 7177 3832 7686
rect 3921 7644 4217 7664
rect 3977 7642 4001 7644
rect 4057 7642 4081 7644
rect 4137 7642 4161 7644
rect 3999 7590 4001 7642
rect 4063 7590 4075 7642
rect 4137 7590 4139 7642
rect 3977 7588 4001 7590
rect 4057 7588 4081 7590
rect 4137 7588 4161 7590
rect 3921 7568 4217 7588
rect 3790 7168 3846 7177
rect 3790 7103 3846 7112
rect 3976 6928 4028 6934
rect 4264 6916 4292 8248
rect 4540 7970 4568 11727
rect 4632 8090 4660 12106
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4724 10470 4752 11630
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4724 9110 4752 10406
rect 4908 10146 4936 12242
rect 5092 12238 5120 12718
rect 5172 12368 5224 12374
rect 5172 12310 5224 12316
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 5000 11218 5028 11494
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5184 10810 5212 12310
rect 5276 11762 5304 13670
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 5368 12646 5396 13330
rect 5460 13326 5488 13874
rect 5552 13802 5580 16520
rect 6886 14716 7182 14736
rect 6942 14714 6966 14716
rect 7022 14714 7046 14716
rect 7102 14714 7126 14716
rect 6964 14662 6966 14714
rect 7028 14662 7040 14714
rect 7102 14662 7104 14714
rect 6942 14660 6966 14662
rect 7022 14660 7046 14662
rect 7102 14660 7126 14662
rect 6886 14640 7182 14660
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6380 13530 6408 13670
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5460 12782 5488 13262
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 4908 10118 5028 10146
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 4802 9752 4858 9761
rect 4802 9687 4858 9696
rect 4816 9382 4844 9687
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4724 8498 4752 8774
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4028 6888 4292 6916
rect 4356 7942 4568 7970
rect 3976 6870 4028 6876
rect 3790 6760 3846 6769
rect 4356 6746 4384 7942
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 3790 6695 3846 6704
rect 4264 6718 4476 6746
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 3700 6112 3752 6118
rect 3698 6080 3700 6089
rect 3752 6080 3754 6089
rect 3698 6015 3754 6024
rect 3804 5574 3832 6695
rect 3921 6556 4217 6576
rect 3977 6554 4001 6556
rect 4057 6554 4081 6556
rect 4137 6554 4161 6556
rect 3999 6502 4001 6554
rect 4063 6502 4075 6554
rect 4137 6502 4139 6554
rect 3977 6500 4001 6502
rect 4057 6500 4081 6502
rect 4137 6500 4161 6502
rect 3921 6480 4217 6500
rect 4264 6440 4292 6718
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4172 6412 4292 6440
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4080 5710 4108 6326
rect 4172 5778 4200 6412
rect 4356 6322 4384 6598
rect 4448 6497 4476 6718
rect 4434 6488 4490 6497
rect 4540 6458 4568 7822
rect 4632 6934 4660 8026
rect 4724 7886 4752 8434
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4724 7410 4752 7822
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4620 6928 4672 6934
rect 4620 6870 4672 6876
rect 4434 6423 4490 6432
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4356 5846 4384 6258
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4356 5642 4384 5782
rect 4344 5636 4396 5642
rect 4344 5578 4396 5584
rect 3792 5568 3844 5574
rect 3698 5536 3754 5545
rect 3792 5510 3844 5516
rect 3698 5471 3754 5480
rect 3712 5370 3740 5471
rect 3921 5468 4217 5488
rect 3977 5466 4001 5468
rect 4057 5466 4081 5468
rect 4137 5466 4161 5468
rect 3999 5414 4001 5466
rect 4063 5414 4075 5466
rect 4137 5414 4139 5466
rect 3977 5412 4001 5414
rect 4057 5412 4081 5414
rect 4137 5412 4161 5414
rect 3921 5392 4217 5412
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 4356 5234 4384 5578
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4448 5114 4476 6326
rect 4264 5086 4476 5114
rect 4540 5098 4568 6394
rect 4724 5778 4752 7142
rect 4816 7002 4844 7346
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4816 5574 4844 6938
rect 4908 6118 4936 9930
rect 5000 7993 5028 10118
rect 5092 9654 5120 10406
rect 5184 10266 5212 10406
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5368 10146 5396 12582
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 10713 5580 12174
rect 6288 11898 6316 13330
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6564 12986 6592 13262
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6656 12866 6684 13806
rect 6886 13628 7182 13648
rect 6942 13626 6966 13628
rect 7022 13626 7046 13628
rect 7102 13626 7126 13628
rect 6964 13574 6966 13626
rect 7028 13574 7040 13626
rect 7102 13574 7104 13626
rect 6942 13572 6966 13574
rect 7022 13572 7046 13574
rect 7102 13572 7126 13574
rect 6886 13552 7182 13572
rect 7484 13530 7512 13874
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 6564 12838 6684 12866
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6380 11558 6408 12242
rect 6564 12073 6592 12838
rect 6932 12714 6960 13262
rect 7484 12782 7512 13466
rect 7760 13462 7788 16520
rect 9496 15224 9548 15230
rect 9496 15166 9548 15172
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 6748 12374 6776 12650
rect 6886 12540 7182 12560
rect 6942 12538 6966 12540
rect 7022 12538 7046 12540
rect 7102 12538 7126 12540
rect 6964 12486 6966 12538
rect 7028 12486 7040 12538
rect 7102 12486 7104 12538
rect 6942 12484 6966 12486
rect 7022 12484 7046 12486
rect 7102 12484 7126 12486
rect 6886 12464 7182 12484
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6550 12064 6606 12073
rect 6550 11999 6606 12008
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6104 11257 6132 11494
rect 6090 11248 6146 11257
rect 6090 11183 6146 11192
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5538 10704 5594 10713
rect 5538 10639 5594 10648
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5276 10118 5396 10146
rect 5172 9988 5224 9994
rect 5172 9930 5224 9936
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 5184 9586 5212 9930
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5184 8362 5212 9522
rect 5276 9450 5304 10118
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 4986 7984 5042 7993
rect 4986 7919 5042 7928
rect 5184 7546 5212 8298
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5276 7426 5304 9046
rect 5368 8090 5396 9998
rect 5460 9518 5488 10406
rect 5552 10198 5580 10639
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5184 7398 5304 7426
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4528 5092 4580 5098
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4080 4690 4108 4762
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3620 2990 3648 4558
rect 3700 4480 3752 4486
rect 3700 4422 3752 4428
rect 3712 4010 3740 4422
rect 3804 4282 3832 4626
rect 3921 4380 4217 4400
rect 3977 4378 4001 4380
rect 4057 4378 4081 4380
rect 4137 4378 4161 4380
rect 3999 4326 4001 4378
rect 4063 4326 4075 4378
rect 4137 4326 4139 4378
rect 3977 4324 4001 4326
rect 4057 4324 4081 4326
rect 4137 4324 4161 4326
rect 3921 4304 4217 4324
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 3700 4004 3752 4010
rect 3700 3946 3752 3952
rect 3792 4004 3844 4010
rect 3792 3946 3844 3952
rect 3712 3058 3740 3946
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3712 2446 3740 2994
rect 3700 2440 3752 2446
rect 3700 2382 3752 2388
rect 3698 2272 3754 2281
rect 3698 2207 3754 2216
rect 3712 2106 3740 2207
rect 3700 2100 3752 2106
rect 3700 2042 3752 2048
rect 3422 1456 3478 1465
rect 3422 1391 3478 1400
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 3344 649 3372 1294
rect 3804 1057 3832 3946
rect 4264 3942 4292 5086
rect 4528 5034 4580 5040
rect 4344 5024 4396 5030
rect 4342 4992 4344 5001
rect 4436 5024 4488 5030
rect 4396 4992 4398 5001
rect 4436 4966 4488 4972
rect 4342 4927 4398 4936
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4356 4282 4384 4626
rect 4448 4282 4476 4966
rect 4816 4826 4844 5510
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4356 3534 4384 4218
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4448 3346 4476 4218
rect 4816 3466 4844 4762
rect 4908 4078 4936 6054
rect 5000 5710 5028 6190
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 5092 5556 5120 6666
rect 5184 6202 5212 7398
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5276 6322 5304 6802
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5448 6248 5500 6254
rect 5262 6216 5318 6225
rect 5184 6174 5262 6202
rect 5448 6190 5500 6196
rect 5262 6151 5318 6160
rect 5276 6118 5304 6151
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5172 5840 5224 5846
rect 5170 5808 5172 5817
rect 5224 5808 5226 5817
rect 5460 5778 5488 6190
rect 5170 5743 5226 5752
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5000 5528 5120 5556
rect 5000 5370 5028 5528
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 4896 4072 4948 4078
rect 4948 4032 5028 4060
rect 4896 4014 4948 4020
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4264 3318 4476 3346
rect 3921 3292 4217 3312
rect 3977 3290 4001 3292
rect 4057 3290 4081 3292
rect 4137 3290 4161 3292
rect 3999 3238 4001 3290
rect 4063 3238 4075 3290
rect 4137 3238 4139 3290
rect 3977 3236 4001 3238
rect 4057 3236 4081 3238
rect 4137 3236 4161 3238
rect 3921 3216 4217 3236
rect 4066 2680 4122 2689
rect 4066 2615 4122 2624
rect 4080 2514 4108 2615
rect 4264 2582 4292 3318
rect 4908 2990 4936 3878
rect 5000 3738 5028 4032
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 5000 3058 5028 3334
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 4252 2576 4304 2582
rect 4252 2518 4304 2524
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4896 2372 4948 2378
rect 4896 2314 4948 2320
rect 3921 2204 4217 2224
rect 3977 2202 4001 2204
rect 4057 2202 4081 2204
rect 4137 2202 4161 2204
rect 3999 2150 4001 2202
rect 4063 2150 4075 2202
rect 4137 2150 4139 2202
rect 3977 2148 4001 2150
rect 4057 2148 4081 2150
rect 4137 2148 4161 2150
rect 3921 2128 4217 2148
rect 3976 1420 4028 1426
rect 3976 1362 4028 1368
rect 3790 1048 3846 1057
rect 3790 983 3846 992
rect 3330 640 3386 649
rect 3330 575 3386 584
rect 3988 480 4016 1362
rect 4908 480 4936 2314
rect 5092 2106 5120 5306
rect 5368 5166 5396 5646
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5184 4146 5212 4966
rect 5552 4842 5580 10134
rect 5736 9654 5764 11086
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5828 10130 5856 11018
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5644 8838 5672 9318
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5736 7886 5764 9454
rect 5920 9110 5948 10610
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 5920 8634 5948 9046
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5736 7274 5764 7822
rect 5724 7268 5776 7274
rect 5724 7210 5776 7216
rect 5908 6180 5960 6186
rect 5908 6122 5960 6128
rect 5920 6089 5948 6122
rect 5906 6080 5962 6089
rect 5906 6015 5962 6024
rect 5368 4814 5580 4842
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 5184 3670 5212 3946
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5184 3058 5212 3334
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5172 2644 5224 2650
rect 5368 2632 5396 4814
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5460 4146 5488 4422
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5460 3670 5488 4082
rect 5632 4072 5684 4078
rect 5736 4060 5764 4422
rect 6012 4078 6040 10678
rect 6104 7954 6132 11183
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6288 9586 6316 10610
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6196 7206 6224 7414
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6104 5914 6132 6054
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6196 4690 6224 7142
rect 6380 6440 6408 11494
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6288 6412 6408 6440
rect 6288 5166 6316 6412
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6380 5370 6408 6258
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6276 5160 6328 5166
rect 6276 5102 6328 5108
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6092 4548 6144 4554
rect 6092 4490 6144 4496
rect 5684 4032 5764 4060
rect 6000 4072 6052 4078
rect 5632 4014 5684 4020
rect 6000 4014 6052 4020
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5552 3194 5580 3538
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5224 2604 5396 2632
rect 5172 2586 5224 2592
rect 5460 2514 5488 3062
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5080 2100 5132 2106
rect 5080 2042 5132 2048
rect 5644 1426 5672 2382
rect 5632 1420 5684 1426
rect 5632 1362 5684 1368
rect 5828 480 5856 3946
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 5920 2854 5948 3062
rect 6104 3058 6132 4490
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6012 2310 6040 2790
rect 6092 2576 6144 2582
rect 6288 2564 6316 5102
rect 6380 4758 6408 5306
rect 6368 4752 6420 4758
rect 6368 4694 6420 4700
rect 6472 4078 6500 11018
rect 6564 10033 6592 11999
rect 6932 11762 6960 12106
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 7024 11694 7052 12174
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 6886 11452 7182 11472
rect 6942 11450 6966 11452
rect 7022 11450 7046 11452
rect 7102 11450 7126 11452
rect 6964 11398 6966 11450
rect 7028 11398 7040 11450
rect 7102 11398 7104 11450
rect 6942 11396 6966 11398
rect 7022 11396 7046 11398
rect 7102 11396 7126 11398
rect 6886 11376 7182 11396
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6550 10024 6606 10033
rect 6550 9959 6606 9968
rect 6656 8566 6684 11154
rect 7024 10810 7052 11222
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6564 7002 6592 7822
rect 6656 7342 6684 8502
rect 6748 8294 6776 10406
rect 6886 10364 7182 10384
rect 6942 10362 6966 10364
rect 7022 10362 7046 10364
rect 7102 10362 7126 10364
rect 6964 10310 6966 10362
rect 7028 10310 7040 10362
rect 7102 10310 7104 10362
rect 6942 10308 6966 10310
rect 7022 10308 7046 10310
rect 7102 10308 7126 10310
rect 6886 10288 7182 10308
rect 6918 10160 6974 10169
rect 6918 10095 6974 10104
rect 6932 9364 6960 10095
rect 7010 10024 7066 10033
rect 7010 9959 7066 9968
rect 7024 9489 7052 9959
rect 7300 9586 7328 12038
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7010 9480 7066 9489
rect 7010 9415 7066 9424
rect 7288 9376 7340 9382
rect 6932 9336 7288 9364
rect 7288 9318 7340 9324
rect 6886 9276 7182 9296
rect 6942 9274 6966 9276
rect 7022 9274 7046 9276
rect 7102 9274 7126 9276
rect 6964 9222 6966 9274
rect 7028 9222 7040 9274
rect 7102 9222 7104 9274
rect 6942 9220 6966 9222
rect 7022 9220 7046 9222
rect 7102 9220 7126 9222
rect 6886 9200 7182 9220
rect 7300 9081 7328 9318
rect 7286 9072 7342 9081
rect 7286 9007 7342 9016
rect 7392 9058 7420 12174
rect 7484 12170 7512 12718
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7484 10452 7512 11766
rect 7576 10606 7604 12174
rect 7668 11694 7696 12718
rect 7944 12646 7972 12786
rect 8128 12646 8156 13806
rect 9508 13705 9536 15166
rect 9968 14634 9996 16520
rect 9968 14606 10364 14634
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10060 14362 10088 14418
rect 10060 14334 10272 14362
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9692 13870 9720 14214
rect 9852 14172 10148 14192
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 9930 14118 9932 14170
rect 9994 14118 10006 14170
rect 10068 14118 10070 14170
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 9852 14096 10148 14116
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 10138 13832 10194 13841
rect 9494 13696 9550 13705
rect 9494 13631 9550 13640
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 8128 12481 8156 12582
rect 7746 12472 7802 12481
rect 7746 12407 7802 12416
rect 8114 12472 8170 12481
rect 8312 12442 8340 13330
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 8574 12744 8630 12753
rect 8574 12679 8630 12688
rect 8114 12407 8170 12416
rect 8300 12436 8352 12442
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7668 11014 7696 11630
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7668 10674 7696 10950
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 7484 10424 7604 10452
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7484 9586 7512 10066
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7576 9518 7604 10424
rect 7668 10198 7696 10610
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7668 9194 7696 10134
rect 7484 9178 7696 9194
rect 7472 9172 7696 9178
rect 7524 9166 7696 9172
rect 7472 9114 7524 9120
rect 7564 9104 7616 9110
rect 7392 9052 7564 9058
rect 7392 9046 7616 9052
rect 7392 9030 7604 9046
rect 7300 8786 7328 9007
rect 7392 8906 7420 9030
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 7300 8758 7512 8786
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6886 8188 7182 8208
rect 6942 8186 6966 8188
rect 7022 8186 7046 8188
rect 7102 8186 7126 8188
rect 6964 8134 6966 8186
rect 7028 8134 7040 8186
rect 7102 8134 7104 8186
rect 6942 8132 6966 8134
rect 7022 8132 7046 8134
rect 7102 8132 7126 8134
rect 6886 8112 7182 8132
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6564 5681 6592 6734
rect 6748 6186 6776 7822
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 7116 7546 7144 7754
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7196 7336 7248 7342
rect 7194 7304 7196 7313
rect 7248 7304 7250 7313
rect 7194 7239 7250 7248
rect 6886 7100 7182 7120
rect 6942 7098 6966 7100
rect 7022 7098 7046 7100
rect 7102 7098 7126 7100
rect 6964 7046 6966 7098
rect 7028 7046 7040 7098
rect 7102 7046 7104 7098
rect 6942 7044 6966 7046
rect 7022 7044 7046 7046
rect 7102 7044 7126 7046
rect 6886 7024 7182 7044
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7116 6458 7144 6802
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6748 5914 6776 6122
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 6886 6012 7182 6032
rect 6942 6010 6966 6012
rect 7022 6010 7046 6012
rect 7102 6010 7126 6012
rect 6964 5958 6966 6010
rect 7028 5958 7040 6010
rect 7102 5958 7104 6010
rect 6942 5956 6966 5958
rect 7022 5956 7046 5958
rect 7102 5956 7126 5958
rect 6886 5936 7182 5956
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 6550 5672 6606 5681
rect 6550 5607 6606 5616
rect 6564 4842 6592 5607
rect 7116 5234 7144 5714
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 6734 4992 6790 5001
rect 6734 4927 6790 4936
rect 6564 4814 6684 4842
rect 6656 4690 6684 4814
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6748 4570 6776 4927
rect 6886 4924 7182 4944
rect 6942 4922 6966 4924
rect 7022 4922 7046 4924
rect 7102 4922 7126 4924
rect 6964 4870 6966 4922
rect 7028 4870 7040 4922
rect 7102 4870 7104 4922
rect 6942 4868 6966 4870
rect 7022 4868 7046 4870
rect 7102 4868 7126 4870
rect 6886 4848 7182 4868
rect 7300 4826 7328 6054
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 6748 4542 6868 4570
rect 6840 4486 6868 4542
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6144 2536 6316 2564
rect 6092 2518 6144 2524
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 6564 626 6592 3946
rect 6748 3942 6776 4422
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6886 3836 7182 3856
rect 6942 3834 6966 3836
rect 7022 3834 7046 3836
rect 7102 3834 7126 3836
rect 6964 3782 6966 3834
rect 7028 3782 7040 3834
rect 7102 3782 7104 3834
rect 6942 3780 6966 3782
rect 7022 3780 7046 3782
rect 7102 3780 7126 3782
rect 6886 3760 7182 3780
rect 6886 2748 7182 2768
rect 6942 2746 6966 2748
rect 7022 2746 7046 2748
rect 7102 2746 7126 2748
rect 6964 2694 6966 2746
rect 7028 2694 7040 2746
rect 7102 2694 7104 2746
rect 6942 2692 6966 2694
rect 7022 2692 7046 2694
rect 7102 2692 7126 2694
rect 6886 2672 7182 2692
rect 7392 2514 7420 7958
rect 7484 7018 7512 8758
rect 7668 8430 7696 9166
rect 7760 8945 7788 12407
rect 8300 12378 8352 12384
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8116 12232 8168 12238
rect 8114 12200 8116 12209
rect 8168 12200 8170 12209
rect 8114 12135 8170 12144
rect 8208 12096 8260 12102
rect 8300 12096 8352 12102
rect 8208 12038 8260 12044
rect 8298 12064 8300 12073
rect 8352 12064 8354 12073
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 8036 10690 8064 10746
rect 7944 10662 8064 10690
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 7746 8936 7802 8945
rect 7746 8871 7802 8880
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7576 7206 7604 8230
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7484 6990 7604 7018
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7484 6254 7512 6802
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7484 5574 7512 6190
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 7484 4690 7512 5238
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7484 2582 7512 4150
rect 7576 4146 7604 6990
rect 7668 6866 7696 7346
rect 7760 7342 7788 8871
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7760 5658 7788 7142
rect 7668 5630 7788 5658
rect 7668 5234 7696 5630
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7668 4078 7696 4626
rect 7760 4622 7788 5510
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7760 3398 7788 4558
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 7852 2514 7880 10542
rect 7944 9450 7972 10662
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 8036 9994 8064 10474
rect 8220 10266 8248 12038
rect 8298 11999 8354 12008
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 8036 9654 8064 9930
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8036 9110 8064 9318
rect 8024 9104 8076 9110
rect 7944 9064 8024 9092
rect 7944 5817 7972 9064
rect 8024 9046 8076 9052
rect 8128 8480 8156 10202
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8220 9586 8248 9998
rect 8300 9920 8352 9926
rect 8352 9897 8432 9908
rect 8352 9888 8446 9897
rect 8352 9880 8390 9888
rect 8300 9862 8352 9868
rect 8390 9823 8446 9832
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8312 9625 8340 9658
rect 8298 9616 8354 9625
rect 8208 9580 8260 9586
rect 8298 9551 8354 9560
rect 8208 9522 8260 9528
rect 8220 9178 8248 9522
rect 8404 9518 8432 9658
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8128 8452 8248 8480
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 8036 7002 8064 7686
rect 8024 6996 8076 7002
rect 8024 6938 8076 6944
rect 8036 5914 8064 6938
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 7930 5808 7986 5817
rect 7930 5743 7986 5752
rect 7944 4078 7972 5743
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8128 2854 8156 8298
rect 8220 7970 8248 8452
rect 8220 7942 8340 7970
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8220 7750 8248 7822
rect 8312 7750 8340 7942
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8220 6458 8248 6802
rect 8298 6488 8354 6497
rect 8208 6452 8260 6458
rect 8298 6423 8300 6432
rect 8208 6394 8260 6400
rect 8352 6423 8354 6432
rect 8300 6394 8352 6400
rect 8404 6338 8432 9318
rect 8496 9042 8524 12310
rect 8588 11830 8616 12679
rect 9048 12442 9076 13262
rect 9140 12986 9168 13262
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 8852 12300 8904 12306
rect 8852 12242 8904 12248
rect 8576 11824 8628 11830
rect 8576 11766 8628 11772
rect 8864 11762 8892 12242
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 9048 11898 9076 12174
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8956 11218 8984 11834
rect 9140 11694 9168 12922
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9232 12238 9260 12650
rect 9310 12336 9366 12345
rect 9310 12271 9366 12280
rect 9404 12300 9456 12306
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9324 12170 9352 12271
rect 9404 12242 9456 12248
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9324 11506 9352 12106
rect 9048 11478 9352 11506
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8956 10742 8984 11154
rect 8944 10736 8996 10742
rect 8944 10678 8996 10684
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8588 8090 8616 10406
rect 8956 10198 8984 10229
rect 8944 10192 8996 10198
rect 8942 10160 8944 10169
rect 8996 10160 8998 10169
rect 8942 10095 8998 10104
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8680 9518 8708 9998
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 8772 9625 8800 9930
rect 8758 9616 8814 9625
rect 8758 9551 8814 9560
rect 8956 9518 8984 10095
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8772 7342 8800 8230
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8864 7857 8892 8026
rect 8944 7880 8996 7886
rect 8850 7848 8906 7857
rect 8944 7822 8996 7828
rect 8850 7783 8906 7792
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8220 6310 8432 6338
rect 8220 5030 8248 6310
rect 8496 6254 8524 7278
rect 8956 7274 8984 7822
rect 8944 7268 8996 7274
rect 8944 7210 8996 7216
rect 8956 7002 8984 7210
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8484 6248 8536 6254
rect 8390 6216 8446 6225
rect 8484 6190 8536 6196
rect 8390 6151 8446 6160
rect 8404 6066 8432 6151
rect 8404 6038 8524 6066
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8220 4214 8248 4966
rect 8312 4826 8340 5170
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8496 3754 8524 6038
rect 8588 3942 8616 6598
rect 8864 5370 8892 6870
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8680 4690 8708 5170
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8680 4146 8708 4626
rect 8864 4554 8892 4762
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 9048 4185 9076 11478
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 9140 10810 9168 11222
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9140 9518 9168 10202
rect 9324 9654 9352 11290
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9416 8838 9444 12242
rect 9508 10810 9536 13631
rect 9600 13410 9628 13806
rect 10138 13767 10140 13776
rect 10192 13767 10194 13776
rect 10140 13738 10192 13744
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9600 13382 9904 13410
rect 9876 13258 9904 13382
rect 9968 13258 9996 13466
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9600 11354 9628 11494
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9508 10062 9536 10746
rect 9600 10266 9628 11154
rect 9692 10674 9720 13126
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9784 10606 9812 13194
rect 9852 13084 10148 13104
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 9930 13030 9932 13082
rect 9994 13030 10006 13082
rect 10068 13030 10070 13082
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 9852 13008 10148 13028
rect 9852 11996 10148 12016
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 9930 11942 9932 11994
rect 9994 11942 10006 11994
rect 10068 11942 10070 11994
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 9852 11920 10148 11940
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10060 11257 10088 11494
rect 10046 11248 10102 11257
rect 10046 11183 10102 11192
rect 9852 10908 10148 10928
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 9930 10854 9932 10906
rect 9994 10854 10006 10906
rect 10068 10854 10070 10906
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 9852 10832 10148 10852
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9862 10568 9918 10577
rect 9862 10503 9918 10512
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9876 9908 9904 10503
rect 9494 9888 9550 9897
rect 9494 9823 9550 9832
rect 9784 9880 9904 9908
rect 9508 9586 9536 9823
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 9232 5302 9260 8502
rect 9508 8362 9536 9318
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9600 8566 9628 8978
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9416 6186 9444 7142
rect 9508 6225 9536 8298
rect 9784 8072 9812 9880
rect 9852 9820 10148 9840
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 9930 9766 9932 9818
rect 9994 9766 10006 9818
rect 10068 9766 10070 9818
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 9852 9744 10148 9764
rect 10244 9654 10272 14334
rect 10336 13802 10364 14606
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 10416 14476 10468 14482
rect 10416 14418 10468 14424
rect 10324 13796 10376 13802
rect 10324 13738 10376 13744
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 10336 12170 10364 12650
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10336 11762 10364 12106
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10336 11354 10364 11698
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10336 10198 10364 10950
rect 10324 10192 10376 10198
rect 10324 10134 10376 10140
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10230 9480 10286 9489
rect 9864 9444 9916 9450
rect 10230 9415 10286 9424
rect 9864 9386 9916 9392
rect 9876 8906 9904 9386
rect 10046 9072 10102 9081
rect 10046 9007 10048 9016
rect 10100 9007 10102 9016
rect 10048 8978 10100 8984
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9852 8732 10148 8752
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 9930 8678 9932 8730
rect 9994 8678 10006 8730
rect 10068 8678 10070 8730
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 9852 8656 10148 8676
rect 9784 8044 9904 8072
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 9692 7274 9720 7958
rect 9876 7954 9904 8044
rect 10048 8016 10100 8022
rect 10046 7984 10048 7993
rect 10100 7984 10102 7993
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9864 7948 9916 7954
rect 10046 7919 10102 7928
rect 10140 7948 10192 7954
rect 9864 7890 9916 7896
rect 10140 7890 10192 7896
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9494 6216 9550 6225
rect 9404 6180 9456 6186
rect 9494 6151 9550 6160
rect 9404 6122 9456 6128
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 9232 5030 9260 5238
rect 9324 5234 9352 5714
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9324 4826 9352 5170
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9324 4214 9352 4762
rect 9312 4208 9364 4214
rect 9034 4176 9090 4185
rect 8668 4140 8720 4146
rect 9312 4150 9364 4156
rect 9034 4111 9090 4120
rect 8668 4082 8720 4088
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8392 3732 8444 3738
rect 8496 3726 8616 3754
rect 8392 3674 8444 3680
rect 8404 2854 8432 3674
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 6564 598 6776 626
rect 6748 480 6776 598
rect 7576 480 7604 2382
rect 8496 480 8524 3470
rect 8588 2854 8616 3726
rect 8680 3398 8708 4082
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8680 3058 8708 3334
rect 8772 3194 8800 3878
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 9048 3126 9076 4111
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9140 3194 9168 3538
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9416 3126 9444 6122
rect 9600 5370 9628 6938
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9692 5166 9720 6734
rect 9784 5370 9812 7890
rect 10152 7857 10180 7890
rect 10138 7848 10194 7857
rect 10138 7783 10194 7792
rect 9852 7644 10148 7664
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 9930 7590 9932 7642
rect 9994 7590 10006 7642
rect 10068 7590 10070 7642
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 9852 7568 10148 7588
rect 10244 7426 10272 9415
rect 10336 8974 10364 10134
rect 10428 9450 10456 14418
rect 10508 14408 10560 14414
rect 11060 14408 11112 14414
rect 10508 14350 10560 14356
rect 10520 13938 10548 14350
rect 10704 14334 11008 14362
rect 11060 14350 11112 14356
rect 10704 14074 10732 14334
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10600 14000 10652 14006
rect 10600 13942 10652 13948
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10324 8968 10376 8974
rect 10322 8936 10324 8945
rect 10416 8968 10468 8974
rect 10376 8936 10378 8945
rect 10416 8910 10468 8916
rect 10322 8871 10378 8880
rect 10428 8650 10456 8910
rect 10520 8906 10548 13670
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10336 8622 10456 8650
rect 10336 8566 10364 8622
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10152 7398 10272 7426
rect 10336 7410 10364 7890
rect 10324 7404 10376 7410
rect 10152 7002 10180 7398
rect 10324 7346 10376 7352
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 9852 6556 10148 6576
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 9930 6502 9932 6554
rect 9994 6502 10006 6554
rect 10068 6502 10070 6554
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 9852 6480 10148 6500
rect 9852 5468 10148 5488
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 9930 5414 9932 5466
rect 9994 5414 10006 5466
rect 10068 5414 10070 5466
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 9852 5392 10148 5412
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 10138 5128 10194 5137
rect 10138 5063 10194 5072
rect 10152 5030 10180 5063
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 9692 4486 9720 4966
rect 9862 4720 9918 4729
rect 9862 4655 9864 4664
rect 9916 4655 9918 4664
rect 9864 4626 9916 4632
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9852 4380 10148 4400
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 9930 4326 9932 4378
rect 9994 4326 10006 4378
rect 10068 4326 10070 4378
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 9852 4304 10148 4324
rect 10244 4146 10272 7278
rect 10336 6934 10364 7346
rect 10324 6928 10376 6934
rect 10324 6870 10376 6876
rect 10336 6458 10364 6870
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10336 5846 10364 6394
rect 10324 5840 10376 5846
rect 10324 5782 10376 5788
rect 10336 4758 10364 5782
rect 10428 5030 10456 7958
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10520 5370 10548 7142
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10324 4752 10376 4758
rect 10428 4729 10456 4966
rect 10324 4694 10376 4700
rect 10414 4720 10470 4729
rect 10336 4146 10364 4694
rect 10414 4655 10470 4664
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 9508 2990 9536 3878
rect 10244 3534 10272 4082
rect 10612 4078 10640 13942
rect 10692 13728 10744 13734
rect 10690 13696 10692 13705
rect 10744 13696 10746 13705
rect 10690 13631 10746 13640
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10704 11830 10732 13330
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10704 11286 10732 11630
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10704 10674 10732 10950
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 10704 9586 10732 10134
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10704 8022 10732 8978
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10704 6934 10732 7822
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10690 5808 10746 5817
rect 10690 5743 10746 5752
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9600 3058 9628 3334
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8772 1018 8800 2790
rect 9784 2650 9812 3402
rect 9852 3292 10148 3312
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 9930 3238 9932 3290
rect 9994 3238 10006 3290
rect 10068 3238 10070 3290
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 9852 3216 10148 3236
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 10336 2446 10364 3674
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10428 3534 10456 3606
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 9852 2204 10148 2224
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 9930 2150 9932 2202
rect 9994 2150 10006 2202
rect 10068 2150 10070 2202
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 9852 2128 10148 2148
rect 9404 2100 9456 2106
rect 9404 2042 9456 2048
rect 8760 1012 8812 1018
rect 8760 954 8812 960
rect 9416 480 9444 2042
rect 10520 1442 10548 3606
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10612 3058 10640 3334
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10704 2990 10732 5743
rect 10796 3602 10824 14214
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10888 9489 10916 12038
rect 10874 9480 10930 9489
rect 10874 9415 10930 9424
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10888 9042 10916 9318
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10888 7342 10916 8570
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10980 7154 11008 14334
rect 11072 13938 11100 14350
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 11072 9926 11100 13874
rect 11164 13530 11192 14554
rect 12176 13938 12204 16520
rect 14278 15464 14334 15473
rect 14278 15399 14334 15408
rect 12817 14716 13113 14736
rect 12873 14714 12897 14716
rect 12953 14714 12977 14716
rect 13033 14714 13057 14716
rect 12895 14662 12897 14714
rect 12959 14662 12971 14714
rect 13033 14662 13035 14714
rect 12873 14660 12897 14662
rect 12953 14660 12977 14662
rect 13033 14660 13057 14662
rect 12817 14640 13113 14660
rect 14292 14550 14320 15399
rect 14280 14544 14332 14550
rect 14280 14486 14332 14492
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12440 13864 12492 13870
rect 11242 13832 11298 13841
rect 11242 13767 11244 13776
rect 11296 13767 11298 13776
rect 11794 13832 11850 13841
rect 12440 13806 12492 13812
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 11794 13767 11850 13776
rect 11244 13738 11296 13744
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11164 12442 11192 13262
rect 11348 12986 11376 13262
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11256 12714 11284 12922
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11348 12442 11376 12922
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11164 11762 11192 12038
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11256 11354 11284 12174
rect 11348 11762 11376 12378
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11440 11014 11468 12718
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 8430 11100 9862
rect 11164 9110 11192 10134
rect 11426 9888 11482 9897
rect 11426 9823 11482 9832
rect 11440 9722 11468 9823
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11348 9178 11376 9318
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 11152 8968 11204 8974
rect 11150 8936 11152 8945
rect 11204 8936 11206 8945
rect 11150 8871 11206 8880
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 11058 7848 11114 7857
rect 11058 7783 11114 7792
rect 10888 7126 11008 7154
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10888 3534 10916 7126
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10980 5914 11008 6190
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 11072 4842 11100 7783
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 11256 5778 11284 6326
rect 11348 6322 11376 7346
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 11532 6186 11560 13466
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11624 12442 11652 12582
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11716 12374 11744 13194
rect 11704 12368 11756 12374
rect 11704 12310 11756 12316
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11624 8906 11652 12174
rect 11808 11898 11836 13767
rect 12452 13462 12480 13806
rect 13280 13734 13308 13806
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 12817 13628 13113 13648
rect 12873 13626 12897 13628
rect 12953 13626 12977 13628
rect 13033 13626 13057 13628
rect 12895 13574 12897 13626
rect 12959 13574 12971 13626
rect 13033 13574 13035 13626
rect 12873 13572 12897 13574
rect 12953 13572 12977 13574
rect 13033 13572 13057 13574
rect 12817 13552 13113 13572
rect 13280 13530 13308 13670
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11900 12782 11928 13262
rect 12624 13184 12676 13190
rect 12676 13132 12756 13138
rect 12624 13126 12756 13132
rect 12636 13110 12756 13126
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 11218 11744 11494
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11704 10532 11756 10538
rect 11704 10474 11756 10480
rect 11716 9722 11744 10474
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11716 9586 11744 9658
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11612 8900 11664 8906
rect 11612 8842 11664 8848
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11624 6730 11652 8298
rect 11716 8022 11744 8434
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11716 7546 11744 7958
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11808 7410 11836 11834
rect 11992 11801 12020 12242
rect 12360 11898 12388 12242
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 11978 11792 12034 11801
rect 11978 11727 12034 11736
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12084 11354 12112 11698
rect 12636 11354 12664 12174
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 11980 11280 12032 11286
rect 11978 11248 11980 11257
rect 12032 11248 12034 11257
rect 11978 11183 12034 11192
rect 11992 10266 12020 11183
rect 12084 10742 12112 11290
rect 12256 11144 12308 11150
rect 12308 11104 12388 11132
rect 12256 11086 12308 11092
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11888 9444 11940 9450
rect 11888 9386 11940 9392
rect 11900 9178 11928 9386
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11992 8786 12020 9862
rect 12084 8974 12112 10678
rect 12256 10532 12308 10538
rect 12256 10474 12308 10480
rect 12268 10266 12296 10474
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 11992 8758 12112 8786
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 12084 6866 12112 8758
rect 12176 7546 12204 10066
rect 12360 9518 12388 11104
rect 12622 10976 12678 10985
rect 12622 10911 12678 10920
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12256 9444 12308 9450
rect 12256 9386 12308 9392
rect 12268 8294 12296 9386
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12346 9072 12402 9081
rect 12346 9007 12402 9016
rect 12360 8974 12388 9007
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12452 8634 12480 9318
rect 12544 9110 12572 10406
rect 12636 10130 12664 10911
rect 12728 10470 12756 13110
rect 13266 12608 13322 12617
rect 12817 12540 13113 12560
rect 13266 12543 13322 12552
rect 12873 12538 12897 12540
rect 12953 12538 12977 12540
rect 13033 12538 13057 12540
rect 12895 12486 12897 12538
rect 12959 12486 12971 12538
rect 13033 12486 13035 12538
rect 12873 12484 12897 12486
rect 12953 12484 12977 12486
rect 13033 12484 13057 12486
rect 12817 12464 13113 12484
rect 13280 12442 13308 12543
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 12817 11452 13113 11472
rect 12873 11450 12897 11452
rect 12953 11450 12977 11452
rect 13033 11450 13057 11452
rect 12895 11398 12897 11450
rect 12959 11398 12971 11450
rect 13033 11398 13035 11450
rect 12873 11396 12897 11398
rect 12953 11396 12977 11398
rect 13033 11396 13057 11398
rect 12817 11376 13113 11396
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 13096 10577 13124 10610
rect 13082 10568 13138 10577
rect 13082 10503 13138 10512
rect 13188 10470 13216 10950
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 12817 10364 13113 10384
rect 12873 10362 12897 10364
rect 12953 10362 12977 10364
rect 13033 10362 13057 10364
rect 12895 10310 12897 10362
rect 12959 10310 12971 10362
rect 13033 10310 13035 10362
rect 12873 10308 12897 10310
rect 12953 10308 12977 10310
rect 13033 10308 13057 10310
rect 12817 10288 13113 10308
rect 13280 10266 13308 11494
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 12624 10124 12676 10130
rect 12676 10084 12756 10112
rect 12624 10066 12676 10072
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12530 8936 12586 8945
rect 12530 8871 12586 8880
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 11612 6724 11664 6730
rect 11612 6666 11664 6672
rect 11716 6322 11744 6802
rect 11900 6458 11928 6802
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11796 6384 11848 6390
rect 11796 6326 11848 6332
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11808 6202 11836 6326
rect 11520 6180 11572 6186
rect 11520 6122 11572 6128
rect 11716 6174 11836 6202
rect 11612 6112 11664 6118
rect 11716 6100 11744 6174
rect 11664 6072 11744 6100
rect 11612 6054 11664 6060
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11164 5098 11192 5306
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 10980 4814 11100 4842
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10782 3088 10838 3097
rect 10782 3023 10838 3032
rect 10692 2984 10744 2990
rect 10692 2926 10744 2932
rect 10796 2514 10824 3023
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10888 2553 10916 2790
rect 10980 2650 11008 4814
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 11072 3058 11100 4694
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 4010 11192 4422
rect 11152 4004 11204 4010
rect 11152 3946 11204 3952
rect 11164 3126 11192 3946
rect 11256 3534 11284 5714
rect 11518 5672 11574 5681
rect 11518 5607 11574 5616
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 11348 4758 11376 5510
rect 11532 5166 11560 5607
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11348 4622 11376 4694
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 10874 2544 10930 2553
rect 10784 2508 10836 2514
rect 10874 2479 10930 2488
rect 10784 2450 10836 2456
rect 11072 2446 11100 2994
rect 11164 2446 11192 3062
rect 11532 2922 11560 5102
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 11624 4282 11652 4490
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11716 4162 11744 6072
rect 12176 5846 12204 7482
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12268 6798 12296 7278
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12268 6662 12296 6734
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 12164 5704 12216 5710
rect 11886 5672 11942 5681
rect 12164 5646 12216 5652
rect 11886 5607 11942 5616
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11808 4826 11836 4966
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11624 4134 11744 4162
rect 11624 3058 11652 4134
rect 11900 3602 11928 5607
rect 12176 5574 12204 5646
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12256 5296 12308 5302
rect 12254 5264 12256 5273
rect 12308 5264 12310 5273
rect 12254 5199 12310 5208
rect 12360 4826 12388 7482
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12452 5234 12480 5510
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 12084 3670 12112 3878
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 12348 3596 12400 3602
rect 12452 3584 12480 5170
rect 12544 4622 12572 8871
rect 12636 6390 12664 9930
rect 12728 9625 12756 10084
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12714 9616 12770 9625
rect 12714 9551 12770 9560
rect 12820 9466 12848 9998
rect 12728 9450 12848 9466
rect 12716 9444 12848 9450
rect 12768 9438 12848 9444
rect 12716 9386 12768 9392
rect 12728 8906 12756 9386
rect 12817 9276 13113 9296
rect 12873 9274 12897 9276
rect 12953 9274 12977 9276
rect 13033 9274 13057 9276
rect 12895 9222 12897 9274
rect 12959 9222 12971 9274
rect 13033 9222 13035 9274
rect 12873 9220 12897 9222
rect 12953 9220 12977 9222
rect 13033 9220 13057 9222
rect 12817 9200 13113 9220
rect 13372 9058 13400 11018
rect 13464 10266 13492 14010
rect 13924 13938 13952 14418
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 13924 13530 13952 13670
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13542 13288 13598 13297
rect 13542 13223 13598 13232
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13556 10198 13584 13223
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13832 12238 13860 12718
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13740 11694 13768 12174
rect 13924 11898 13952 13330
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 14016 12442 14044 13262
rect 14108 12714 14136 13262
rect 14200 13258 14228 13874
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14200 12918 14228 13194
rect 14188 12912 14240 12918
rect 14188 12854 14240 12860
rect 14096 12708 14148 12714
rect 14096 12650 14148 12656
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 14004 11892 14056 11898
rect 14004 11834 14056 11840
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13912 11620 13964 11626
rect 13912 11562 13964 11568
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13544 10192 13596 10198
rect 13544 10134 13596 10140
rect 13188 9030 13400 9058
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 12728 8498 12756 8842
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12728 8090 12756 8434
rect 12817 8188 13113 8208
rect 12873 8186 12897 8188
rect 12953 8186 12977 8188
rect 13033 8186 13057 8188
rect 12895 8134 12897 8186
rect 12959 8134 12971 8186
rect 13033 8134 13035 8186
rect 12873 8132 12897 8134
rect 12953 8132 12977 8134
rect 13033 8132 13057 8134
rect 12817 8112 13113 8132
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 13188 7970 13216 9030
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 12728 7942 13216 7970
rect 12728 6458 12756 7942
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13188 7410 13216 7754
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 12817 7100 13113 7120
rect 12873 7098 12897 7100
rect 12953 7098 12977 7100
rect 13033 7098 13057 7100
rect 12895 7046 12897 7098
rect 12959 7046 12971 7098
rect 13033 7046 13035 7098
rect 12873 7044 12897 7046
rect 12953 7044 12977 7046
rect 13033 7044 13057 7046
rect 12817 7024 13113 7044
rect 13188 7002 13216 7346
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12912 6458 12940 6802
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 12624 6384 12676 6390
rect 12624 6326 12676 6332
rect 12636 6254 12664 6326
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12728 6118 12756 6394
rect 13004 6390 13032 6734
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 13096 6322 13124 6734
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12817 6012 13113 6032
rect 12873 6010 12897 6012
rect 12953 6010 12977 6012
rect 13033 6010 13057 6012
rect 12895 5958 12897 6010
rect 12959 5958 12971 6010
rect 13033 5958 13035 6010
rect 12873 5956 12897 5958
rect 12953 5956 12977 5958
rect 13033 5956 13057 5958
rect 12817 5936 13113 5956
rect 12817 4924 13113 4944
rect 12873 4922 12897 4924
rect 12953 4922 12977 4924
rect 13033 4922 13057 4924
rect 12895 4870 12897 4922
rect 12959 4870 12971 4922
rect 13033 4870 13035 4922
rect 12873 4868 12897 4870
rect 12953 4868 12977 4870
rect 13033 4868 13057 4870
rect 12817 4848 13113 4868
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12400 3556 12480 3584
rect 12348 3538 12400 3544
rect 12254 3496 12310 3505
rect 12254 3431 12256 3440
rect 12308 3431 12310 3440
rect 12256 3402 12308 3408
rect 11796 3392 11848 3398
rect 12072 3392 12124 3398
rect 11848 3340 11928 3346
rect 11796 3334 11928 3340
rect 12072 3334 12124 3340
rect 11808 3318 11928 3334
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11244 2916 11296 2922
rect 11244 2858 11296 2864
rect 11520 2916 11572 2922
rect 11520 2858 11572 2864
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11256 1562 11284 2858
rect 11716 2650 11744 3130
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11440 2310 11468 2450
rect 11428 2304 11480 2310
rect 11428 2246 11480 2252
rect 11244 1556 11296 1562
rect 11244 1498 11296 1504
rect 11808 1442 11836 3130
rect 11900 3126 11928 3318
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 11888 2576 11940 2582
rect 11888 2518 11940 2524
rect 11900 2106 11928 2518
rect 11888 2100 11940 2106
rect 11888 2042 11940 2048
rect 10336 1414 10548 1442
rect 11256 1414 11836 1442
rect 10336 480 10364 1414
rect 11256 480 11284 1414
rect 12084 1358 12112 3334
rect 12544 2922 12572 4422
rect 12728 4146 12756 4422
rect 12820 4185 12848 4422
rect 13188 4282 13216 4490
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 12806 4176 12862 4185
rect 12716 4140 12768 4146
rect 12806 4111 12862 4120
rect 12716 4082 12768 4088
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12728 3670 12756 3878
rect 12817 3836 13113 3856
rect 12873 3834 12897 3836
rect 12953 3834 12977 3836
rect 13033 3834 13057 3836
rect 12895 3782 12897 3834
rect 12959 3782 12971 3834
rect 13033 3782 13035 3834
rect 12873 3780 12897 3782
rect 12953 3780 12977 3782
rect 13033 3780 13057 3782
rect 12817 3760 13113 3780
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 13280 3534 13308 8502
rect 13372 8090 13400 8910
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13372 6118 13400 7890
rect 13464 7478 13492 8366
rect 13544 8288 13596 8294
rect 13542 8256 13544 8265
rect 13596 8256 13598 8265
rect 13542 8191 13598 8200
rect 13648 7954 13676 11494
rect 13924 11354 13952 11562
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13740 10606 13768 11290
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13832 10538 13860 11222
rect 14016 11218 14044 11834
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13924 10577 13952 11086
rect 13910 10568 13966 10577
rect 13820 10532 13872 10538
rect 13910 10503 13966 10512
rect 13820 10474 13872 10480
rect 13832 9994 13860 10474
rect 13924 10062 13952 10503
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13924 9654 13952 9998
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 14016 9042 14044 11154
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 13924 8022 13952 8774
rect 14016 8498 14044 8774
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 14002 8256 14058 8265
rect 14002 8191 14058 8200
rect 13912 8016 13964 8022
rect 13912 7958 13964 7964
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13636 7812 13688 7818
rect 13556 7772 13636 7800
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13452 6860 13504 6866
rect 13556 6848 13584 7772
rect 13636 7754 13688 7760
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13832 7274 13860 7686
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13504 6820 13584 6848
rect 13820 6860 13872 6866
rect 13452 6802 13504 6808
rect 13820 6802 13872 6808
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13464 5574 13492 6802
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13556 5642 13584 6258
rect 13740 6254 13768 6394
rect 13832 6322 13860 6802
rect 13910 6488 13966 6497
rect 13910 6423 13966 6432
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13924 6254 13952 6423
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 13636 5636 13688 5642
rect 13636 5578 13688 5584
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13464 5234 13492 5510
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13372 4622 13400 4966
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13464 4078 13492 5170
rect 13648 5166 13676 5578
rect 13740 5370 13768 5714
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 13740 4298 13768 5306
rect 13832 5166 13860 6054
rect 13924 5817 13952 6054
rect 13910 5808 13966 5817
rect 13910 5743 13966 5752
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13648 4270 13768 4298
rect 13648 4214 13676 4270
rect 13636 4208 13688 4214
rect 13636 4150 13688 4156
rect 14016 4128 14044 8191
rect 14108 7206 14136 12310
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 10146 14228 12038
rect 14292 11558 14320 14486
rect 14384 14482 14412 16520
rect 14554 16280 14610 16289
rect 14554 16215 14610 16224
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14464 12708 14516 12714
rect 14464 12650 14516 12656
rect 14476 12238 14504 12650
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14464 12232 14516 12238
rect 14568 12209 14596 16215
rect 15014 15872 15070 15881
rect 15014 15807 15070 15816
rect 14646 15056 14702 15065
rect 14646 14991 14702 15000
rect 14464 12174 14516 12180
rect 14554 12200 14610 12209
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 14292 10266 14320 11154
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14200 10118 14320 10146
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 14200 9722 14228 9930
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14108 6866 14136 7142
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14200 6118 14228 8978
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14096 5840 14148 5846
rect 14096 5782 14148 5788
rect 14108 5370 14136 5782
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14016 4100 14136 4128
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13924 3466 13952 3946
rect 14108 3602 14136 4100
rect 14200 3738 14228 4558
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 13912 3460 13964 3466
rect 13912 3402 13964 3408
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 12532 2916 12584 2922
rect 12532 2858 12584 2864
rect 12817 2748 13113 2768
rect 12873 2746 12897 2748
rect 12953 2746 12977 2748
rect 13033 2746 13057 2748
rect 12895 2694 12897 2746
rect 12959 2694 12971 2746
rect 13033 2694 13035 2746
rect 12873 2692 12897 2694
rect 12953 2692 12977 2694
rect 13033 2692 13057 2694
rect 12817 2672 13113 2692
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 12164 2372 12216 2378
rect 12164 2314 12216 2320
rect 12072 1352 12124 1358
rect 12072 1294 12124 1300
rect 12176 480 12204 2314
rect 13096 480 13124 2382
rect 13924 480 13952 2994
rect 14188 2508 14240 2514
rect 14292 2496 14320 10118
rect 14384 8090 14412 12174
rect 14476 11762 14504 12174
rect 14554 12135 14610 12144
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14476 9194 14504 10610
rect 14568 10554 14596 12135
rect 14660 10674 14688 14991
rect 14740 14000 14792 14006
rect 14740 13942 14792 13948
rect 14924 14000 14976 14006
rect 14924 13942 14976 13948
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14568 10526 14688 10554
rect 14476 9166 14596 9194
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14568 7018 14596 9166
rect 14660 7206 14688 10526
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14568 6990 14688 7018
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 14384 4622 14412 5034
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14476 2514 14504 4762
rect 14568 3942 14596 6054
rect 14660 5846 14688 6990
rect 14648 5840 14700 5846
rect 14648 5782 14700 5788
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14648 2984 14700 2990
rect 14752 2972 14780 13942
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14844 12374 14872 13670
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 14936 11898 14964 13942
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 15028 11830 15056 15807
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15106 12880 15162 12889
rect 15106 12815 15162 12824
rect 15120 12306 15148 12815
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 15016 11824 15068 11830
rect 15016 11766 15068 11772
rect 15028 11354 15056 11766
rect 15212 11370 15240 13806
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 15304 13530 15332 13738
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15304 12306 15332 12718
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15304 11762 15332 12242
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15120 11342 15240 11370
rect 14830 11248 14886 11257
rect 14830 11183 14832 11192
rect 14884 11183 14886 11192
rect 14832 11154 14884 11160
rect 15120 10996 15148 11342
rect 15198 11248 15254 11257
rect 15304 11218 15332 11698
rect 15198 11183 15254 11192
rect 15292 11212 15344 11218
rect 15212 11150 15240 11183
rect 15292 11154 15344 11160
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15120 10968 15240 10996
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14844 10062 14872 10406
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 14844 9518 14872 9998
rect 14936 9761 14964 10542
rect 15106 10296 15162 10305
rect 15106 10231 15162 10240
rect 15120 9897 15148 10231
rect 15106 9888 15162 9897
rect 15106 9823 15162 9832
rect 14922 9752 14978 9761
rect 14922 9687 14978 9696
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 15016 9512 15068 9518
rect 15212 9489 15240 10968
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15198 9480 15254 9489
rect 15016 9454 15068 9460
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14844 8974 14872 9318
rect 15028 9110 15056 9454
rect 15120 9438 15198 9466
rect 15016 9104 15068 9110
rect 15016 9046 15068 9052
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14844 8498 14872 8910
rect 14924 8900 14976 8906
rect 14924 8842 14976 8848
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14844 7886 14872 8434
rect 14936 8294 14964 8842
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14936 7993 14964 8230
rect 14922 7984 14978 7993
rect 14922 7919 14978 7928
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14844 7410 14872 7822
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14936 7290 14964 7919
rect 14844 7262 14964 7290
rect 14844 5370 14872 7262
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 14936 5914 14964 6054
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 15028 5794 15056 9046
rect 15120 8362 15148 9438
rect 15198 9415 15254 9424
rect 15304 9178 15332 9862
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15108 8356 15160 8362
rect 15108 8298 15160 8304
rect 15120 7857 15148 8298
rect 15106 7848 15162 7857
rect 15106 7783 15162 7792
rect 15120 6497 15148 7783
rect 15106 6488 15162 6497
rect 15106 6423 15162 6432
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 14936 5766 15056 5794
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 14844 4010 14872 5102
rect 14936 4826 14964 5766
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 14924 4820 14976 4826
rect 14924 4762 14976 4768
rect 15028 4554 15056 5646
rect 15120 5030 15148 6258
rect 15108 5024 15160 5030
rect 15108 4966 15160 4972
rect 15212 4622 15240 8774
rect 15304 7342 15332 8910
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15016 4548 15068 4554
rect 15016 4490 15068 4496
rect 15028 4282 15056 4490
rect 15016 4276 15068 4282
rect 15016 4218 15068 4224
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 14832 4004 14884 4010
rect 14832 3946 14884 3952
rect 14844 3097 14872 3946
rect 14830 3088 14886 3097
rect 14830 3023 14886 3032
rect 14700 2944 14780 2972
rect 14648 2926 14700 2932
rect 15212 2922 15240 4082
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 14240 2468 14320 2496
rect 14464 2508 14516 2514
rect 14188 2450 14240 2456
rect 14464 2450 14516 2456
rect 14844 480 14872 2858
rect 15304 2582 15332 6598
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 15396 1986 15424 14350
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 16210 14240 16266 14249
rect 15672 13870 15700 14214
rect 15782 14172 16078 14192
rect 16210 14175 16266 14184
rect 15838 14170 15862 14172
rect 15918 14170 15942 14172
rect 15998 14170 16022 14172
rect 15860 14118 15862 14170
rect 15924 14118 15936 14170
rect 15998 14118 16000 14170
rect 15838 14116 15862 14118
rect 15918 14116 15942 14118
rect 15998 14116 16022 14118
rect 15782 14096 16078 14116
rect 16224 14074 16252 14175
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16592 13938 16620 16520
rect 16670 14648 16726 14657
rect 16670 14583 16726 14592
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15488 6746 15516 13126
rect 15580 12986 15608 13330
rect 16118 13288 16174 13297
rect 15660 13252 15712 13258
rect 16118 13223 16174 13232
rect 15660 13194 15712 13200
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15672 12442 15700 13194
rect 15782 13084 16078 13104
rect 15838 13082 15862 13084
rect 15918 13082 15942 13084
rect 15998 13082 16022 13084
rect 15860 13030 15862 13082
rect 15924 13030 15936 13082
rect 15998 13030 16000 13082
rect 15838 13028 15862 13030
rect 15918 13028 15942 13030
rect 15998 13028 16022 13030
rect 15782 13008 16078 13028
rect 15750 12472 15806 12481
rect 15660 12436 15712 12442
rect 15750 12407 15806 12416
rect 15660 12378 15712 12384
rect 15764 12084 15792 12407
rect 15672 12056 15792 12084
rect 15566 11656 15622 11665
rect 15566 11591 15622 11600
rect 15580 11121 15608 11591
rect 15566 11112 15622 11121
rect 15566 11047 15622 11056
rect 15566 10568 15622 10577
rect 15566 10503 15622 10512
rect 15580 8906 15608 10503
rect 15672 9450 15700 12056
rect 15782 11996 16078 12016
rect 15838 11994 15862 11996
rect 15918 11994 15942 11996
rect 15998 11994 16022 11996
rect 15860 11942 15862 11994
rect 15924 11942 15936 11994
rect 15998 11942 16000 11994
rect 15838 11940 15862 11942
rect 15918 11940 15942 11942
rect 15998 11940 16022 11942
rect 15782 11920 16078 11940
rect 15782 10908 16078 10928
rect 15838 10906 15862 10908
rect 15918 10906 15942 10908
rect 15998 10906 16022 10908
rect 15860 10854 15862 10906
rect 15924 10854 15936 10906
rect 15998 10854 16000 10906
rect 15838 10852 15862 10854
rect 15918 10852 15942 10854
rect 15998 10852 16022 10854
rect 15782 10832 16078 10852
rect 16132 10606 16160 13223
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16304 12708 16356 12714
rect 16304 12650 16356 12656
rect 16316 12288 16344 12650
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 16224 12260 16344 12288
rect 16224 10962 16252 12260
rect 16304 12164 16356 12170
rect 16304 12106 16356 12112
rect 16316 12073 16344 12106
rect 16302 12064 16358 12073
rect 16302 11999 16358 12008
rect 16408 11898 16436 12582
rect 16500 12238 16528 12786
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16486 11792 16542 11801
rect 16486 11727 16488 11736
rect 16540 11727 16542 11736
rect 16488 11698 16540 11704
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16224 10934 16344 10962
rect 16210 10840 16266 10849
rect 16210 10775 16212 10784
rect 16264 10775 16266 10784
rect 16212 10746 16264 10752
rect 16316 10690 16344 10934
rect 16224 10662 16344 10690
rect 16120 10600 16172 10606
rect 16224 10577 16252 10662
rect 16304 10600 16356 10606
rect 16120 10542 16172 10548
rect 16210 10568 16266 10577
rect 16304 10542 16356 10548
rect 16210 10503 16266 10512
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16120 10192 16172 10198
rect 16120 10134 16172 10140
rect 15782 9820 16078 9840
rect 15838 9818 15862 9820
rect 15918 9818 15942 9820
rect 15998 9818 16022 9820
rect 15860 9766 15862 9818
rect 15924 9766 15936 9818
rect 15998 9766 16000 9818
rect 15838 9764 15862 9766
rect 15918 9764 15942 9766
rect 15998 9764 16022 9766
rect 15782 9744 16078 9764
rect 16132 9450 16160 10134
rect 15660 9444 15712 9450
rect 15660 9386 15712 9392
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 16224 9058 16252 10202
rect 16316 10130 16344 10542
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16316 9722 16344 10066
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 16316 9178 16344 9658
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16120 9036 16172 9042
rect 16224 9030 16344 9058
rect 16120 8978 16172 8984
rect 15568 8900 15620 8906
rect 15568 8842 15620 8848
rect 15782 8732 16078 8752
rect 15838 8730 15862 8732
rect 15918 8730 15942 8732
rect 15998 8730 16022 8732
rect 15860 8678 15862 8730
rect 15924 8678 15936 8730
rect 15998 8678 16000 8730
rect 15838 8676 15862 8678
rect 15918 8676 15942 8678
rect 15998 8676 16022 8678
rect 15782 8656 16078 8676
rect 16132 8634 16160 8978
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 15568 8560 15620 8566
rect 15568 8502 15620 8508
rect 15580 6866 15608 8502
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15672 7410 15700 7686
rect 15782 7644 16078 7664
rect 15838 7642 15862 7644
rect 15918 7642 15942 7644
rect 15998 7642 16022 7644
rect 15860 7590 15862 7642
rect 15924 7590 15936 7642
rect 15998 7590 16000 7642
rect 15838 7588 15862 7590
rect 15918 7588 15942 7590
rect 15998 7588 16022 7590
rect 15782 7568 16078 7588
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15672 7002 15700 7142
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 16224 6798 16252 8570
rect 16316 7426 16344 9030
rect 16408 7546 16436 11154
rect 16500 10198 16528 11698
rect 16592 10810 16620 12582
rect 16684 11218 16712 14583
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16684 10266 16712 10746
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16488 10192 16540 10198
rect 16580 10192 16632 10198
rect 16488 10134 16540 10140
rect 16578 10160 16580 10169
rect 16632 10160 16634 10169
rect 16578 10095 16634 10104
rect 16486 9888 16542 9897
rect 16486 9823 16542 9832
rect 16500 8838 16528 9823
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16500 8090 16528 8298
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16316 7398 16436 7426
rect 16500 7410 16528 8026
rect 16212 6792 16264 6798
rect 15488 6718 15608 6746
rect 16212 6734 16264 6740
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15488 5370 15516 6054
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15580 4146 15608 6718
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 15782 6556 16078 6576
rect 15838 6554 15862 6556
rect 15918 6554 15942 6556
rect 15998 6554 16022 6556
rect 15860 6502 15862 6554
rect 15924 6502 15936 6554
rect 15998 6502 16000 6554
rect 15838 6500 15862 6502
rect 15918 6500 15942 6502
rect 15998 6500 16022 6502
rect 15782 6480 16078 6500
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15672 4826 15700 6394
rect 15936 6384 15988 6390
rect 15936 6326 15988 6332
rect 15948 6118 15976 6326
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15948 5681 15976 6054
rect 15934 5672 15990 5681
rect 15934 5607 15990 5616
rect 15782 5468 16078 5488
rect 15838 5466 15862 5468
rect 15918 5466 15942 5468
rect 15998 5466 16022 5468
rect 15860 5414 15862 5466
rect 15924 5414 15936 5466
rect 15998 5414 16000 5466
rect 15838 5412 15862 5414
rect 15918 5412 15942 5414
rect 15998 5412 16022 5414
rect 15782 5392 16078 5412
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 15672 4214 15700 4762
rect 15948 4622 15976 5170
rect 16118 5128 16174 5137
rect 16118 5063 16120 5072
rect 16172 5063 16174 5072
rect 16120 5034 16172 5040
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 15782 4380 16078 4400
rect 15838 4378 15862 4380
rect 15918 4378 15942 4380
rect 15998 4378 16022 4380
rect 15860 4326 15862 4378
rect 15924 4326 15936 4378
rect 15998 4326 16000 4378
rect 15838 4324 15862 4326
rect 15918 4324 15942 4326
rect 15998 4324 16022 4326
rect 15782 4304 16078 4324
rect 16224 4282 16252 4966
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 15660 4208 15712 4214
rect 15660 4150 15712 4156
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 16316 4078 16344 6598
rect 16408 6118 16436 7398
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16592 6798 16620 10095
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16684 7410 16712 9318
rect 16776 7546 16804 13262
rect 16868 11694 16896 13262
rect 16960 12986 16988 13330
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17052 12442 17080 14214
rect 17132 14000 17184 14006
rect 17132 13942 17184 13948
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 17144 12374 17172 13942
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 17132 12368 17184 12374
rect 17132 12310 17184 12316
rect 17144 11830 17172 12310
rect 17132 11824 17184 11830
rect 17132 11766 17184 11772
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 16868 11354 16896 11630
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16868 8090 16896 9318
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16960 7342 16988 11018
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 17052 6254 17080 10950
rect 17144 10305 17172 11154
rect 17130 10296 17186 10305
rect 17130 10231 17186 10240
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 17144 8634 17172 8978
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17144 7886 17172 8366
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 15474 3496 15530 3505
rect 15474 3431 15530 3440
rect 15488 3194 15516 3431
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15580 2990 15608 3538
rect 15782 3292 16078 3312
rect 15838 3290 15862 3292
rect 15918 3290 15942 3292
rect 15998 3290 16022 3292
rect 15860 3238 15862 3290
rect 15924 3238 15936 3290
rect 15998 3238 16000 3290
rect 15838 3236 15862 3238
rect 15918 3236 15942 3238
rect 15998 3236 16022 3238
rect 15782 3216 16078 3236
rect 16408 3194 16436 6054
rect 17038 5808 17094 5817
rect 17038 5743 17094 5752
rect 16580 4752 16632 4758
rect 16580 4694 16632 4700
rect 16592 3602 16620 4694
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16684 2990 16712 3878
rect 17052 2990 17080 5743
rect 17144 3738 17172 7822
rect 17132 3732 17184 3738
rect 17132 3674 17184 3680
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 16396 2848 16448 2854
rect 16396 2790 16448 2796
rect 16408 2553 16436 2790
rect 16394 2544 16450 2553
rect 16394 2479 16450 2488
rect 15782 2204 16078 2224
rect 15838 2202 15862 2204
rect 15918 2202 15942 2204
rect 15998 2202 16022 2204
rect 15860 2150 15862 2202
rect 15924 2150 15936 2202
rect 15998 2150 16000 2202
rect 15838 2148 15862 2150
rect 15918 2148 15942 2150
rect 15998 2148 16022 2150
rect 15782 2128 16078 2148
rect 15396 1958 15792 1986
rect 15764 480 15792 1958
rect 16684 480 16712 2926
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17052 1873 17080 2790
rect 17038 1864 17094 1873
rect 17038 1799 17094 1808
rect 17236 1306 17264 13806
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17328 12782 17356 13126
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 17420 11762 17448 14418
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17512 12617 17540 14350
rect 17696 14006 17724 14350
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17498 12608 17554 12617
rect 17498 12543 17554 12552
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17328 9897 17356 11018
rect 17420 10713 17448 11494
rect 17512 10810 17540 12543
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17406 10704 17462 10713
rect 17406 10639 17462 10648
rect 17604 10554 17632 13874
rect 17972 13530 18000 16623
rect 18786 16520 18842 17000
rect 18800 14550 18828 16520
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18052 14340 18104 14346
rect 18052 14282 18104 14288
rect 18064 13870 18092 14282
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 17696 11150 17724 13194
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17788 11286 17816 12786
rect 17776 11280 17828 11286
rect 17776 11222 17828 11228
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17696 10606 17724 11086
rect 17420 10526 17632 10554
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17314 9888 17370 9897
rect 17314 9823 17370 9832
rect 17314 9072 17370 9081
rect 17314 9007 17370 9016
rect 17328 8265 17356 9007
rect 17314 8256 17370 8265
rect 17314 8191 17370 8200
rect 17328 8090 17356 8191
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17316 6180 17368 6186
rect 17316 6122 17368 6128
rect 17328 5778 17356 6122
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 17314 5264 17370 5273
rect 17314 5199 17370 5208
rect 17328 4690 17356 5199
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17420 3942 17448 10526
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17512 9178 17540 10066
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17512 7886 17540 9114
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17604 7410 17632 10406
rect 17696 10266 17724 10542
rect 17788 10470 17816 11222
rect 17880 10674 17908 13330
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17866 10568 17922 10577
rect 17866 10503 17922 10512
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17696 9586 17724 10202
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17880 9194 17908 10503
rect 17972 10198 18000 13466
rect 18144 11620 18196 11626
rect 18144 11562 18196 11568
rect 18052 10532 18104 10538
rect 18052 10474 18104 10480
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17696 9166 17908 9194
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17604 5681 17632 6054
rect 17590 5672 17646 5681
rect 17590 5607 17646 5616
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 17512 5273 17540 5510
rect 17498 5264 17554 5273
rect 17498 5199 17554 5208
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17500 4480 17552 4486
rect 17604 4457 17632 4966
rect 17500 4422 17552 4428
rect 17590 4448 17646 4457
rect 17512 4049 17540 4422
rect 17590 4383 17646 4392
rect 17498 4040 17554 4049
rect 17498 3975 17554 3984
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17512 2281 17540 3334
rect 17604 3097 17632 3878
rect 17590 3088 17646 3097
rect 17696 3058 17724 9166
rect 17868 8560 17920 8566
rect 17868 8502 17920 8508
rect 17880 8265 17908 8502
rect 17866 8256 17922 8265
rect 17866 8191 17922 8200
rect 17972 7342 18000 9862
rect 18064 8430 18092 10474
rect 18156 10441 18184 11562
rect 18142 10432 18198 10441
rect 18142 10367 18198 10376
rect 18326 10296 18382 10305
rect 18326 10231 18382 10240
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 18156 8673 18184 9386
rect 18142 8664 18198 8673
rect 18142 8599 18198 8608
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 18156 7936 18184 8599
rect 18064 7908 18184 7936
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 18064 7154 18092 7908
rect 18142 7848 18198 7857
rect 18142 7783 18144 7792
rect 18196 7783 18198 7792
rect 18144 7754 18196 7760
rect 18236 7472 18288 7478
rect 18234 7440 18236 7449
rect 18288 7440 18290 7449
rect 18234 7375 18290 7384
rect 17972 7126 18092 7154
rect 17972 6390 18000 7126
rect 18050 7032 18106 7041
rect 18050 6967 18106 6976
rect 18064 6730 18092 6967
rect 18052 6724 18104 6730
rect 18052 6666 18104 6672
rect 18234 6488 18290 6497
rect 18234 6423 18236 6432
rect 18288 6423 18290 6432
rect 18236 6394 18288 6400
rect 17960 6384 18012 6390
rect 17960 6326 18012 6332
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17788 5098 17816 6190
rect 18050 6080 18106 6089
rect 18050 6015 18106 6024
rect 18064 5914 18092 6015
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18340 5166 18368 10231
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 17776 5092 17828 5098
rect 17776 5034 17828 5040
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18248 4865 18276 4966
rect 18234 4856 18290 4865
rect 18234 4791 18290 4800
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17880 3641 17908 4422
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 17866 3632 17922 3641
rect 17866 3567 17922 3576
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 17590 3023 17646 3032
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 17592 2304 17644 2310
rect 17498 2272 17554 2281
rect 17592 2246 17644 2252
rect 17498 2207 17554 2216
rect 17604 1465 17632 2246
rect 17590 1456 17646 1465
rect 17590 1391 17646 1400
rect 17236 1278 17632 1306
rect 17604 480 17632 1278
rect 17696 1057 17724 2790
rect 17682 1048 17738 1057
rect 17682 983 17738 992
rect 18064 649 18092 3334
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 18050 640 18106 649
rect 18050 575 18106 584
rect 2778 232 2834 241
rect 2778 167 2834 176
rect 3054 0 3110 480
rect 3974 0 4030 480
rect 4894 0 4950 480
rect 5814 0 5870 480
rect 6734 0 6790 480
rect 7562 0 7618 480
rect 8482 0 8538 480
rect 9402 0 9458 480
rect 10322 0 10378 480
rect 11242 0 11298 480
rect 12162 0 12218 480
rect 13082 0 13138 480
rect 13910 0 13966 480
rect 14830 0 14886 480
rect 15750 0 15806 480
rect 16670 0 16726 480
rect 17590 0 17646 480
rect 18248 241 18276 2790
rect 18340 2689 18368 3878
rect 18326 2680 18382 2689
rect 18326 2615 18382 2624
rect 18524 480 18552 13942
rect 19432 1556 19484 1562
rect 19432 1498 19484 1504
rect 19444 480 19472 1498
rect 18234 232 18290 241
rect 18234 167 18290 176
rect 18510 0 18566 480
rect 19430 0 19486 480
<< via2 >>
rect 4066 16632 4122 16688
rect 2870 15816 2926 15872
rect 1398 7520 1454 7576
rect 1398 4664 1454 4720
rect 2318 12708 2374 12744
rect 2318 12688 2320 12708
rect 2320 12688 2372 12708
rect 2372 12688 2374 12708
rect 2870 13368 2926 13424
rect 3790 15408 3846 15464
rect 3698 15000 3754 15056
rect 3514 14592 3570 14648
rect 3422 13776 3478 13832
rect 3606 14184 3662 14240
rect 2778 9696 2834 9752
rect 2778 7248 2834 7304
rect 1674 4256 1730 4312
rect 1858 3440 1914 3496
rect 2962 8064 3018 8120
rect 2870 5888 2926 5944
rect 2778 3848 2834 3904
rect 3606 11328 3662 11384
rect 3422 10920 3478 10976
rect 3422 10124 3478 10160
rect 3422 10104 3424 10124
rect 3424 10104 3476 10124
rect 3476 10104 3478 10124
rect 3330 9696 3386 9752
rect 3422 8916 3424 8936
rect 3424 8916 3476 8936
rect 3476 8916 3478 8936
rect 3422 8880 3478 8916
rect 3238 7928 3294 7984
rect 3330 6296 3386 6352
rect 17958 16632 18014 16688
rect 3921 14170 3977 14172
rect 4001 14170 4057 14172
rect 4081 14170 4137 14172
rect 4161 14170 4217 14172
rect 3921 14118 3947 14170
rect 3947 14118 3977 14170
rect 4001 14118 4011 14170
rect 4011 14118 4057 14170
rect 4081 14118 4127 14170
rect 4127 14118 4137 14170
rect 4161 14118 4191 14170
rect 4191 14118 4217 14170
rect 3921 14116 3977 14118
rect 4001 14116 4057 14118
rect 4081 14116 4137 14118
rect 4161 14116 4217 14118
rect 4066 13232 4122 13288
rect 3921 13082 3977 13084
rect 4001 13082 4057 13084
rect 4081 13082 4137 13084
rect 4161 13082 4217 13084
rect 3921 13030 3947 13082
rect 3947 13030 3977 13082
rect 4001 13030 4011 13082
rect 4011 13030 4057 13082
rect 4081 13030 4127 13082
rect 4127 13030 4137 13082
rect 4161 13030 4191 13082
rect 4191 13030 4217 13082
rect 3921 13028 3977 13030
rect 4001 13028 4057 13030
rect 4081 13028 4137 13030
rect 4161 13028 4217 13030
rect 4066 12824 4122 12880
rect 3974 12588 3976 12608
rect 3976 12588 4028 12608
rect 4028 12588 4030 12608
rect 3974 12552 4030 12588
rect 3921 11994 3977 11996
rect 4001 11994 4057 11996
rect 4081 11994 4137 11996
rect 4161 11994 4217 11996
rect 3921 11942 3947 11994
rect 3947 11942 3977 11994
rect 4001 11942 4011 11994
rect 4011 11942 4057 11994
rect 4081 11942 4127 11994
rect 4127 11942 4137 11994
rect 4161 11942 4191 11994
rect 4191 11942 4217 11994
rect 3921 11940 3977 11942
rect 4001 11940 4057 11942
rect 4081 11940 4137 11942
rect 4161 11940 4217 11942
rect 4526 11736 4582 11792
rect 3921 10906 3977 10908
rect 4001 10906 4057 10908
rect 4081 10906 4137 10908
rect 4161 10906 4217 10908
rect 3921 10854 3947 10906
rect 3947 10854 3977 10906
rect 4001 10854 4011 10906
rect 4011 10854 4057 10906
rect 4081 10854 4127 10906
rect 4127 10854 4137 10906
rect 4161 10854 4191 10906
rect 4191 10854 4217 10906
rect 3921 10852 3977 10854
rect 4001 10852 4057 10854
rect 4081 10852 4137 10854
rect 4161 10852 4217 10854
rect 3974 10512 4030 10568
rect 3698 10104 3754 10160
rect 3921 9818 3977 9820
rect 4001 9818 4057 9820
rect 4081 9818 4137 9820
rect 4161 9818 4217 9820
rect 3921 9766 3947 9818
rect 3947 9766 3977 9818
rect 4001 9766 4011 9818
rect 4011 9766 4057 9818
rect 4081 9766 4127 9818
rect 4127 9766 4137 9818
rect 4161 9766 4191 9818
rect 4191 9766 4217 9818
rect 3921 9764 3977 9766
rect 4001 9764 4057 9766
rect 4081 9764 4137 9766
rect 4161 9764 4217 9766
rect 4066 9288 4122 9344
rect 3790 9016 3846 9072
rect 3921 8730 3977 8732
rect 4001 8730 4057 8732
rect 4081 8730 4137 8732
rect 4161 8730 4217 8732
rect 3921 8678 3947 8730
rect 3947 8678 3977 8730
rect 4001 8678 4011 8730
rect 4011 8678 4057 8730
rect 4081 8678 4127 8730
rect 4127 8678 4137 8730
rect 4161 8678 4191 8730
rect 4191 8678 4217 8730
rect 3921 8676 3977 8678
rect 4001 8676 4057 8678
rect 4081 8676 4137 8678
rect 4161 8676 4217 8678
rect 3606 8064 3662 8120
rect 3054 5072 3110 5128
rect 3238 3032 3294 3088
rect 2962 1808 3018 1864
rect 3606 7656 3662 7712
rect 4066 8336 4122 8392
rect 3790 7928 3846 7984
rect 3921 7642 3977 7644
rect 4001 7642 4057 7644
rect 4081 7642 4137 7644
rect 4161 7642 4217 7644
rect 3921 7590 3947 7642
rect 3947 7590 3977 7642
rect 4001 7590 4011 7642
rect 4011 7590 4057 7642
rect 4081 7590 4127 7642
rect 4127 7590 4137 7642
rect 4161 7590 4191 7642
rect 4191 7590 4217 7642
rect 3921 7588 3977 7590
rect 4001 7588 4057 7590
rect 4081 7588 4137 7590
rect 4161 7588 4217 7590
rect 3790 7112 3846 7168
rect 6886 14714 6942 14716
rect 6966 14714 7022 14716
rect 7046 14714 7102 14716
rect 7126 14714 7182 14716
rect 6886 14662 6912 14714
rect 6912 14662 6942 14714
rect 6966 14662 6976 14714
rect 6976 14662 7022 14714
rect 7046 14662 7092 14714
rect 7092 14662 7102 14714
rect 7126 14662 7156 14714
rect 7156 14662 7182 14714
rect 6886 14660 6942 14662
rect 6966 14660 7022 14662
rect 7046 14660 7102 14662
rect 7126 14660 7182 14662
rect 4802 9696 4858 9752
rect 3790 6704 3846 6760
rect 3698 6060 3700 6080
rect 3700 6060 3752 6080
rect 3752 6060 3754 6080
rect 3698 6024 3754 6060
rect 3921 6554 3977 6556
rect 4001 6554 4057 6556
rect 4081 6554 4137 6556
rect 4161 6554 4217 6556
rect 3921 6502 3947 6554
rect 3947 6502 3977 6554
rect 4001 6502 4011 6554
rect 4011 6502 4057 6554
rect 4081 6502 4127 6554
rect 4127 6502 4137 6554
rect 4161 6502 4191 6554
rect 4191 6502 4217 6554
rect 3921 6500 3977 6502
rect 4001 6500 4057 6502
rect 4081 6500 4137 6502
rect 4161 6500 4217 6502
rect 4434 6432 4490 6488
rect 3698 5480 3754 5536
rect 3921 5466 3977 5468
rect 4001 5466 4057 5468
rect 4081 5466 4137 5468
rect 4161 5466 4217 5468
rect 3921 5414 3947 5466
rect 3947 5414 3977 5466
rect 4001 5414 4011 5466
rect 4011 5414 4057 5466
rect 4081 5414 4127 5466
rect 4127 5414 4137 5466
rect 4161 5414 4191 5466
rect 4191 5414 4217 5466
rect 3921 5412 3977 5414
rect 4001 5412 4057 5414
rect 4081 5412 4137 5414
rect 4161 5412 4217 5414
rect 6886 13626 6942 13628
rect 6966 13626 7022 13628
rect 7046 13626 7102 13628
rect 7126 13626 7182 13628
rect 6886 13574 6912 13626
rect 6912 13574 6942 13626
rect 6966 13574 6976 13626
rect 6976 13574 7022 13626
rect 7046 13574 7092 13626
rect 7092 13574 7102 13626
rect 7126 13574 7156 13626
rect 7156 13574 7182 13626
rect 6886 13572 6942 13574
rect 6966 13572 7022 13574
rect 7046 13572 7102 13574
rect 7126 13572 7182 13574
rect 6886 12538 6942 12540
rect 6966 12538 7022 12540
rect 7046 12538 7102 12540
rect 7126 12538 7182 12540
rect 6886 12486 6912 12538
rect 6912 12486 6942 12538
rect 6966 12486 6976 12538
rect 6976 12486 7022 12538
rect 7046 12486 7092 12538
rect 7092 12486 7102 12538
rect 7126 12486 7156 12538
rect 7156 12486 7182 12538
rect 6886 12484 6942 12486
rect 6966 12484 7022 12486
rect 7046 12484 7102 12486
rect 7126 12484 7182 12486
rect 6550 12008 6606 12064
rect 6090 11192 6146 11248
rect 5538 10648 5594 10704
rect 4986 7928 5042 7984
rect 3921 4378 3977 4380
rect 4001 4378 4057 4380
rect 4081 4378 4137 4380
rect 4161 4378 4217 4380
rect 3921 4326 3947 4378
rect 3947 4326 3977 4378
rect 4001 4326 4011 4378
rect 4011 4326 4057 4378
rect 4081 4326 4127 4378
rect 4127 4326 4137 4378
rect 4161 4326 4191 4378
rect 4191 4326 4217 4378
rect 3921 4324 3977 4326
rect 4001 4324 4057 4326
rect 4081 4324 4137 4326
rect 4161 4324 4217 4326
rect 3698 2216 3754 2272
rect 3422 1400 3478 1456
rect 4342 4972 4344 4992
rect 4344 4972 4396 4992
rect 4396 4972 4398 4992
rect 4342 4936 4398 4972
rect 5262 6160 5318 6216
rect 5170 5788 5172 5808
rect 5172 5788 5224 5808
rect 5224 5788 5226 5808
rect 5170 5752 5226 5788
rect 3921 3290 3977 3292
rect 4001 3290 4057 3292
rect 4081 3290 4137 3292
rect 4161 3290 4217 3292
rect 3921 3238 3947 3290
rect 3947 3238 3977 3290
rect 4001 3238 4011 3290
rect 4011 3238 4057 3290
rect 4081 3238 4127 3290
rect 4127 3238 4137 3290
rect 4161 3238 4191 3290
rect 4191 3238 4217 3290
rect 3921 3236 3977 3238
rect 4001 3236 4057 3238
rect 4081 3236 4137 3238
rect 4161 3236 4217 3238
rect 4066 2624 4122 2680
rect 3921 2202 3977 2204
rect 4001 2202 4057 2204
rect 4081 2202 4137 2204
rect 4161 2202 4217 2204
rect 3921 2150 3947 2202
rect 3947 2150 3977 2202
rect 4001 2150 4011 2202
rect 4011 2150 4057 2202
rect 4081 2150 4127 2202
rect 4127 2150 4137 2202
rect 4161 2150 4191 2202
rect 4191 2150 4217 2202
rect 3921 2148 3977 2150
rect 4001 2148 4057 2150
rect 4081 2148 4137 2150
rect 4161 2148 4217 2150
rect 3790 992 3846 1048
rect 3330 584 3386 640
rect 5906 6024 5962 6080
rect 6886 11450 6942 11452
rect 6966 11450 7022 11452
rect 7046 11450 7102 11452
rect 7126 11450 7182 11452
rect 6886 11398 6912 11450
rect 6912 11398 6942 11450
rect 6966 11398 6976 11450
rect 6976 11398 7022 11450
rect 7046 11398 7092 11450
rect 7092 11398 7102 11450
rect 7126 11398 7156 11450
rect 7156 11398 7182 11450
rect 6886 11396 6942 11398
rect 6966 11396 7022 11398
rect 7046 11396 7102 11398
rect 7126 11396 7182 11398
rect 6550 9968 6606 10024
rect 6886 10362 6942 10364
rect 6966 10362 7022 10364
rect 7046 10362 7102 10364
rect 7126 10362 7182 10364
rect 6886 10310 6912 10362
rect 6912 10310 6942 10362
rect 6966 10310 6976 10362
rect 6976 10310 7022 10362
rect 7046 10310 7092 10362
rect 7092 10310 7102 10362
rect 7126 10310 7156 10362
rect 7156 10310 7182 10362
rect 6886 10308 6942 10310
rect 6966 10308 7022 10310
rect 7046 10308 7102 10310
rect 7126 10308 7182 10310
rect 6918 10104 6974 10160
rect 7010 9968 7066 10024
rect 7010 9424 7066 9480
rect 6886 9274 6942 9276
rect 6966 9274 7022 9276
rect 7046 9274 7102 9276
rect 7126 9274 7182 9276
rect 6886 9222 6912 9274
rect 6912 9222 6942 9274
rect 6966 9222 6976 9274
rect 6976 9222 7022 9274
rect 7046 9222 7092 9274
rect 7092 9222 7102 9274
rect 7126 9222 7156 9274
rect 7156 9222 7182 9274
rect 6886 9220 6942 9222
rect 6966 9220 7022 9222
rect 7046 9220 7102 9222
rect 7126 9220 7182 9222
rect 7286 9016 7342 9072
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9878 14170
rect 9878 14118 9908 14170
rect 9932 14118 9942 14170
rect 9942 14118 9988 14170
rect 10012 14118 10058 14170
rect 10058 14118 10068 14170
rect 10092 14118 10122 14170
rect 10122 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 9494 13640 9550 13696
rect 7746 12416 7802 12472
rect 8114 12416 8170 12472
rect 8574 12688 8630 12744
rect 6886 8186 6942 8188
rect 6966 8186 7022 8188
rect 7046 8186 7102 8188
rect 7126 8186 7182 8188
rect 6886 8134 6912 8186
rect 6912 8134 6942 8186
rect 6966 8134 6976 8186
rect 6976 8134 7022 8186
rect 7046 8134 7092 8186
rect 7092 8134 7102 8186
rect 7126 8134 7156 8186
rect 7156 8134 7182 8186
rect 6886 8132 6942 8134
rect 6966 8132 7022 8134
rect 7046 8132 7102 8134
rect 7126 8132 7182 8134
rect 7194 7284 7196 7304
rect 7196 7284 7248 7304
rect 7248 7284 7250 7304
rect 7194 7248 7250 7284
rect 6886 7098 6942 7100
rect 6966 7098 7022 7100
rect 7046 7098 7102 7100
rect 7126 7098 7182 7100
rect 6886 7046 6912 7098
rect 6912 7046 6942 7098
rect 6966 7046 6976 7098
rect 6976 7046 7022 7098
rect 7046 7046 7092 7098
rect 7092 7046 7102 7098
rect 7126 7046 7156 7098
rect 7156 7046 7182 7098
rect 6886 7044 6942 7046
rect 6966 7044 7022 7046
rect 7046 7044 7102 7046
rect 7126 7044 7182 7046
rect 6886 6010 6942 6012
rect 6966 6010 7022 6012
rect 7046 6010 7102 6012
rect 7126 6010 7182 6012
rect 6886 5958 6912 6010
rect 6912 5958 6942 6010
rect 6966 5958 6976 6010
rect 6976 5958 7022 6010
rect 7046 5958 7092 6010
rect 7092 5958 7102 6010
rect 7126 5958 7156 6010
rect 7156 5958 7182 6010
rect 6886 5956 6942 5958
rect 6966 5956 7022 5958
rect 7046 5956 7102 5958
rect 7126 5956 7182 5958
rect 6550 5616 6606 5672
rect 6734 4936 6790 4992
rect 6886 4922 6942 4924
rect 6966 4922 7022 4924
rect 7046 4922 7102 4924
rect 7126 4922 7182 4924
rect 6886 4870 6912 4922
rect 6912 4870 6942 4922
rect 6966 4870 6976 4922
rect 6976 4870 7022 4922
rect 7046 4870 7092 4922
rect 7092 4870 7102 4922
rect 7126 4870 7156 4922
rect 7156 4870 7182 4922
rect 6886 4868 6942 4870
rect 6966 4868 7022 4870
rect 7046 4868 7102 4870
rect 7126 4868 7182 4870
rect 6886 3834 6942 3836
rect 6966 3834 7022 3836
rect 7046 3834 7102 3836
rect 7126 3834 7182 3836
rect 6886 3782 6912 3834
rect 6912 3782 6942 3834
rect 6966 3782 6976 3834
rect 6976 3782 7022 3834
rect 7046 3782 7092 3834
rect 7092 3782 7102 3834
rect 7126 3782 7156 3834
rect 7156 3782 7182 3834
rect 6886 3780 6942 3782
rect 6966 3780 7022 3782
rect 7046 3780 7102 3782
rect 7126 3780 7182 3782
rect 6886 2746 6942 2748
rect 6966 2746 7022 2748
rect 7046 2746 7102 2748
rect 7126 2746 7182 2748
rect 6886 2694 6912 2746
rect 6912 2694 6942 2746
rect 6966 2694 6976 2746
rect 6976 2694 7022 2746
rect 7046 2694 7092 2746
rect 7092 2694 7102 2746
rect 7126 2694 7156 2746
rect 7156 2694 7182 2746
rect 6886 2692 6942 2694
rect 6966 2692 7022 2694
rect 7046 2692 7102 2694
rect 7126 2692 7182 2694
rect 8114 12180 8116 12200
rect 8116 12180 8168 12200
rect 8168 12180 8170 12200
rect 8114 12144 8170 12180
rect 8298 12044 8300 12064
rect 8300 12044 8352 12064
rect 8352 12044 8354 12064
rect 7746 8880 7802 8936
rect 8298 12008 8354 12044
rect 8390 9832 8446 9888
rect 8298 9560 8354 9616
rect 7930 5752 7986 5808
rect 8298 6452 8354 6488
rect 8298 6432 8300 6452
rect 8300 6432 8352 6452
rect 8352 6432 8354 6452
rect 9310 12280 9366 12336
rect 8942 10140 8944 10160
rect 8944 10140 8996 10160
rect 8996 10140 8998 10160
rect 8942 10104 8998 10140
rect 8758 9560 8814 9616
rect 8850 7792 8906 7848
rect 8390 6160 8446 6216
rect 10138 13796 10194 13832
rect 10138 13776 10140 13796
rect 10140 13776 10192 13796
rect 10192 13776 10194 13796
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9878 13082
rect 9878 13030 9908 13082
rect 9932 13030 9942 13082
rect 9942 13030 9988 13082
rect 10012 13030 10058 13082
rect 10058 13030 10068 13082
rect 10092 13030 10122 13082
rect 10122 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9878 11994
rect 9878 11942 9908 11994
rect 9932 11942 9942 11994
rect 9942 11942 9988 11994
rect 10012 11942 10058 11994
rect 10058 11942 10068 11994
rect 10092 11942 10122 11994
rect 10122 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 10046 11192 10102 11248
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9878 10906
rect 9878 10854 9908 10906
rect 9932 10854 9942 10906
rect 9942 10854 9988 10906
rect 10012 10854 10058 10906
rect 10058 10854 10068 10906
rect 10092 10854 10122 10906
rect 10122 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 9862 10512 9918 10568
rect 9494 9832 9550 9888
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9878 9818
rect 9878 9766 9908 9818
rect 9932 9766 9942 9818
rect 9942 9766 9988 9818
rect 10012 9766 10058 9818
rect 10058 9766 10068 9818
rect 10092 9766 10122 9818
rect 10122 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 10230 9424 10286 9480
rect 10046 9036 10102 9072
rect 10046 9016 10048 9036
rect 10048 9016 10100 9036
rect 10100 9016 10102 9036
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9878 8730
rect 9878 8678 9908 8730
rect 9932 8678 9942 8730
rect 9942 8678 9988 8730
rect 10012 8678 10058 8730
rect 10058 8678 10068 8730
rect 10092 8678 10122 8730
rect 10122 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 10046 7964 10048 7984
rect 10048 7964 10100 7984
rect 10100 7964 10102 7984
rect 10046 7928 10102 7964
rect 9494 6160 9550 6216
rect 9034 4120 9090 4176
rect 10138 7792 10194 7848
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9878 7642
rect 9878 7590 9908 7642
rect 9932 7590 9942 7642
rect 9942 7590 9988 7642
rect 10012 7590 10058 7642
rect 10058 7590 10068 7642
rect 10092 7590 10122 7642
rect 10122 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 10322 8916 10324 8936
rect 10324 8916 10376 8936
rect 10376 8916 10378 8936
rect 10322 8880 10378 8916
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9878 6554
rect 9878 6502 9908 6554
rect 9932 6502 9942 6554
rect 9942 6502 9988 6554
rect 10012 6502 10058 6554
rect 10058 6502 10068 6554
rect 10092 6502 10122 6554
rect 10122 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9878 5466
rect 9878 5414 9908 5466
rect 9932 5414 9942 5466
rect 9942 5414 9988 5466
rect 10012 5414 10058 5466
rect 10058 5414 10068 5466
rect 10092 5414 10122 5466
rect 10122 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 10138 5072 10194 5128
rect 9862 4684 9918 4720
rect 9862 4664 9864 4684
rect 9864 4664 9916 4684
rect 9916 4664 9918 4684
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9878 4378
rect 9878 4326 9908 4378
rect 9932 4326 9942 4378
rect 9942 4326 9988 4378
rect 10012 4326 10058 4378
rect 10058 4326 10068 4378
rect 10092 4326 10122 4378
rect 10122 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 10414 4664 10470 4720
rect 10690 13676 10692 13696
rect 10692 13676 10744 13696
rect 10744 13676 10746 13696
rect 10690 13640 10746 13676
rect 10690 5752 10746 5808
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9878 3290
rect 9878 3238 9908 3290
rect 9932 3238 9942 3290
rect 9942 3238 9988 3290
rect 10012 3238 10058 3290
rect 10058 3238 10068 3290
rect 10092 3238 10122 3290
rect 10122 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9878 2202
rect 9878 2150 9908 2202
rect 9932 2150 9942 2202
rect 9942 2150 9988 2202
rect 10012 2150 10058 2202
rect 10058 2150 10068 2202
rect 10092 2150 10122 2202
rect 10122 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 10874 9424 10930 9480
rect 14278 15408 14334 15464
rect 12817 14714 12873 14716
rect 12897 14714 12953 14716
rect 12977 14714 13033 14716
rect 13057 14714 13113 14716
rect 12817 14662 12843 14714
rect 12843 14662 12873 14714
rect 12897 14662 12907 14714
rect 12907 14662 12953 14714
rect 12977 14662 13023 14714
rect 13023 14662 13033 14714
rect 13057 14662 13087 14714
rect 13087 14662 13113 14714
rect 12817 14660 12873 14662
rect 12897 14660 12953 14662
rect 12977 14660 13033 14662
rect 13057 14660 13113 14662
rect 11242 13796 11298 13832
rect 11242 13776 11244 13796
rect 11244 13776 11296 13796
rect 11296 13776 11298 13796
rect 11794 13776 11850 13832
rect 11426 9832 11482 9888
rect 11150 8916 11152 8936
rect 11152 8916 11204 8936
rect 11204 8916 11206 8936
rect 11150 8880 11206 8916
rect 11058 7792 11114 7848
rect 12817 13626 12873 13628
rect 12897 13626 12953 13628
rect 12977 13626 13033 13628
rect 13057 13626 13113 13628
rect 12817 13574 12843 13626
rect 12843 13574 12873 13626
rect 12897 13574 12907 13626
rect 12907 13574 12953 13626
rect 12977 13574 13023 13626
rect 13023 13574 13033 13626
rect 13057 13574 13087 13626
rect 13087 13574 13113 13626
rect 12817 13572 12873 13574
rect 12897 13572 12953 13574
rect 12977 13572 13033 13574
rect 13057 13572 13113 13574
rect 11978 11736 12034 11792
rect 11978 11228 11980 11248
rect 11980 11228 12032 11248
rect 12032 11228 12034 11248
rect 11978 11192 12034 11228
rect 12622 10920 12678 10976
rect 12346 9016 12402 9072
rect 13266 12552 13322 12608
rect 12817 12538 12873 12540
rect 12897 12538 12953 12540
rect 12977 12538 13033 12540
rect 13057 12538 13113 12540
rect 12817 12486 12843 12538
rect 12843 12486 12873 12538
rect 12897 12486 12907 12538
rect 12907 12486 12953 12538
rect 12977 12486 13023 12538
rect 13023 12486 13033 12538
rect 13057 12486 13087 12538
rect 13087 12486 13113 12538
rect 12817 12484 12873 12486
rect 12897 12484 12953 12486
rect 12977 12484 13033 12486
rect 13057 12484 13113 12486
rect 12817 11450 12873 11452
rect 12897 11450 12953 11452
rect 12977 11450 13033 11452
rect 13057 11450 13113 11452
rect 12817 11398 12843 11450
rect 12843 11398 12873 11450
rect 12897 11398 12907 11450
rect 12907 11398 12953 11450
rect 12977 11398 13023 11450
rect 13023 11398 13033 11450
rect 13057 11398 13087 11450
rect 13087 11398 13113 11450
rect 12817 11396 12873 11398
rect 12897 11396 12953 11398
rect 12977 11396 13033 11398
rect 13057 11396 13113 11398
rect 13082 10512 13138 10568
rect 12817 10362 12873 10364
rect 12897 10362 12953 10364
rect 12977 10362 13033 10364
rect 13057 10362 13113 10364
rect 12817 10310 12843 10362
rect 12843 10310 12873 10362
rect 12897 10310 12907 10362
rect 12907 10310 12953 10362
rect 12977 10310 13023 10362
rect 13023 10310 13033 10362
rect 13057 10310 13087 10362
rect 13087 10310 13113 10362
rect 12817 10308 12873 10310
rect 12897 10308 12953 10310
rect 12977 10308 13033 10310
rect 13057 10308 13113 10310
rect 12530 8880 12586 8936
rect 10782 3032 10838 3088
rect 11518 5616 11574 5672
rect 10874 2488 10930 2544
rect 11886 5616 11942 5672
rect 12254 5244 12256 5264
rect 12256 5244 12308 5264
rect 12308 5244 12310 5264
rect 12254 5208 12310 5244
rect 12714 9560 12770 9616
rect 12817 9274 12873 9276
rect 12897 9274 12953 9276
rect 12977 9274 13033 9276
rect 13057 9274 13113 9276
rect 12817 9222 12843 9274
rect 12843 9222 12873 9274
rect 12897 9222 12907 9274
rect 12907 9222 12953 9274
rect 12977 9222 13023 9274
rect 13023 9222 13033 9274
rect 13057 9222 13087 9274
rect 13087 9222 13113 9274
rect 12817 9220 12873 9222
rect 12897 9220 12953 9222
rect 12977 9220 13033 9222
rect 13057 9220 13113 9222
rect 13542 13232 13598 13288
rect 12817 8186 12873 8188
rect 12897 8186 12953 8188
rect 12977 8186 13033 8188
rect 13057 8186 13113 8188
rect 12817 8134 12843 8186
rect 12843 8134 12873 8186
rect 12897 8134 12907 8186
rect 12907 8134 12953 8186
rect 12977 8134 13023 8186
rect 13023 8134 13033 8186
rect 13057 8134 13087 8186
rect 13087 8134 13113 8186
rect 12817 8132 12873 8134
rect 12897 8132 12953 8134
rect 12977 8132 13033 8134
rect 13057 8132 13113 8134
rect 12817 7098 12873 7100
rect 12897 7098 12953 7100
rect 12977 7098 13033 7100
rect 13057 7098 13113 7100
rect 12817 7046 12843 7098
rect 12843 7046 12873 7098
rect 12897 7046 12907 7098
rect 12907 7046 12953 7098
rect 12977 7046 13023 7098
rect 13023 7046 13033 7098
rect 13057 7046 13087 7098
rect 13087 7046 13113 7098
rect 12817 7044 12873 7046
rect 12897 7044 12953 7046
rect 12977 7044 13033 7046
rect 13057 7044 13113 7046
rect 12817 6010 12873 6012
rect 12897 6010 12953 6012
rect 12977 6010 13033 6012
rect 13057 6010 13113 6012
rect 12817 5958 12843 6010
rect 12843 5958 12873 6010
rect 12897 5958 12907 6010
rect 12907 5958 12953 6010
rect 12977 5958 13023 6010
rect 13023 5958 13033 6010
rect 13057 5958 13087 6010
rect 13087 5958 13113 6010
rect 12817 5956 12873 5958
rect 12897 5956 12953 5958
rect 12977 5956 13033 5958
rect 13057 5956 13113 5958
rect 12817 4922 12873 4924
rect 12897 4922 12953 4924
rect 12977 4922 13033 4924
rect 13057 4922 13113 4924
rect 12817 4870 12843 4922
rect 12843 4870 12873 4922
rect 12897 4870 12907 4922
rect 12907 4870 12953 4922
rect 12977 4870 13023 4922
rect 13023 4870 13033 4922
rect 13057 4870 13087 4922
rect 13087 4870 13113 4922
rect 12817 4868 12873 4870
rect 12897 4868 12953 4870
rect 12977 4868 13033 4870
rect 13057 4868 13113 4870
rect 12254 3460 12310 3496
rect 12254 3440 12256 3460
rect 12256 3440 12308 3460
rect 12308 3440 12310 3460
rect 12806 4120 12862 4176
rect 12817 3834 12873 3836
rect 12897 3834 12953 3836
rect 12977 3834 13033 3836
rect 13057 3834 13113 3836
rect 12817 3782 12843 3834
rect 12843 3782 12873 3834
rect 12897 3782 12907 3834
rect 12907 3782 12953 3834
rect 12977 3782 13023 3834
rect 13023 3782 13033 3834
rect 13057 3782 13087 3834
rect 13087 3782 13113 3834
rect 12817 3780 12873 3782
rect 12897 3780 12953 3782
rect 12977 3780 13033 3782
rect 13057 3780 13113 3782
rect 13542 8236 13544 8256
rect 13544 8236 13596 8256
rect 13596 8236 13598 8256
rect 13542 8200 13598 8236
rect 13910 10512 13966 10568
rect 14002 8200 14058 8256
rect 13910 6432 13966 6488
rect 13910 5752 13966 5808
rect 14554 16224 14610 16280
rect 15014 15816 15070 15872
rect 14646 15000 14702 15056
rect 12817 2746 12873 2748
rect 12897 2746 12953 2748
rect 12977 2746 13033 2748
rect 13057 2746 13113 2748
rect 12817 2694 12843 2746
rect 12843 2694 12873 2746
rect 12897 2694 12907 2746
rect 12907 2694 12953 2746
rect 12977 2694 13023 2746
rect 13023 2694 13033 2746
rect 13057 2694 13087 2746
rect 13087 2694 13113 2746
rect 12817 2692 12873 2694
rect 12897 2692 12953 2694
rect 12977 2692 13033 2694
rect 13057 2692 13113 2694
rect 14554 12144 14610 12200
rect 15106 12824 15162 12880
rect 14830 11212 14886 11248
rect 14830 11192 14832 11212
rect 14832 11192 14884 11212
rect 14884 11192 14886 11212
rect 15198 11192 15254 11248
rect 15106 10240 15162 10296
rect 15106 9832 15162 9888
rect 14922 9696 14978 9752
rect 14922 7928 14978 7984
rect 15198 9424 15254 9480
rect 15106 7792 15162 7848
rect 15106 6432 15162 6488
rect 14830 3032 14886 3088
rect 16210 14184 16266 14240
rect 15782 14170 15838 14172
rect 15862 14170 15918 14172
rect 15942 14170 15998 14172
rect 16022 14170 16078 14172
rect 15782 14118 15808 14170
rect 15808 14118 15838 14170
rect 15862 14118 15872 14170
rect 15872 14118 15918 14170
rect 15942 14118 15988 14170
rect 15988 14118 15998 14170
rect 16022 14118 16052 14170
rect 16052 14118 16078 14170
rect 15782 14116 15838 14118
rect 15862 14116 15918 14118
rect 15942 14116 15998 14118
rect 16022 14116 16078 14118
rect 16670 14592 16726 14648
rect 16118 13232 16174 13288
rect 15782 13082 15838 13084
rect 15862 13082 15918 13084
rect 15942 13082 15998 13084
rect 16022 13082 16078 13084
rect 15782 13030 15808 13082
rect 15808 13030 15838 13082
rect 15862 13030 15872 13082
rect 15872 13030 15918 13082
rect 15942 13030 15988 13082
rect 15988 13030 15998 13082
rect 16022 13030 16052 13082
rect 16052 13030 16078 13082
rect 15782 13028 15838 13030
rect 15862 13028 15918 13030
rect 15942 13028 15998 13030
rect 16022 13028 16078 13030
rect 15750 12416 15806 12472
rect 15566 11600 15622 11656
rect 15566 11056 15622 11112
rect 15566 10512 15622 10568
rect 15782 11994 15838 11996
rect 15862 11994 15918 11996
rect 15942 11994 15998 11996
rect 16022 11994 16078 11996
rect 15782 11942 15808 11994
rect 15808 11942 15838 11994
rect 15862 11942 15872 11994
rect 15872 11942 15918 11994
rect 15942 11942 15988 11994
rect 15988 11942 15998 11994
rect 16022 11942 16052 11994
rect 16052 11942 16078 11994
rect 15782 11940 15838 11942
rect 15862 11940 15918 11942
rect 15942 11940 15998 11942
rect 16022 11940 16078 11942
rect 15782 10906 15838 10908
rect 15862 10906 15918 10908
rect 15942 10906 15998 10908
rect 16022 10906 16078 10908
rect 15782 10854 15808 10906
rect 15808 10854 15838 10906
rect 15862 10854 15872 10906
rect 15872 10854 15918 10906
rect 15942 10854 15988 10906
rect 15988 10854 15998 10906
rect 16022 10854 16052 10906
rect 16052 10854 16078 10906
rect 15782 10852 15838 10854
rect 15862 10852 15918 10854
rect 15942 10852 15998 10854
rect 16022 10852 16078 10854
rect 16302 12008 16358 12064
rect 16486 11756 16542 11792
rect 16486 11736 16488 11756
rect 16488 11736 16540 11756
rect 16540 11736 16542 11756
rect 16210 10804 16266 10840
rect 16210 10784 16212 10804
rect 16212 10784 16264 10804
rect 16264 10784 16266 10804
rect 16210 10512 16266 10568
rect 15782 9818 15838 9820
rect 15862 9818 15918 9820
rect 15942 9818 15998 9820
rect 16022 9818 16078 9820
rect 15782 9766 15808 9818
rect 15808 9766 15838 9818
rect 15862 9766 15872 9818
rect 15872 9766 15918 9818
rect 15942 9766 15988 9818
rect 15988 9766 15998 9818
rect 16022 9766 16052 9818
rect 16052 9766 16078 9818
rect 15782 9764 15838 9766
rect 15862 9764 15918 9766
rect 15942 9764 15998 9766
rect 16022 9764 16078 9766
rect 15782 8730 15838 8732
rect 15862 8730 15918 8732
rect 15942 8730 15998 8732
rect 16022 8730 16078 8732
rect 15782 8678 15808 8730
rect 15808 8678 15838 8730
rect 15862 8678 15872 8730
rect 15872 8678 15918 8730
rect 15942 8678 15988 8730
rect 15988 8678 15998 8730
rect 16022 8678 16052 8730
rect 16052 8678 16078 8730
rect 15782 8676 15838 8678
rect 15862 8676 15918 8678
rect 15942 8676 15998 8678
rect 16022 8676 16078 8678
rect 15782 7642 15838 7644
rect 15862 7642 15918 7644
rect 15942 7642 15998 7644
rect 16022 7642 16078 7644
rect 15782 7590 15808 7642
rect 15808 7590 15838 7642
rect 15862 7590 15872 7642
rect 15872 7590 15918 7642
rect 15942 7590 15988 7642
rect 15988 7590 15998 7642
rect 16022 7590 16052 7642
rect 16052 7590 16078 7642
rect 15782 7588 15838 7590
rect 15862 7588 15918 7590
rect 15942 7588 15998 7590
rect 16022 7588 16078 7590
rect 16578 10140 16580 10160
rect 16580 10140 16632 10160
rect 16632 10140 16634 10160
rect 16578 10104 16634 10140
rect 16486 9832 16542 9888
rect 15782 6554 15838 6556
rect 15862 6554 15918 6556
rect 15942 6554 15998 6556
rect 16022 6554 16078 6556
rect 15782 6502 15808 6554
rect 15808 6502 15838 6554
rect 15862 6502 15872 6554
rect 15872 6502 15918 6554
rect 15942 6502 15988 6554
rect 15988 6502 15998 6554
rect 16022 6502 16052 6554
rect 16052 6502 16078 6554
rect 15782 6500 15838 6502
rect 15862 6500 15918 6502
rect 15942 6500 15998 6502
rect 16022 6500 16078 6502
rect 15934 5616 15990 5672
rect 15782 5466 15838 5468
rect 15862 5466 15918 5468
rect 15942 5466 15998 5468
rect 16022 5466 16078 5468
rect 15782 5414 15808 5466
rect 15808 5414 15838 5466
rect 15862 5414 15872 5466
rect 15872 5414 15918 5466
rect 15942 5414 15988 5466
rect 15988 5414 15998 5466
rect 16022 5414 16052 5466
rect 16052 5414 16078 5466
rect 15782 5412 15838 5414
rect 15862 5412 15918 5414
rect 15942 5412 15998 5414
rect 16022 5412 16078 5414
rect 16118 5092 16174 5128
rect 16118 5072 16120 5092
rect 16120 5072 16172 5092
rect 16172 5072 16174 5092
rect 15782 4378 15838 4380
rect 15862 4378 15918 4380
rect 15942 4378 15998 4380
rect 16022 4378 16078 4380
rect 15782 4326 15808 4378
rect 15808 4326 15838 4378
rect 15862 4326 15872 4378
rect 15872 4326 15918 4378
rect 15942 4326 15988 4378
rect 15988 4326 15998 4378
rect 16022 4326 16052 4378
rect 16052 4326 16078 4378
rect 15782 4324 15838 4326
rect 15862 4324 15918 4326
rect 15942 4324 15998 4326
rect 16022 4324 16078 4326
rect 17130 10240 17186 10296
rect 15474 3440 15530 3496
rect 15782 3290 15838 3292
rect 15862 3290 15918 3292
rect 15942 3290 15998 3292
rect 16022 3290 16078 3292
rect 15782 3238 15808 3290
rect 15808 3238 15838 3290
rect 15862 3238 15872 3290
rect 15872 3238 15918 3290
rect 15942 3238 15988 3290
rect 15988 3238 15998 3290
rect 16022 3238 16052 3290
rect 16052 3238 16078 3290
rect 15782 3236 15838 3238
rect 15862 3236 15918 3238
rect 15942 3236 15998 3238
rect 16022 3236 16078 3238
rect 17038 5752 17094 5808
rect 16394 2488 16450 2544
rect 15782 2202 15838 2204
rect 15862 2202 15918 2204
rect 15942 2202 15998 2204
rect 16022 2202 16078 2204
rect 15782 2150 15808 2202
rect 15808 2150 15838 2202
rect 15862 2150 15872 2202
rect 15872 2150 15918 2202
rect 15942 2150 15988 2202
rect 15988 2150 15998 2202
rect 16022 2150 16052 2202
rect 16052 2150 16078 2202
rect 15782 2148 15838 2150
rect 15862 2148 15918 2150
rect 15942 2148 15998 2150
rect 16022 2148 16078 2150
rect 17038 1808 17094 1864
rect 17498 12552 17554 12608
rect 17406 10648 17462 10704
rect 17314 9832 17370 9888
rect 17314 9016 17370 9072
rect 17314 8200 17370 8256
rect 17314 5208 17370 5264
rect 17866 10512 17922 10568
rect 17590 5616 17646 5672
rect 17498 5208 17554 5264
rect 17590 4392 17646 4448
rect 17498 3984 17554 4040
rect 17590 3032 17646 3088
rect 17866 8200 17922 8256
rect 18142 10376 18198 10432
rect 18326 10240 18382 10296
rect 18142 8608 18198 8664
rect 18142 7812 18198 7848
rect 18142 7792 18144 7812
rect 18144 7792 18196 7812
rect 18196 7792 18198 7812
rect 18234 7420 18236 7440
rect 18236 7420 18288 7440
rect 18288 7420 18290 7440
rect 18234 7384 18290 7420
rect 18050 6976 18106 7032
rect 18234 6452 18290 6488
rect 18234 6432 18236 6452
rect 18236 6432 18288 6452
rect 18288 6432 18290 6452
rect 18050 6024 18106 6080
rect 18234 4800 18290 4856
rect 17866 3576 17922 3632
rect 17498 2216 17554 2272
rect 17590 1400 17646 1456
rect 17682 992 17738 1048
rect 18050 584 18106 640
rect 2778 176 2834 232
rect 18326 2624 18382 2680
rect 18234 176 18290 232
<< metal3 >>
rect 0 16690 480 16720
rect 4061 16690 4127 16693
rect 0 16688 4127 16690
rect 0 16632 4066 16688
rect 4122 16632 4127 16688
rect 0 16630 4127 16632
rect 0 16600 480 16630
rect 4061 16627 4127 16630
rect 17953 16690 18019 16693
rect 19520 16690 20000 16720
rect 17953 16688 20000 16690
rect 17953 16632 17958 16688
rect 18014 16632 20000 16688
rect 17953 16630 20000 16632
rect 17953 16627 18019 16630
rect 19520 16600 20000 16630
rect 0 16282 480 16312
rect 4654 16282 4660 16284
rect 0 16222 4660 16282
rect 0 16192 480 16222
rect 4654 16220 4660 16222
rect 4724 16220 4730 16284
rect 14549 16282 14615 16285
rect 19520 16282 20000 16312
rect 14549 16280 20000 16282
rect 14549 16224 14554 16280
rect 14610 16224 20000 16280
rect 14549 16222 20000 16224
rect 14549 16219 14615 16222
rect 19520 16192 20000 16222
rect 0 15874 480 15904
rect 2865 15874 2931 15877
rect 0 15872 2931 15874
rect 0 15816 2870 15872
rect 2926 15816 2931 15872
rect 0 15814 2931 15816
rect 0 15784 480 15814
rect 2865 15811 2931 15814
rect 15009 15874 15075 15877
rect 19520 15874 20000 15904
rect 15009 15872 20000 15874
rect 15009 15816 15014 15872
rect 15070 15816 20000 15872
rect 15009 15814 20000 15816
rect 15009 15811 15075 15814
rect 19520 15784 20000 15814
rect 0 15466 480 15496
rect 3785 15466 3851 15469
rect 0 15464 3851 15466
rect 0 15408 3790 15464
rect 3846 15408 3851 15464
rect 0 15406 3851 15408
rect 0 15376 480 15406
rect 3785 15403 3851 15406
rect 14273 15466 14339 15469
rect 19520 15466 20000 15496
rect 14273 15464 20000 15466
rect 14273 15408 14278 15464
rect 14334 15408 20000 15464
rect 14273 15406 20000 15408
rect 14273 15403 14339 15406
rect 19520 15376 20000 15406
rect 0 15058 480 15088
rect 3693 15058 3759 15061
rect 0 15056 3759 15058
rect 0 15000 3698 15056
rect 3754 15000 3759 15056
rect 0 14998 3759 15000
rect 0 14968 480 14998
rect 3693 14995 3759 14998
rect 14641 15058 14707 15061
rect 19520 15058 20000 15088
rect 14641 15056 20000 15058
rect 14641 15000 14646 15056
rect 14702 15000 20000 15056
rect 14641 14998 20000 15000
rect 14641 14995 14707 14998
rect 19520 14968 20000 14998
rect 6874 14720 7194 14721
rect 0 14650 480 14680
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7194 14720
rect 6874 14655 7194 14656
rect 12805 14720 13125 14721
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 14655 13125 14656
rect 3509 14650 3575 14653
rect 0 14648 3575 14650
rect 0 14592 3514 14648
rect 3570 14592 3575 14648
rect 0 14590 3575 14592
rect 0 14560 480 14590
rect 3509 14587 3575 14590
rect 16665 14650 16731 14653
rect 19520 14650 20000 14680
rect 16665 14648 20000 14650
rect 16665 14592 16670 14648
rect 16726 14592 20000 14648
rect 16665 14590 20000 14592
rect 16665 14587 16731 14590
rect 19520 14560 20000 14590
rect 0 14242 480 14272
rect 3601 14242 3667 14245
rect 0 14240 3667 14242
rect 0 14184 3606 14240
rect 3662 14184 3667 14240
rect 0 14182 3667 14184
rect 0 14152 480 14182
rect 3601 14179 3667 14182
rect 16205 14242 16271 14245
rect 19520 14242 20000 14272
rect 16205 14240 20000 14242
rect 16205 14184 16210 14240
rect 16266 14184 20000 14240
rect 16205 14182 20000 14184
rect 16205 14179 16271 14182
rect 3909 14176 4229 14177
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 14111 4229 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 15770 14176 16090 14177
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 19520 14152 20000 14182
rect 15770 14111 16090 14112
rect 0 13834 480 13864
rect 3417 13834 3483 13837
rect 0 13832 3483 13834
rect 0 13776 3422 13832
rect 3478 13776 3483 13832
rect 0 13774 3483 13776
rect 0 13744 480 13774
rect 3417 13771 3483 13774
rect 10133 13834 10199 13837
rect 11237 13834 11303 13837
rect 10133 13832 11303 13834
rect 10133 13776 10138 13832
rect 10194 13776 11242 13832
rect 11298 13776 11303 13832
rect 10133 13774 11303 13776
rect 10133 13771 10199 13774
rect 11237 13771 11303 13774
rect 11789 13834 11855 13837
rect 19520 13834 20000 13864
rect 11789 13832 20000 13834
rect 11789 13776 11794 13832
rect 11850 13776 20000 13832
rect 11789 13774 20000 13776
rect 11789 13771 11855 13774
rect 19520 13744 20000 13774
rect 9489 13698 9555 13701
rect 10685 13698 10751 13701
rect 9489 13696 10751 13698
rect 9489 13640 9494 13696
rect 9550 13640 10690 13696
rect 10746 13640 10751 13696
rect 9489 13638 10751 13640
rect 9489 13635 9555 13638
rect 10685 13635 10751 13638
rect 6874 13632 7194 13633
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7194 13632
rect 6874 13567 7194 13568
rect 12805 13632 13125 13633
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 13567 13125 13568
rect 0 13426 480 13456
rect 2865 13426 2931 13429
rect 0 13424 2931 13426
rect 0 13368 2870 13424
rect 2926 13368 2931 13424
rect 0 13366 2931 13368
rect 0 13336 480 13366
rect 2865 13363 2931 13366
rect 4061 13290 4127 13293
rect 13537 13290 13603 13293
rect 4061 13288 13603 13290
rect 4061 13232 4066 13288
rect 4122 13232 13542 13288
rect 13598 13232 13603 13288
rect 4061 13230 13603 13232
rect 4061 13227 4127 13230
rect 13537 13227 13603 13230
rect 16113 13290 16179 13293
rect 19520 13290 20000 13320
rect 16113 13288 20000 13290
rect 16113 13232 16118 13288
rect 16174 13232 20000 13288
rect 16113 13230 20000 13232
rect 16113 13227 16179 13230
rect 19520 13200 20000 13230
rect 3909 13088 4229 13089
rect 0 13018 480 13048
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 13023 4229 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 15770 13088 16090 13089
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 13023 16090 13024
rect 0 12958 3434 13018
rect 0 12928 480 12958
rect 3374 12882 3434 12958
rect 4061 12882 4127 12885
rect 3374 12880 4127 12882
rect 3374 12824 4066 12880
rect 4122 12824 4127 12880
rect 3374 12822 4127 12824
rect 4061 12819 4127 12822
rect 15101 12882 15167 12885
rect 19520 12882 20000 12912
rect 15101 12880 20000 12882
rect 15101 12824 15106 12880
rect 15162 12824 20000 12880
rect 15101 12822 20000 12824
rect 15101 12819 15167 12822
rect 19520 12792 20000 12822
rect 2313 12746 2379 12749
rect 8569 12746 8635 12749
rect 2313 12744 8635 12746
rect 2313 12688 2318 12744
rect 2374 12688 8574 12744
rect 8630 12688 8635 12744
rect 2313 12686 8635 12688
rect 2313 12683 2379 12686
rect 8569 12683 8635 12686
rect 0 12610 480 12640
rect 3969 12610 4035 12613
rect 0 12608 4035 12610
rect 0 12552 3974 12608
rect 4030 12552 4035 12608
rect 0 12550 4035 12552
rect 0 12520 480 12550
rect 3969 12547 4035 12550
rect 13261 12610 13327 12613
rect 17493 12610 17559 12613
rect 13261 12608 17559 12610
rect 13261 12552 13266 12608
rect 13322 12552 17498 12608
rect 17554 12552 17559 12608
rect 13261 12550 17559 12552
rect 13261 12547 13327 12550
rect 17493 12547 17559 12550
rect 6874 12544 7194 12545
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7194 12544
rect 6874 12479 7194 12480
rect 12805 12544 13125 12545
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 12479 13125 12480
rect 7741 12474 7807 12477
rect 8109 12474 8175 12477
rect 7741 12472 8175 12474
rect 7741 12416 7746 12472
rect 7802 12416 8114 12472
rect 8170 12416 8175 12472
rect 7741 12414 8175 12416
rect 7741 12411 7807 12414
rect 8109 12411 8175 12414
rect 15745 12474 15811 12477
rect 19520 12474 20000 12504
rect 15745 12472 20000 12474
rect 15745 12416 15750 12472
rect 15806 12416 20000 12472
rect 15745 12414 20000 12416
rect 15745 12411 15811 12414
rect 19520 12384 20000 12414
rect 2638 12338 2882 12372
rect 9305 12338 9371 12341
rect 2638 12336 9371 12338
rect 2638 12312 9310 12336
rect 0 12202 480 12232
rect 2638 12202 2698 12312
rect 2822 12280 9310 12312
rect 9366 12280 9371 12336
rect 2822 12278 9371 12280
rect 9305 12275 9371 12278
rect 0 12142 2698 12202
rect 8109 12202 8175 12205
rect 14549 12202 14615 12205
rect 8109 12200 14615 12202
rect 8109 12144 8114 12200
rect 8170 12144 14554 12200
rect 14610 12144 14615 12200
rect 8109 12142 14615 12144
rect 0 12112 480 12142
rect 8109 12139 8175 12142
rect 14549 12139 14615 12142
rect 6545 12066 6611 12069
rect 8293 12066 8359 12069
rect 6545 12064 8359 12066
rect 6545 12008 6550 12064
rect 6606 12008 8298 12064
rect 8354 12008 8359 12064
rect 6545 12006 8359 12008
rect 6545 12003 6611 12006
rect 8293 12003 8359 12006
rect 16297 12066 16363 12069
rect 19520 12066 20000 12096
rect 16297 12064 20000 12066
rect 16297 12008 16302 12064
rect 16358 12008 20000 12064
rect 16297 12006 20000 12008
rect 16297 12003 16363 12006
rect 3909 12000 4229 12001
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 11935 4229 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 15770 12000 16090 12001
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 19520 11976 20000 12006
rect 15770 11935 16090 11936
rect 0 11794 480 11824
rect 4521 11794 4587 11797
rect 0 11792 4587 11794
rect 0 11736 4526 11792
rect 4582 11736 4587 11792
rect 0 11734 4587 11736
rect 0 11704 480 11734
rect 4521 11731 4587 11734
rect 11973 11794 12039 11797
rect 16481 11794 16547 11797
rect 11973 11792 16547 11794
rect 11973 11736 11978 11792
rect 12034 11736 16486 11792
rect 16542 11736 16547 11792
rect 11973 11734 16547 11736
rect 11973 11731 12039 11734
rect 16481 11731 16547 11734
rect 15561 11658 15627 11661
rect 19520 11658 20000 11688
rect 15561 11656 20000 11658
rect 15561 11600 15566 11656
rect 15622 11600 20000 11656
rect 15561 11598 20000 11600
rect 15561 11595 15627 11598
rect 19520 11568 20000 11598
rect 6874 11456 7194 11457
rect 0 11386 480 11416
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7194 11456
rect 6874 11391 7194 11392
rect 12805 11456 13125 11457
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 11391 13125 11392
rect 3601 11386 3667 11389
rect 0 11384 3667 11386
rect 0 11328 3606 11384
rect 3662 11328 3667 11384
rect 0 11326 3667 11328
rect 0 11296 480 11326
rect 3601 11323 3667 11326
rect 6085 11250 6151 11253
rect 9622 11250 9628 11252
rect 6085 11248 9628 11250
rect 6085 11192 6090 11248
rect 6146 11192 9628 11248
rect 6085 11190 9628 11192
rect 6085 11187 6151 11190
rect 9622 11188 9628 11190
rect 9692 11250 9698 11252
rect 10041 11250 10107 11253
rect 9692 11248 10107 11250
rect 9692 11192 10046 11248
rect 10102 11192 10107 11248
rect 9692 11190 10107 11192
rect 9692 11188 9698 11190
rect 10041 11187 10107 11190
rect 11973 11250 12039 11253
rect 14825 11250 14891 11253
rect 11973 11248 14891 11250
rect 11973 11192 11978 11248
rect 12034 11192 14830 11248
rect 14886 11192 14891 11248
rect 11973 11190 14891 11192
rect 11973 11187 12039 11190
rect 14825 11187 14891 11190
rect 15193 11250 15259 11253
rect 19520 11250 20000 11280
rect 15193 11248 20000 11250
rect 15193 11192 15198 11248
rect 15254 11192 20000 11248
rect 15193 11190 20000 11192
rect 15193 11187 15259 11190
rect 19520 11160 20000 11190
rect 15561 11114 15627 11117
rect 15150 11112 15627 11114
rect 15150 11056 15566 11112
rect 15622 11056 15627 11112
rect 15150 11054 15627 11056
rect 0 10978 480 11008
rect 3417 10978 3483 10981
rect 0 10976 3483 10978
rect 0 10920 3422 10976
rect 3478 10920 3483 10976
rect 0 10918 3483 10920
rect 0 10888 480 10918
rect 3417 10915 3483 10918
rect 12617 10978 12683 10981
rect 15150 10978 15210 11054
rect 15561 11051 15627 11054
rect 12617 10976 15210 10978
rect 12617 10920 12622 10976
rect 12678 10920 15210 10976
rect 12617 10918 15210 10920
rect 12617 10915 12683 10918
rect 3909 10912 4229 10913
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 10847 4229 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 15770 10912 16090 10913
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 10847 16090 10848
rect 16205 10842 16271 10845
rect 19520 10842 20000 10872
rect 16205 10840 20000 10842
rect 16205 10784 16210 10840
rect 16266 10784 20000 10840
rect 16205 10782 20000 10784
rect 16205 10779 16271 10782
rect 19520 10752 20000 10782
rect 5533 10706 5599 10709
rect 17401 10706 17467 10709
rect 5533 10704 17924 10706
rect 5533 10648 5538 10704
rect 5594 10648 17406 10704
rect 17462 10648 17924 10704
rect 5533 10646 17924 10648
rect 5533 10643 5599 10646
rect 17401 10643 17467 10646
rect 0 10570 480 10600
rect 17864 10573 17924 10646
rect 3969 10570 4035 10573
rect 0 10568 4035 10570
rect 0 10512 3974 10568
rect 4030 10512 4035 10568
rect 0 10510 4035 10512
rect 0 10480 480 10510
rect 3969 10507 4035 10510
rect 9622 10508 9628 10572
rect 9692 10570 9698 10572
rect 9857 10570 9923 10573
rect 9692 10568 9923 10570
rect 9692 10512 9862 10568
rect 9918 10512 9923 10568
rect 9692 10510 9923 10512
rect 9692 10508 9698 10510
rect 9857 10507 9923 10510
rect 13077 10570 13143 10573
rect 13905 10570 13971 10573
rect 13077 10568 13971 10570
rect 13077 10512 13082 10568
rect 13138 10512 13910 10568
rect 13966 10512 13971 10568
rect 13077 10510 13971 10512
rect 13077 10507 13143 10510
rect 13905 10507 13971 10510
rect 15561 10570 15627 10573
rect 16205 10570 16271 10573
rect 15561 10568 16271 10570
rect 15561 10512 15566 10568
rect 15622 10512 16210 10568
rect 16266 10512 16271 10568
rect 15561 10510 16271 10512
rect 15561 10507 15627 10510
rect 16205 10507 16271 10510
rect 17861 10568 17927 10573
rect 17861 10512 17866 10568
rect 17922 10512 17927 10568
rect 17861 10507 17927 10512
rect 18137 10434 18203 10437
rect 19520 10434 20000 10464
rect 18137 10432 20000 10434
rect 18137 10376 18142 10432
rect 18198 10376 20000 10432
rect 18137 10374 20000 10376
rect 18137 10371 18203 10374
rect 6874 10368 7194 10369
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7194 10368
rect 6874 10303 7194 10304
rect 12805 10368 13125 10369
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 19520 10344 20000 10374
rect 12805 10303 13125 10304
rect 15101 10298 15167 10301
rect 17125 10298 17191 10301
rect 18321 10298 18387 10301
rect 15101 10296 18387 10298
rect 15101 10240 15106 10296
rect 15162 10240 17130 10296
rect 17186 10240 18326 10296
rect 18382 10240 18387 10296
rect 15101 10238 18387 10240
rect 15101 10235 15167 10238
rect 17125 10235 17191 10238
rect 18321 10235 18387 10238
rect 0 10162 480 10192
rect 3417 10162 3483 10165
rect 3693 10162 3759 10165
rect 6913 10162 6979 10165
rect 0 10160 6979 10162
rect 0 10104 3422 10160
rect 3478 10104 3698 10160
rect 3754 10104 6918 10160
rect 6974 10104 6979 10160
rect 0 10102 6979 10104
rect 0 10072 480 10102
rect 3417 10099 3483 10102
rect 3693 10099 3759 10102
rect 6913 10099 6979 10102
rect 8937 10162 9003 10165
rect 16573 10162 16639 10165
rect 8937 10160 16639 10162
rect 8937 10104 8942 10160
rect 8998 10104 16578 10160
rect 16634 10104 16639 10160
rect 8937 10102 16639 10104
rect 8937 10099 9003 10102
rect 16573 10099 16639 10102
rect 6545 10026 6611 10029
rect 7005 10026 7071 10029
rect 6545 10024 7071 10026
rect 6545 9968 6550 10024
rect 6606 9968 7010 10024
rect 7066 9968 7071 10024
rect 6545 9966 7071 9968
rect 6545 9963 6611 9966
rect 7005 9963 7071 9966
rect 8385 9890 8451 9893
rect 9489 9890 9555 9893
rect 8385 9888 9555 9890
rect 8385 9832 8390 9888
rect 8446 9832 9494 9888
rect 9550 9832 9555 9888
rect 8385 9830 9555 9832
rect 8385 9827 8451 9830
rect 9489 9827 9555 9830
rect 11421 9890 11487 9893
rect 15101 9890 15167 9893
rect 11421 9888 15167 9890
rect 11421 9832 11426 9888
rect 11482 9832 15106 9888
rect 15162 9832 15167 9888
rect 11421 9830 15167 9832
rect 11421 9827 11487 9830
rect 15101 9827 15167 9830
rect 16481 9890 16547 9893
rect 17309 9890 17375 9893
rect 19520 9890 20000 9920
rect 16481 9888 20000 9890
rect 16481 9832 16486 9888
rect 16542 9832 17314 9888
rect 17370 9832 20000 9888
rect 16481 9830 20000 9832
rect 16481 9827 16547 9830
rect 17309 9827 17375 9830
rect 3909 9824 4229 9825
rect 0 9754 480 9784
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 9759 4229 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 15770 9824 16090 9825
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 19520 9800 20000 9830
rect 15770 9759 16090 9760
rect 2773 9754 2839 9757
rect 3325 9754 3391 9757
rect 0 9752 3391 9754
rect 0 9696 2778 9752
rect 2834 9696 3330 9752
rect 3386 9696 3391 9752
rect 0 9694 3391 9696
rect 0 9664 480 9694
rect 2773 9691 2839 9694
rect 3325 9691 3391 9694
rect 4654 9692 4660 9756
rect 4724 9754 4730 9756
rect 4797 9754 4863 9757
rect 14917 9754 14983 9757
rect 4724 9752 4863 9754
rect 4724 9696 4802 9752
rect 4858 9696 4863 9752
rect 4724 9694 4863 9696
rect 4724 9692 4730 9694
rect 4797 9691 4863 9694
rect 10228 9752 14983 9754
rect 10228 9696 14922 9752
rect 14978 9696 14983 9752
rect 10228 9694 14983 9696
rect 8293 9618 8359 9621
rect 8753 9618 8819 9621
rect 10228 9618 10288 9694
rect 14917 9691 14983 9694
rect 12709 9618 12775 9621
rect 8293 9616 10288 9618
rect 8293 9560 8298 9616
rect 8354 9560 8758 9616
rect 8814 9560 10288 9616
rect 8293 9558 10288 9560
rect 12574 9616 12775 9618
rect 12574 9560 12714 9616
rect 12770 9560 12775 9616
rect 12574 9558 12775 9560
rect 8293 9555 8359 9558
rect 8753 9555 8819 9558
rect 6678 9420 6684 9484
rect 6748 9482 6754 9484
rect 7005 9482 7071 9485
rect 6748 9480 7071 9482
rect 6748 9424 7010 9480
rect 7066 9424 7071 9480
rect 6748 9422 7071 9424
rect 6748 9420 6754 9422
rect 7005 9419 7071 9422
rect 10225 9482 10291 9485
rect 10869 9482 10935 9485
rect 10225 9480 10935 9482
rect 10225 9424 10230 9480
rect 10286 9424 10874 9480
rect 10930 9424 10935 9480
rect 10225 9422 10935 9424
rect 10225 9419 10291 9422
rect 10869 9419 10935 9422
rect 0 9346 480 9376
rect 4061 9346 4127 9349
rect 0 9344 4127 9346
rect 0 9288 4066 9344
rect 4122 9288 4127 9344
rect 0 9286 4127 9288
rect 0 9256 480 9286
rect 4061 9283 4127 9286
rect 6874 9280 7194 9281
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7194 9280
rect 6874 9215 7194 9216
rect 3785 9074 3851 9077
rect 4286 9074 4292 9076
rect 3785 9072 4292 9074
rect 3785 9016 3790 9072
rect 3846 9016 4292 9072
rect 3785 9014 4292 9016
rect 3785 9011 3851 9014
rect 4286 9012 4292 9014
rect 4356 9012 4362 9076
rect 7281 9074 7347 9077
rect 10041 9074 10107 9077
rect 12341 9074 12407 9077
rect 7281 9072 12407 9074
rect 7281 9016 7286 9072
rect 7342 9016 10046 9072
rect 10102 9016 12346 9072
rect 12402 9016 12407 9072
rect 7281 9014 12407 9016
rect 7281 9011 7347 9014
rect 10041 9011 10107 9014
rect 12341 9011 12407 9014
rect 0 8938 480 8968
rect 12574 8941 12634 9558
rect 12709 9555 12775 9558
rect 15193 9482 15259 9485
rect 19520 9482 20000 9512
rect 15193 9480 20000 9482
rect 15193 9424 15198 9480
rect 15254 9424 20000 9480
rect 15193 9422 20000 9424
rect 15193 9419 15259 9422
rect 19520 9392 20000 9422
rect 12805 9280 13125 9281
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 9215 13125 9216
rect 17309 9074 17375 9077
rect 19520 9074 20000 9104
rect 17309 9072 20000 9074
rect 17309 9016 17314 9072
rect 17370 9016 20000 9072
rect 17309 9014 20000 9016
rect 17309 9011 17375 9014
rect 19520 8984 20000 9014
rect 3417 8938 3483 8941
rect 7741 8938 7807 8941
rect 0 8936 7807 8938
rect 0 8880 3422 8936
rect 3478 8880 7746 8936
rect 7802 8880 7807 8936
rect 0 8878 7807 8880
rect 0 8848 480 8878
rect 3417 8875 3483 8878
rect 7741 8875 7807 8878
rect 10317 8938 10383 8941
rect 11145 8938 11211 8941
rect 10317 8936 11211 8938
rect 10317 8880 10322 8936
rect 10378 8880 11150 8936
rect 11206 8880 11211 8936
rect 10317 8878 11211 8880
rect 10317 8875 10383 8878
rect 11145 8875 11211 8878
rect 12525 8936 12634 8941
rect 12525 8880 12530 8936
rect 12586 8880 12634 8936
rect 12525 8878 12634 8880
rect 12525 8875 12591 8878
rect 3909 8736 4229 8737
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 8671 4229 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 15770 8736 16090 8737
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15770 8671 16090 8672
rect 18137 8666 18203 8669
rect 19520 8666 20000 8696
rect 18137 8664 20000 8666
rect 18137 8608 18142 8664
rect 18198 8608 20000 8664
rect 18137 8606 20000 8608
rect 18137 8603 18203 8606
rect 19520 8576 20000 8606
rect 0 8394 480 8424
rect 4061 8394 4127 8397
rect 0 8392 4127 8394
rect 0 8336 4066 8392
rect 4122 8336 4127 8392
rect 0 8334 4127 8336
rect 0 8304 480 8334
rect 4061 8331 4127 8334
rect 13537 8258 13603 8261
rect 13997 8258 14063 8261
rect 17309 8258 17375 8261
rect 13537 8256 17375 8258
rect 13537 8200 13542 8256
rect 13598 8200 14002 8256
rect 14058 8200 17314 8256
rect 17370 8200 17375 8256
rect 13537 8198 17375 8200
rect 13537 8195 13603 8198
rect 13997 8195 14063 8198
rect 17309 8195 17375 8198
rect 17861 8258 17927 8261
rect 19520 8258 20000 8288
rect 17861 8256 20000 8258
rect 17861 8200 17866 8256
rect 17922 8200 20000 8256
rect 17861 8198 20000 8200
rect 17861 8195 17927 8198
rect 6874 8192 7194 8193
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7194 8192
rect 6874 8127 7194 8128
rect 12805 8192 13125 8193
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 19520 8168 20000 8198
rect 12805 8127 13125 8128
rect 2957 8122 3023 8125
rect 3601 8122 3667 8125
rect 2957 8120 3986 8122
rect 2957 8064 2962 8120
rect 3018 8064 3606 8120
rect 3662 8064 3986 8120
rect 2957 8062 3986 8064
rect 2957 8059 3023 8062
rect 3601 8059 3667 8062
rect 0 7986 480 8016
rect 3233 7986 3299 7989
rect 3785 7986 3851 7989
rect 0 7984 3299 7986
rect 0 7928 3238 7984
rect 3294 7928 3299 7984
rect 0 7926 3299 7928
rect 0 7896 480 7926
rect 3233 7923 3299 7926
rect 3420 7984 3851 7986
rect 3420 7928 3790 7984
rect 3846 7928 3851 7984
rect 3420 7926 3851 7928
rect 3420 7714 3480 7926
rect 3785 7923 3851 7926
rect 3926 7850 3986 8062
rect 4981 7986 5047 7989
rect 10041 7986 10107 7989
rect 14917 7986 14983 7989
rect 4981 7984 14983 7986
rect 4981 7928 4986 7984
rect 5042 7928 10046 7984
rect 10102 7928 14922 7984
rect 14978 7928 14983 7984
rect 4981 7926 14983 7928
rect 4981 7923 5047 7926
rect 10041 7923 10107 7926
rect 14917 7923 14983 7926
rect 8845 7850 8911 7853
rect 3926 7848 8911 7850
rect 3926 7792 8850 7848
rect 8906 7792 8911 7848
rect 3926 7790 8911 7792
rect 8845 7787 8911 7790
rect 10133 7850 10199 7853
rect 11053 7850 11119 7853
rect 15101 7850 15167 7853
rect 10133 7848 15167 7850
rect 10133 7792 10138 7848
rect 10194 7792 11058 7848
rect 11114 7792 15106 7848
rect 15162 7792 15167 7848
rect 10133 7790 15167 7792
rect 10133 7787 10199 7790
rect 11053 7787 11119 7790
rect 15101 7787 15167 7790
rect 18137 7850 18203 7853
rect 19520 7850 20000 7880
rect 18137 7848 20000 7850
rect 18137 7792 18142 7848
rect 18198 7792 20000 7848
rect 18137 7790 20000 7792
rect 18137 7787 18203 7790
rect 19520 7760 20000 7790
rect 3601 7714 3667 7717
rect 3420 7712 3667 7714
rect 3420 7656 3606 7712
rect 3662 7656 3667 7712
rect 3420 7654 3667 7656
rect 3601 7651 3667 7654
rect 3909 7648 4229 7649
rect 0 7578 480 7608
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 7583 4229 7584
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 15770 7648 16090 7649
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 7583 16090 7584
rect 1393 7578 1459 7581
rect 0 7576 1459 7578
rect 0 7520 1398 7576
rect 1454 7520 1459 7576
rect 0 7518 1459 7520
rect 0 7488 480 7518
rect 1393 7515 1459 7518
rect 18229 7442 18295 7445
rect 19520 7442 20000 7472
rect 18229 7440 20000 7442
rect 18229 7384 18234 7440
rect 18290 7384 20000 7440
rect 18229 7382 20000 7384
rect 18229 7379 18295 7382
rect 19520 7352 20000 7382
rect 2773 7306 2839 7309
rect 6678 7306 6684 7308
rect 2773 7304 6684 7306
rect 2773 7248 2778 7304
rect 2834 7248 6684 7304
rect 2773 7246 6684 7248
rect 2773 7243 2839 7246
rect 6678 7244 6684 7246
rect 6748 7306 6754 7308
rect 7189 7306 7255 7309
rect 6748 7304 7255 7306
rect 6748 7248 7194 7304
rect 7250 7248 7255 7304
rect 6748 7246 7255 7248
rect 6748 7244 6754 7246
rect 7189 7243 7255 7246
rect 0 7170 480 7200
rect 3785 7170 3851 7173
rect 0 7168 3851 7170
rect 0 7112 3790 7168
rect 3846 7112 3851 7168
rect 0 7110 3851 7112
rect 0 7080 480 7110
rect 3785 7107 3851 7110
rect 6874 7104 7194 7105
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7194 7104
rect 6874 7039 7194 7040
rect 12805 7104 13125 7105
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 7039 13125 7040
rect 18045 7034 18111 7037
rect 19520 7034 20000 7064
rect 18045 7032 20000 7034
rect 18045 6976 18050 7032
rect 18106 6976 20000 7032
rect 18045 6974 20000 6976
rect 18045 6971 18111 6974
rect 19520 6944 20000 6974
rect 0 6762 480 6792
rect 3785 6762 3851 6765
rect 0 6760 3851 6762
rect 0 6704 3790 6760
rect 3846 6704 3851 6760
rect 0 6702 3851 6704
rect 0 6672 480 6702
rect 3785 6699 3851 6702
rect 3909 6560 4229 6561
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 6495 4229 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 15770 6560 16090 6561
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 6495 16090 6496
rect 4429 6490 4495 6493
rect 8293 6490 8359 6493
rect 4429 6488 8359 6490
rect 4429 6432 4434 6488
rect 4490 6432 8298 6488
rect 8354 6432 8359 6488
rect 4429 6430 8359 6432
rect 4429 6427 4495 6430
rect 8293 6427 8359 6430
rect 13905 6490 13971 6493
rect 15101 6490 15167 6493
rect 13905 6488 15167 6490
rect 13905 6432 13910 6488
rect 13966 6432 15106 6488
rect 15162 6432 15167 6488
rect 13905 6430 15167 6432
rect 13905 6427 13971 6430
rect 15101 6427 15167 6430
rect 18229 6490 18295 6493
rect 19520 6490 20000 6520
rect 18229 6488 20000 6490
rect 18229 6432 18234 6488
rect 18290 6432 20000 6488
rect 18229 6430 20000 6432
rect 18229 6427 18295 6430
rect 19520 6400 20000 6430
rect 0 6354 480 6384
rect 3325 6354 3391 6357
rect 0 6352 3391 6354
rect 0 6296 3330 6352
rect 3386 6296 3391 6352
rect 0 6294 3391 6296
rect 0 6264 480 6294
rect 3325 6291 3391 6294
rect 5257 6218 5323 6221
rect 8385 6218 8451 6221
rect 9489 6218 9555 6221
rect 5257 6216 9555 6218
rect 5257 6160 5262 6216
rect 5318 6160 8390 6216
rect 8446 6160 9494 6216
rect 9550 6160 9555 6216
rect 5257 6158 9555 6160
rect 5257 6155 5323 6158
rect 8385 6155 8451 6158
rect 9489 6155 9555 6158
rect 3693 6082 3759 6085
rect 5901 6082 5967 6085
rect 3693 6080 5967 6082
rect 3693 6024 3698 6080
rect 3754 6024 5906 6080
rect 5962 6024 5967 6080
rect 3693 6022 5967 6024
rect 3693 6019 3759 6022
rect 5901 6019 5967 6022
rect 18045 6082 18111 6085
rect 19520 6082 20000 6112
rect 18045 6080 20000 6082
rect 18045 6024 18050 6080
rect 18106 6024 20000 6080
rect 18045 6022 20000 6024
rect 18045 6019 18111 6022
rect 6874 6016 7194 6017
rect 0 5946 480 5976
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7194 6016
rect 6874 5951 7194 5952
rect 12805 6016 13125 6017
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 19520 5992 20000 6022
rect 12805 5951 13125 5952
rect 2865 5946 2931 5949
rect 0 5944 2931 5946
rect 0 5888 2870 5944
rect 2926 5888 2931 5944
rect 0 5886 2931 5888
rect 0 5856 480 5886
rect 2865 5883 2931 5886
rect 5165 5810 5231 5813
rect 7925 5810 7991 5813
rect 5165 5808 7991 5810
rect 5165 5752 5170 5808
rect 5226 5752 7930 5808
rect 7986 5752 7991 5808
rect 5165 5750 7991 5752
rect 5165 5747 5231 5750
rect 7925 5747 7991 5750
rect 10685 5810 10751 5813
rect 13905 5810 13971 5813
rect 17033 5810 17099 5813
rect 10685 5808 17099 5810
rect 10685 5752 10690 5808
rect 10746 5752 13910 5808
rect 13966 5752 17038 5808
rect 17094 5752 17099 5808
rect 10685 5750 17099 5752
rect 10685 5747 10751 5750
rect 13905 5747 13971 5750
rect 17033 5747 17099 5750
rect 6545 5674 6611 5677
rect 11513 5674 11579 5677
rect 6545 5672 11579 5674
rect 6545 5616 6550 5672
rect 6606 5616 11518 5672
rect 11574 5616 11579 5672
rect 6545 5614 11579 5616
rect 6545 5611 6611 5614
rect 11513 5611 11579 5614
rect 11881 5674 11947 5677
rect 15929 5674 15995 5677
rect 11881 5672 15995 5674
rect 11881 5616 11886 5672
rect 11942 5616 15934 5672
rect 15990 5616 15995 5672
rect 11881 5614 15995 5616
rect 11881 5611 11947 5614
rect 15929 5611 15995 5614
rect 17585 5674 17651 5677
rect 19520 5674 20000 5704
rect 17585 5672 20000 5674
rect 17585 5616 17590 5672
rect 17646 5616 20000 5672
rect 17585 5614 20000 5616
rect 17585 5611 17651 5614
rect 19520 5584 20000 5614
rect 0 5538 480 5568
rect 3693 5538 3759 5541
rect 0 5536 3759 5538
rect 0 5480 3698 5536
rect 3754 5480 3759 5536
rect 0 5478 3759 5480
rect 0 5448 480 5478
rect 3693 5475 3759 5478
rect 3909 5472 4229 5473
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 5407 4229 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 15770 5472 16090 5473
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 5407 16090 5408
rect 12249 5266 12315 5269
rect 17309 5266 17375 5269
rect 12249 5264 17375 5266
rect 12249 5208 12254 5264
rect 12310 5208 17314 5264
rect 17370 5208 17375 5264
rect 12249 5206 17375 5208
rect 12249 5203 12315 5206
rect 17309 5203 17375 5206
rect 17493 5266 17559 5269
rect 19520 5266 20000 5296
rect 17493 5264 20000 5266
rect 17493 5208 17498 5264
rect 17554 5208 20000 5264
rect 17493 5206 20000 5208
rect 17493 5203 17559 5206
rect 19520 5176 20000 5206
rect 0 5130 480 5160
rect 3049 5130 3115 5133
rect 0 5128 3115 5130
rect 0 5072 3054 5128
rect 3110 5072 3115 5128
rect 0 5070 3115 5072
rect 0 5040 480 5070
rect 3049 5067 3115 5070
rect 10133 5130 10199 5133
rect 16113 5130 16179 5133
rect 10133 5128 16179 5130
rect 10133 5072 10138 5128
rect 10194 5072 16118 5128
rect 16174 5072 16179 5128
rect 10133 5070 16179 5072
rect 10133 5067 10199 5070
rect 16113 5067 16179 5070
rect 4337 4996 4403 4997
rect 4286 4932 4292 4996
rect 4356 4994 4403 4996
rect 6729 4994 6795 4997
rect 4356 4992 6795 4994
rect 4398 4936 6734 4992
rect 6790 4936 6795 4992
rect 4356 4934 6795 4936
rect 4356 4932 4403 4934
rect 4337 4931 4403 4932
rect 6729 4931 6795 4934
rect 6874 4928 7194 4929
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7194 4928
rect 6874 4863 7194 4864
rect 12805 4928 13125 4929
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 4863 13125 4864
rect 18229 4858 18295 4861
rect 19520 4858 20000 4888
rect 18229 4856 20000 4858
rect 18229 4800 18234 4856
rect 18290 4800 20000 4856
rect 18229 4798 20000 4800
rect 18229 4795 18295 4798
rect 19520 4768 20000 4798
rect 0 4722 480 4752
rect 1393 4722 1459 4725
rect 0 4720 1459 4722
rect 0 4664 1398 4720
rect 1454 4664 1459 4720
rect 0 4662 1459 4664
rect 0 4632 480 4662
rect 1393 4659 1459 4662
rect 9857 4722 9923 4725
rect 10409 4722 10475 4725
rect 9857 4720 10475 4722
rect 9857 4664 9862 4720
rect 9918 4664 10414 4720
rect 10470 4664 10475 4720
rect 9857 4662 10475 4664
rect 9857 4659 9923 4662
rect 10409 4659 10475 4662
rect 17585 4450 17651 4453
rect 19520 4450 20000 4480
rect 17585 4448 20000 4450
rect 17585 4392 17590 4448
rect 17646 4392 20000 4448
rect 17585 4390 20000 4392
rect 17585 4387 17651 4390
rect 3909 4384 4229 4385
rect 0 4314 480 4344
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 4319 4229 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 15770 4384 16090 4385
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 19520 4360 20000 4390
rect 15770 4319 16090 4320
rect 1669 4314 1735 4317
rect 0 4312 1735 4314
rect 0 4256 1674 4312
rect 1730 4256 1735 4312
rect 0 4254 1735 4256
rect 0 4224 480 4254
rect 1669 4251 1735 4254
rect 9029 4178 9095 4181
rect 12801 4178 12867 4181
rect 9029 4176 12867 4178
rect 9029 4120 9034 4176
rect 9090 4120 12806 4176
rect 12862 4120 12867 4176
rect 9029 4118 12867 4120
rect 9029 4115 9095 4118
rect 12801 4115 12867 4118
rect 17493 4042 17559 4045
rect 19520 4042 20000 4072
rect 17493 4040 20000 4042
rect 17493 3984 17498 4040
rect 17554 3984 20000 4040
rect 17493 3982 20000 3984
rect 17493 3979 17559 3982
rect 19520 3952 20000 3982
rect 0 3906 480 3936
rect 2773 3906 2839 3909
rect 0 3904 2839 3906
rect 0 3848 2778 3904
rect 2834 3848 2839 3904
rect 0 3846 2839 3848
rect 0 3816 480 3846
rect 2773 3843 2839 3846
rect 6874 3840 7194 3841
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7194 3840
rect 6874 3775 7194 3776
rect 12805 3840 13125 3841
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 3775 13125 3776
rect 17861 3634 17927 3637
rect 19520 3634 20000 3664
rect 17861 3632 20000 3634
rect 17861 3576 17866 3632
rect 17922 3576 20000 3632
rect 17861 3574 20000 3576
rect 17861 3571 17927 3574
rect 19520 3544 20000 3574
rect 0 3498 480 3528
rect 1853 3498 1919 3501
rect 0 3496 1919 3498
rect 0 3440 1858 3496
rect 1914 3440 1919 3496
rect 0 3438 1919 3440
rect 0 3408 480 3438
rect 1853 3435 1919 3438
rect 12249 3498 12315 3501
rect 15469 3498 15535 3501
rect 12249 3496 15535 3498
rect 12249 3440 12254 3496
rect 12310 3440 15474 3496
rect 15530 3440 15535 3496
rect 12249 3438 15535 3440
rect 12249 3435 12315 3438
rect 15469 3435 15535 3438
rect 3909 3296 4229 3297
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 3231 4229 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 15770 3296 16090 3297
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 3231 16090 3232
rect 0 3090 480 3120
rect 3233 3090 3299 3093
rect 0 3088 3299 3090
rect 0 3032 3238 3088
rect 3294 3032 3299 3088
rect 0 3030 3299 3032
rect 0 3000 480 3030
rect 3233 3027 3299 3030
rect 10777 3090 10843 3093
rect 14825 3090 14891 3093
rect 10777 3088 14891 3090
rect 10777 3032 10782 3088
rect 10838 3032 14830 3088
rect 14886 3032 14891 3088
rect 10777 3030 14891 3032
rect 10777 3027 10843 3030
rect 14825 3027 14891 3030
rect 17585 3090 17651 3093
rect 19520 3090 20000 3120
rect 17585 3088 20000 3090
rect 17585 3032 17590 3088
rect 17646 3032 20000 3088
rect 17585 3030 20000 3032
rect 17585 3027 17651 3030
rect 19520 3000 20000 3030
rect 6874 2752 7194 2753
rect 0 2682 480 2712
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7194 2752
rect 6874 2687 7194 2688
rect 12805 2752 13125 2753
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2687 13125 2688
rect 4061 2682 4127 2685
rect 0 2680 4127 2682
rect 0 2624 4066 2680
rect 4122 2624 4127 2680
rect 0 2622 4127 2624
rect 0 2592 480 2622
rect 4061 2619 4127 2622
rect 18321 2682 18387 2685
rect 19520 2682 20000 2712
rect 18321 2680 20000 2682
rect 18321 2624 18326 2680
rect 18382 2624 20000 2680
rect 18321 2622 20000 2624
rect 18321 2619 18387 2622
rect 19520 2592 20000 2622
rect 10869 2546 10935 2549
rect 16389 2546 16455 2549
rect 10869 2544 16455 2546
rect 10869 2488 10874 2544
rect 10930 2488 16394 2544
rect 16450 2488 16455 2544
rect 10869 2486 16455 2488
rect 10869 2483 10935 2486
rect 16389 2483 16455 2486
rect 0 2274 480 2304
rect 3693 2274 3759 2277
rect 0 2272 3759 2274
rect 0 2216 3698 2272
rect 3754 2216 3759 2272
rect 0 2214 3759 2216
rect 0 2184 480 2214
rect 3693 2211 3759 2214
rect 17493 2274 17559 2277
rect 19520 2274 20000 2304
rect 17493 2272 20000 2274
rect 17493 2216 17498 2272
rect 17554 2216 20000 2272
rect 17493 2214 20000 2216
rect 17493 2211 17559 2214
rect 3909 2208 4229 2209
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2143 4229 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 15770 2208 16090 2209
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 19520 2184 20000 2214
rect 15770 2143 16090 2144
rect 0 1866 480 1896
rect 2957 1866 3023 1869
rect 0 1864 3023 1866
rect 0 1808 2962 1864
rect 3018 1808 3023 1864
rect 0 1806 3023 1808
rect 0 1776 480 1806
rect 2957 1803 3023 1806
rect 17033 1866 17099 1869
rect 19520 1866 20000 1896
rect 17033 1864 20000 1866
rect 17033 1808 17038 1864
rect 17094 1808 20000 1864
rect 17033 1806 20000 1808
rect 17033 1803 17099 1806
rect 19520 1776 20000 1806
rect 0 1458 480 1488
rect 3417 1458 3483 1461
rect 0 1456 3483 1458
rect 0 1400 3422 1456
rect 3478 1400 3483 1456
rect 0 1398 3483 1400
rect 0 1368 480 1398
rect 3417 1395 3483 1398
rect 17585 1458 17651 1461
rect 19520 1458 20000 1488
rect 17585 1456 20000 1458
rect 17585 1400 17590 1456
rect 17646 1400 20000 1456
rect 17585 1398 20000 1400
rect 17585 1395 17651 1398
rect 19520 1368 20000 1398
rect 0 1050 480 1080
rect 3785 1050 3851 1053
rect 0 1048 3851 1050
rect 0 992 3790 1048
rect 3846 992 3851 1048
rect 0 990 3851 992
rect 0 960 480 990
rect 3785 987 3851 990
rect 17677 1050 17743 1053
rect 19520 1050 20000 1080
rect 17677 1048 20000 1050
rect 17677 992 17682 1048
rect 17738 992 20000 1048
rect 17677 990 20000 992
rect 17677 987 17743 990
rect 19520 960 20000 990
rect 0 642 480 672
rect 3325 642 3391 645
rect 0 640 3391 642
rect 0 584 3330 640
rect 3386 584 3391 640
rect 0 582 3391 584
rect 0 552 480 582
rect 3325 579 3391 582
rect 18045 642 18111 645
rect 19520 642 20000 672
rect 18045 640 20000 642
rect 18045 584 18050 640
rect 18106 584 20000 640
rect 18045 582 20000 584
rect 18045 579 18111 582
rect 19520 552 20000 582
rect 0 234 480 264
rect 2773 234 2839 237
rect 0 232 2839 234
rect 0 176 2778 232
rect 2834 176 2839 232
rect 0 174 2839 176
rect 0 144 480 174
rect 2773 171 2839 174
rect 18229 234 18295 237
rect 19520 234 20000 264
rect 18229 232 20000 234
rect 18229 176 18234 232
rect 18290 176 20000 232
rect 18229 174 20000 176
rect 18229 171 18295 174
rect 19520 144 20000 174
<< via3 >>
rect 4660 16220 4724 16284
rect 6882 14716 6946 14720
rect 6882 14660 6886 14716
rect 6886 14660 6942 14716
rect 6942 14660 6946 14716
rect 6882 14656 6946 14660
rect 6962 14716 7026 14720
rect 6962 14660 6966 14716
rect 6966 14660 7022 14716
rect 7022 14660 7026 14716
rect 6962 14656 7026 14660
rect 7042 14716 7106 14720
rect 7042 14660 7046 14716
rect 7046 14660 7102 14716
rect 7102 14660 7106 14716
rect 7042 14656 7106 14660
rect 7122 14716 7186 14720
rect 7122 14660 7126 14716
rect 7126 14660 7182 14716
rect 7182 14660 7186 14716
rect 7122 14656 7186 14660
rect 12813 14716 12877 14720
rect 12813 14660 12817 14716
rect 12817 14660 12873 14716
rect 12873 14660 12877 14716
rect 12813 14656 12877 14660
rect 12893 14716 12957 14720
rect 12893 14660 12897 14716
rect 12897 14660 12953 14716
rect 12953 14660 12957 14716
rect 12893 14656 12957 14660
rect 12973 14716 13037 14720
rect 12973 14660 12977 14716
rect 12977 14660 13033 14716
rect 13033 14660 13037 14716
rect 12973 14656 13037 14660
rect 13053 14716 13117 14720
rect 13053 14660 13057 14716
rect 13057 14660 13113 14716
rect 13113 14660 13117 14716
rect 13053 14656 13117 14660
rect 3917 14172 3981 14176
rect 3917 14116 3921 14172
rect 3921 14116 3977 14172
rect 3977 14116 3981 14172
rect 3917 14112 3981 14116
rect 3997 14172 4061 14176
rect 3997 14116 4001 14172
rect 4001 14116 4057 14172
rect 4057 14116 4061 14172
rect 3997 14112 4061 14116
rect 4077 14172 4141 14176
rect 4077 14116 4081 14172
rect 4081 14116 4137 14172
rect 4137 14116 4141 14172
rect 4077 14112 4141 14116
rect 4157 14172 4221 14176
rect 4157 14116 4161 14172
rect 4161 14116 4217 14172
rect 4217 14116 4221 14172
rect 4157 14112 4221 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 15778 14172 15842 14176
rect 15778 14116 15782 14172
rect 15782 14116 15838 14172
rect 15838 14116 15842 14172
rect 15778 14112 15842 14116
rect 15858 14172 15922 14176
rect 15858 14116 15862 14172
rect 15862 14116 15918 14172
rect 15918 14116 15922 14172
rect 15858 14112 15922 14116
rect 15938 14172 16002 14176
rect 15938 14116 15942 14172
rect 15942 14116 15998 14172
rect 15998 14116 16002 14172
rect 15938 14112 16002 14116
rect 16018 14172 16082 14176
rect 16018 14116 16022 14172
rect 16022 14116 16078 14172
rect 16078 14116 16082 14172
rect 16018 14112 16082 14116
rect 6882 13628 6946 13632
rect 6882 13572 6886 13628
rect 6886 13572 6942 13628
rect 6942 13572 6946 13628
rect 6882 13568 6946 13572
rect 6962 13628 7026 13632
rect 6962 13572 6966 13628
rect 6966 13572 7022 13628
rect 7022 13572 7026 13628
rect 6962 13568 7026 13572
rect 7042 13628 7106 13632
rect 7042 13572 7046 13628
rect 7046 13572 7102 13628
rect 7102 13572 7106 13628
rect 7042 13568 7106 13572
rect 7122 13628 7186 13632
rect 7122 13572 7126 13628
rect 7126 13572 7182 13628
rect 7182 13572 7186 13628
rect 7122 13568 7186 13572
rect 12813 13628 12877 13632
rect 12813 13572 12817 13628
rect 12817 13572 12873 13628
rect 12873 13572 12877 13628
rect 12813 13568 12877 13572
rect 12893 13628 12957 13632
rect 12893 13572 12897 13628
rect 12897 13572 12953 13628
rect 12953 13572 12957 13628
rect 12893 13568 12957 13572
rect 12973 13628 13037 13632
rect 12973 13572 12977 13628
rect 12977 13572 13033 13628
rect 13033 13572 13037 13628
rect 12973 13568 13037 13572
rect 13053 13628 13117 13632
rect 13053 13572 13057 13628
rect 13057 13572 13113 13628
rect 13113 13572 13117 13628
rect 13053 13568 13117 13572
rect 3917 13084 3981 13088
rect 3917 13028 3921 13084
rect 3921 13028 3977 13084
rect 3977 13028 3981 13084
rect 3917 13024 3981 13028
rect 3997 13084 4061 13088
rect 3997 13028 4001 13084
rect 4001 13028 4057 13084
rect 4057 13028 4061 13084
rect 3997 13024 4061 13028
rect 4077 13084 4141 13088
rect 4077 13028 4081 13084
rect 4081 13028 4137 13084
rect 4137 13028 4141 13084
rect 4077 13024 4141 13028
rect 4157 13084 4221 13088
rect 4157 13028 4161 13084
rect 4161 13028 4217 13084
rect 4217 13028 4221 13084
rect 4157 13024 4221 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 15778 13084 15842 13088
rect 15778 13028 15782 13084
rect 15782 13028 15838 13084
rect 15838 13028 15842 13084
rect 15778 13024 15842 13028
rect 15858 13084 15922 13088
rect 15858 13028 15862 13084
rect 15862 13028 15918 13084
rect 15918 13028 15922 13084
rect 15858 13024 15922 13028
rect 15938 13084 16002 13088
rect 15938 13028 15942 13084
rect 15942 13028 15998 13084
rect 15998 13028 16002 13084
rect 15938 13024 16002 13028
rect 16018 13084 16082 13088
rect 16018 13028 16022 13084
rect 16022 13028 16078 13084
rect 16078 13028 16082 13084
rect 16018 13024 16082 13028
rect 6882 12540 6946 12544
rect 6882 12484 6886 12540
rect 6886 12484 6942 12540
rect 6942 12484 6946 12540
rect 6882 12480 6946 12484
rect 6962 12540 7026 12544
rect 6962 12484 6966 12540
rect 6966 12484 7022 12540
rect 7022 12484 7026 12540
rect 6962 12480 7026 12484
rect 7042 12540 7106 12544
rect 7042 12484 7046 12540
rect 7046 12484 7102 12540
rect 7102 12484 7106 12540
rect 7042 12480 7106 12484
rect 7122 12540 7186 12544
rect 7122 12484 7126 12540
rect 7126 12484 7182 12540
rect 7182 12484 7186 12540
rect 7122 12480 7186 12484
rect 12813 12540 12877 12544
rect 12813 12484 12817 12540
rect 12817 12484 12873 12540
rect 12873 12484 12877 12540
rect 12813 12480 12877 12484
rect 12893 12540 12957 12544
rect 12893 12484 12897 12540
rect 12897 12484 12953 12540
rect 12953 12484 12957 12540
rect 12893 12480 12957 12484
rect 12973 12540 13037 12544
rect 12973 12484 12977 12540
rect 12977 12484 13033 12540
rect 13033 12484 13037 12540
rect 12973 12480 13037 12484
rect 13053 12540 13117 12544
rect 13053 12484 13057 12540
rect 13057 12484 13113 12540
rect 13113 12484 13117 12540
rect 13053 12480 13117 12484
rect 3917 11996 3981 12000
rect 3917 11940 3921 11996
rect 3921 11940 3977 11996
rect 3977 11940 3981 11996
rect 3917 11936 3981 11940
rect 3997 11996 4061 12000
rect 3997 11940 4001 11996
rect 4001 11940 4057 11996
rect 4057 11940 4061 11996
rect 3997 11936 4061 11940
rect 4077 11996 4141 12000
rect 4077 11940 4081 11996
rect 4081 11940 4137 11996
rect 4137 11940 4141 11996
rect 4077 11936 4141 11940
rect 4157 11996 4221 12000
rect 4157 11940 4161 11996
rect 4161 11940 4217 11996
rect 4217 11940 4221 11996
rect 4157 11936 4221 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 15778 11996 15842 12000
rect 15778 11940 15782 11996
rect 15782 11940 15838 11996
rect 15838 11940 15842 11996
rect 15778 11936 15842 11940
rect 15858 11996 15922 12000
rect 15858 11940 15862 11996
rect 15862 11940 15918 11996
rect 15918 11940 15922 11996
rect 15858 11936 15922 11940
rect 15938 11996 16002 12000
rect 15938 11940 15942 11996
rect 15942 11940 15998 11996
rect 15998 11940 16002 11996
rect 15938 11936 16002 11940
rect 16018 11996 16082 12000
rect 16018 11940 16022 11996
rect 16022 11940 16078 11996
rect 16078 11940 16082 11996
rect 16018 11936 16082 11940
rect 6882 11452 6946 11456
rect 6882 11396 6886 11452
rect 6886 11396 6942 11452
rect 6942 11396 6946 11452
rect 6882 11392 6946 11396
rect 6962 11452 7026 11456
rect 6962 11396 6966 11452
rect 6966 11396 7022 11452
rect 7022 11396 7026 11452
rect 6962 11392 7026 11396
rect 7042 11452 7106 11456
rect 7042 11396 7046 11452
rect 7046 11396 7102 11452
rect 7102 11396 7106 11452
rect 7042 11392 7106 11396
rect 7122 11452 7186 11456
rect 7122 11396 7126 11452
rect 7126 11396 7182 11452
rect 7182 11396 7186 11452
rect 7122 11392 7186 11396
rect 12813 11452 12877 11456
rect 12813 11396 12817 11452
rect 12817 11396 12873 11452
rect 12873 11396 12877 11452
rect 12813 11392 12877 11396
rect 12893 11452 12957 11456
rect 12893 11396 12897 11452
rect 12897 11396 12953 11452
rect 12953 11396 12957 11452
rect 12893 11392 12957 11396
rect 12973 11452 13037 11456
rect 12973 11396 12977 11452
rect 12977 11396 13033 11452
rect 13033 11396 13037 11452
rect 12973 11392 13037 11396
rect 13053 11452 13117 11456
rect 13053 11396 13057 11452
rect 13057 11396 13113 11452
rect 13113 11396 13117 11452
rect 13053 11392 13117 11396
rect 9628 11188 9692 11252
rect 3917 10908 3981 10912
rect 3917 10852 3921 10908
rect 3921 10852 3977 10908
rect 3977 10852 3981 10908
rect 3917 10848 3981 10852
rect 3997 10908 4061 10912
rect 3997 10852 4001 10908
rect 4001 10852 4057 10908
rect 4057 10852 4061 10908
rect 3997 10848 4061 10852
rect 4077 10908 4141 10912
rect 4077 10852 4081 10908
rect 4081 10852 4137 10908
rect 4137 10852 4141 10908
rect 4077 10848 4141 10852
rect 4157 10908 4221 10912
rect 4157 10852 4161 10908
rect 4161 10852 4217 10908
rect 4217 10852 4221 10908
rect 4157 10848 4221 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 15778 10908 15842 10912
rect 15778 10852 15782 10908
rect 15782 10852 15838 10908
rect 15838 10852 15842 10908
rect 15778 10848 15842 10852
rect 15858 10908 15922 10912
rect 15858 10852 15862 10908
rect 15862 10852 15918 10908
rect 15918 10852 15922 10908
rect 15858 10848 15922 10852
rect 15938 10908 16002 10912
rect 15938 10852 15942 10908
rect 15942 10852 15998 10908
rect 15998 10852 16002 10908
rect 15938 10848 16002 10852
rect 16018 10908 16082 10912
rect 16018 10852 16022 10908
rect 16022 10852 16078 10908
rect 16078 10852 16082 10908
rect 16018 10848 16082 10852
rect 9628 10508 9692 10572
rect 6882 10364 6946 10368
rect 6882 10308 6886 10364
rect 6886 10308 6942 10364
rect 6942 10308 6946 10364
rect 6882 10304 6946 10308
rect 6962 10364 7026 10368
rect 6962 10308 6966 10364
rect 6966 10308 7022 10364
rect 7022 10308 7026 10364
rect 6962 10304 7026 10308
rect 7042 10364 7106 10368
rect 7042 10308 7046 10364
rect 7046 10308 7102 10364
rect 7102 10308 7106 10364
rect 7042 10304 7106 10308
rect 7122 10364 7186 10368
rect 7122 10308 7126 10364
rect 7126 10308 7182 10364
rect 7182 10308 7186 10364
rect 7122 10304 7186 10308
rect 12813 10364 12877 10368
rect 12813 10308 12817 10364
rect 12817 10308 12873 10364
rect 12873 10308 12877 10364
rect 12813 10304 12877 10308
rect 12893 10364 12957 10368
rect 12893 10308 12897 10364
rect 12897 10308 12953 10364
rect 12953 10308 12957 10364
rect 12893 10304 12957 10308
rect 12973 10364 13037 10368
rect 12973 10308 12977 10364
rect 12977 10308 13033 10364
rect 13033 10308 13037 10364
rect 12973 10304 13037 10308
rect 13053 10364 13117 10368
rect 13053 10308 13057 10364
rect 13057 10308 13113 10364
rect 13113 10308 13117 10364
rect 13053 10304 13117 10308
rect 3917 9820 3981 9824
rect 3917 9764 3921 9820
rect 3921 9764 3977 9820
rect 3977 9764 3981 9820
rect 3917 9760 3981 9764
rect 3997 9820 4061 9824
rect 3997 9764 4001 9820
rect 4001 9764 4057 9820
rect 4057 9764 4061 9820
rect 3997 9760 4061 9764
rect 4077 9820 4141 9824
rect 4077 9764 4081 9820
rect 4081 9764 4137 9820
rect 4137 9764 4141 9820
rect 4077 9760 4141 9764
rect 4157 9820 4221 9824
rect 4157 9764 4161 9820
rect 4161 9764 4217 9820
rect 4217 9764 4221 9820
rect 4157 9760 4221 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 15778 9820 15842 9824
rect 15778 9764 15782 9820
rect 15782 9764 15838 9820
rect 15838 9764 15842 9820
rect 15778 9760 15842 9764
rect 15858 9820 15922 9824
rect 15858 9764 15862 9820
rect 15862 9764 15918 9820
rect 15918 9764 15922 9820
rect 15858 9760 15922 9764
rect 15938 9820 16002 9824
rect 15938 9764 15942 9820
rect 15942 9764 15998 9820
rect 15998 9764 16002 9820
rect 15938 9760 16002 9764
rect 16018 9820 16082 9824
rect 16018 9764 16022 9820
rect 16022 9764 16078 9820
rect 16078 9764 16082 9820
rect 16018 9760 16082 9764
rect 4660 9692 4724 9756
rect 6684 9420 6748 9484
rect 6882 9276 6946 9280
rect 6882 9220 6886 9276
rect 6886 9220 6942 9276
rect 6942 9220 6946 9276
rect 6882 9216 6946 9220
rect 6962 9276 7026 9280
rect 6962 9220 6966 9276
rect 6966 9220 7022 9276
rect 7022 9220 7026 9276
rect 6962 9216 7026 9220
rect 7042 9276 7106 9280
rect 7042 9220 7046 9276
rect 7046 9220 7102 9276
rect 7102 9220 7106 9276
rect 7042 9216 7106 9220
rect 7122 9276 7186 9280
rect 7122 9220 7126 9276
rect 7126 9220 7182 9276
rect 7182 9220 7186 9276
rect 7122 9216 7186 9220
rect 4292 9012 4356 9076
rect 12813 9276 12877 9280
rect 12813 9220 12817 9276
rect 12817 9220 12873 9276
rect 12873 9220 12877 9276
rect 12813 9216 12877 9220
rect 12893 9276 12957 9280
rect 12893 9220 12897 9276
rect 12897 9220 12953 9276
rect 12953 9220 12957 9276
rect 12893 9216 12957 9220
rect 12973 9276 13037 9280
rect 12973 9220 12977 9276
rect 12977 9220 13033 9276
rect 13033 9220 13037 9276
rect 12973 9216 13037 9220
rect 13053 9276 13117 9280
rect 13053 9220 13057 9276
rect 13057 9220 13113 9276
rect 13113 9220 13117 9276
rect 13053 9216 13117 9220
rect 3917 8732 3981 8736
rect 3917 8676 3921 8732
rect 3921 8676 3977 8732
rect 3977 8676 3981 8732
rect 3917 8672 3981 8676
rect 3997 8732 4061 8736
rect 3997 8676 4001 8732
rect 4001 8676 4057 8732
rect 4057 8676 4061 8732
rect 3997 8672 4061 8676
rect 4077 8732 4141 8736
rect 4077 8676 4081 8732
rect 4081 8676 4137 8732
rect 4137 8676 4141 8732
rect 4077 8672 4141 8676
rect 4157 8732 4221 8736
rect 4157 8676 4161 8732
rect 4161 8676 4217 8732
rect 4217 8676 4221 8732
rect 4157 8672 4221 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 15778 8732 15842 8736
rect 15778 8676 15782 8732
rect 15782 8676 15838 8732
rect 15838 8676 15842 8732
rect 15778 8672 15842 8676
rect 15858 8732 15922 8736
rect 15858 8676 15862 8732
rect 15862 8676 15918 8732
rect 15918 8676 15922 8732
rect 15858 8672 15922 8676
rect 15938 8732 16002 8736
rect 15938 8676 15942 8732
rect 15942 8676 15998 8732
rect 15998 8676 16002 8732
rect 15938 8672 16002 8676
rect 16018 8732 16082 8736
rect 16018 8676 16022 8732
rect 16022 8676 16078 8732
rect 16078 8676 16082 8732
rect 16018 8672 16082 8676
rect 6882 8188 6946 8192
rect 6882 8132 6886 8188
rect 6886 8132 6942 8188
rect 6942 8132 6946 8188
rect 6882 8128 6946 8132
rect 6962 8188 7026 8192
rect 6962 8132 6966 8188
rect 6966 8132 7022 8188
rect 7022 8132 7026 8188
rect 6962 8128 7026 8132
rect 7042 8188 7106 8192
rect 7042 8132 7046 8188
rect 7046 8132 7102 8188
rect 7102 8132 7106 8188
rect 7042 8128 7106 8132
rect 7122 8188 7186 8192
rect 7122 8132 7126 8188
rect 7126 8132 7182 8188
rect 7182 8132 7186 8188
rect 7122 8128 7186 8132
rect 12813 8188 12877 8192
rect 12813 8132 12817 8188
rect 12817 8132 12873 8188
rect 12873 8132 12877 8188
rect 12813 8128 12877 8132
rect 12893 8188 12957 8192
rect 12893 8132 12897 8188
rect 12897 8132 12953 8188
rect 12953 8132 12957 8188
rect 12893 8128 12957 8132
rect 12973 8188 13037 8192
rect 12973 8132 12977 8188
rect 12977 8132 13033 8188
rect 13033 8132 13037 8188
rect 12973 8128 13037 8132
rect 13053 8188 13117 8192
rect 13053 8132 13057 8188
rect 13057 8132 13113 8188
rect 13113 8132 13117 8188
rect 13053 8128 13117 8132
rect 3917 7644 3981 7648
rect 3917 7588 3921 7644
rect 3921 7588 3977 7644
rect 3977 7588 3981 7644
rect 3917 7584 3981 7588
rect 3997 7644 4061 7648
rect 3997 7588 4001 7644
rect 4001 7588 4057 7644
rect 4057 7588 4061 7644
rect 3997 7584 4061 7588
rect 4077 7644 4141 7648
rect 4077 7588 4081 7644
rect 4081 7588 4137 7644
rect 4137 7588 4141 7644
rect 4077 7584 4141 7588
rect 4157 7644 4221 7648
rect 4157 7588 4161 7644
rect 4161 7588 4217 7644
rect 4217 7588 4221 7644
rect 4157 7584 4221 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 15778 7644 15842 7648
rect 15778 7588 15782 7644
rect 15782 7588 15838 7644
rect 15838 7588 15842 7644
rect 15778 7584 15842 7588
rect 15858 7644 15922 7648
rect 15858 7588 15862 7644
rect 15862 7588 15918 7644
rect 15918 7588 15922 7644
rect 15858 7584 15922 7588
rect 15938 7644 16002 7648
rect 15938 7588 15942 7644
rect 15942 7588 15998 7644
rect 15998 7588 16002 7644
rect 15938 7584 16002 7588
rect 16018 7644 16082 7648
rect 16018 7588 16022 7644
rect 16022 7588 16078 7644
rect 16078 7588 16082 7644
rect 16018 7584 16082 7588
rect 6684 7244 6748 7308
rect 6882 7100 6946 7104
rect 6882 7044 6886 7100
rect 6886 7044 6942 7100
rect 6942 7044 6946 7100
rect 6882 7040 6946 7044
rect 6962 7100 7026 7104
rect 6962 7044 6966 7100
rect 6966 7044 7022 7100
rect 7022 7044 7026 7100
rect 6962 7040 7026 7044
rect 7042 7100 7106 7104
rect 7042 7044 7046 7100
rect 7046 7044 7102 7100
rect 7102 7044 7106 7100
rect 7042 7040 7106 7044
rect 7122 7100 7186 7104
rect 7122 7044 7126 7100
rect 7126 7044 7182 7100
rect 7182 7044 7186 7100
rect 7122 7040 7186 7044
rect 12813 7100 12877 7104
rect 12813 7044 12817 7100
rect 12817 7044 12873 7100
rect 12873 7044 12877 7100
rect 12813 7040 12877 7044
rect 12893 7100 12957 7104
rect 12893 7044 12897 7100
rect 12897 7044 12953 7100
rect 12953 7044 12957 7100
rect 12893 7040 12957 7044
rect 12973 7100 13037 7104
rect 12973 7044 12977 7100
rect 12977 7044 13033 7100
rect 13033 7044 13037 7100
rect 12973 7040 13037 7044
rect 13053 7100 13117 7104
rect 13053 7044 13057 7100
rect 13057 7044 13113 7100
rect 13113 7044 13117 7100
rect 13053 7040 13117 7044
rect 3917 6556 3981 6560
rect 3917 6500 3921 6556
rect 3921 6500 3977 6556
rect 3977 6500 3981 6556
rect 3917 6496 3981 6500
rect 3997 6556 4061 6560
rect 3997 6500 4001 6556
rect 4001 6500 4057 6556
rect 4057 6500 4061 6556
rect 3997 6496 4061 6500
rect 4077 6556 4141 6560
rect 4077 6500 4081 6556
rect 4081 6500 4137 6556
rect 4137 6500 4141 6556
rect 4077 6496 4141 6500
rect 4157 6556 4221 6560
rect 4157 6500 4161 6556
rect 4161 6500 4217 6556
rect 4217 6500 4221 6556
rect 4157 6496 4221 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 15778 6556 15842 6560
rect 15778 6500 15782 6556
rect 15782 6500 15838 6556
rect 15838 6500 15842 6556
rect 15778 6496 15842 6500
rect 15858 6556 15922 6560
rect 15858 6500 15862 6556
rect 15862 6500 15918 6556
rect 15918 6500 15922 6556
rect 15858 6496 15922 6500
rect 15938 6556 16002 6560
rect 15938 6500 15942 6556
rect 15942 6500 15998 6556
rect 15998 6500 16002 6556
rect 15938 6496 16002 6500
rect 16018 6556 16082 6560
rect 16018 6500 16022 6556
rect 16022 6500 16078 6556
rect 16078 6500 16082 6556
rect 16018 6496 16082 6500
rect 6882 6012 6946 6016
rect 6882 5956 6886 6012
rect 6886 5956 6942 6012
rect 6942 5956 6946 6012
rect 6882 5952 6946 5956
rect 6962 6012 7026 6016
rect 6962 5956 6966 6012
rect 6966 5956 7022 6012
rect 7022 5956 7026 6012
rect 6962 5952 7026 5956
rect 7042 6012 7106 6016
rect 7042 5956 7046 6012
rect 7046 5956 7102 6012
rect 7102 5956 7106 6012
rect 7042 5952 7106 5956
rect 7122 6012 7186 6016
rect 7122 5956 7126 6012
rect 7126 5956 7182 6012
rect 7182 5956 7186 6012
rect 7122 5952 7186 5956
rect 12813 6012 12877 6016
rect 12813 5956 12817 6012
rect 12817 5956 12873 6012
rect 12873 5956 12877 6012
rect 12813 5952 12877 5956
rect 12893 6012 12957 6016
rect 12893 5956 12897 6012
rect 12897 5956 12953 6012
rect 12953 5956 12957 6012
rect 12893 5952 12957 5956
rect 12973 6012 13037 6016
rect 12973 5956 12977 6012
rect 12977 5956 13033 6012
rect 13033 5956 13037 6012
rect 12973 5952 13037 5956
rect 13053 6012 13117 6016
rect 13053 5956 13057 6012
rect 13057 5956 13113 6012
rect 13113 5956 13117 6012
rect 13053 5952 13117 5956
rect 3917 5468 3981 5472
rect 3917 5412 3921 5468
rect 3921 5412 3977 5468
rect 3977 5412 3981 5468
rect 3917 5408 3981 5412
rect 3997 5468 4061 5472
rect 3997 5412 4001 5468
rect 4001 5412 4057 5468
rect 4057 5412 4061 5468
rect 3997 5408 4061 5412
rect 4077 5468 4141 5472
rect 4077 5412 4081 5468
rect 4081 5412 4137 5468
rect 4137 5412 4141 5468
rect 4077 5408 4141 5412
rect 4157 5468 4221 5472
rect 4157 5412 4161 5468
rect 4161 5412 4217 5468
rect 4217 5412 4221 5468
rect 4157 5408 4221 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 15778 5468 15842 5472
rect 15778 5412 15782 5468
rect 15782 5412 15838 5468
rect 15838 5412 15842 5468
rect 15778 5408 15842 5412
rect 15858 5468 15922 5472
rect 15858 5412 15862 5468
rect 15862 5412 15918 5468
rect 15918 5412 15922 5468
rect 15858 5408 15922 5412
rect 15938 5468 16002 5472
rect 15938 5412 15942 5468
rect 15942 5412 15998 5468
rect 15998 5412 16002 5468
rect 15938 5408 16002 5412
rect 16018 5468 16082 5472
rect 16018 5412 16022 5468
rect 16022 5412 16078 5468
rect 16078 5412 16082 5468
rect 16018 5408 16082 5412
rect 4292 4992 4356 4996
rect 4292 4936 4342 4992
rect 4342 4936 4356 4992
rect 4292 4932 4356 4936
rect 6882 4924 6946 4928
rect 6882 4868 6886 4924
rect 6886 4868 6942 4924
rect 6942 4868 6946 4924
rect 6882 4864 6946 4868
rect 6962 4924 7026 4928
rect 6962 4868 6966 4924
rect 6966 4868 7022 4924
rect 7022 4868 7026 4924
rect 6962 4864 7026 4868
rect 7042 4924 7106 4928
rect 7042 4868 7046 4924
rect 7046 4868 7102 4924
rect 7102 4868 7106 4924
rect 7042 4864 7106 4868
rect 7122 4924 7186 4928
rect 7122 4868 7126 4924
rect 7126 4868 7182 4924
rect 7182 4868 7186 4924
rect 7122 4864 7186 4868
rect 12813 4924 12877 4928
rect 12813 4868 12817 4924
rect 12817 4868 12873 4924
rect 12873 4868 12877 4924
rect 12813 4864 12877 4868
rect 12893 4924 12957 4928
rect 12893 4868 12897 4924
rect 12897 4868 12953 4924
rect 12953 4868 12957 4924
rect 12893 4864 12957 4868
rect 12973 4924 13037 4928
rect 12973 4868 12977 4924
rect 12977 4868 13033 4924
rect 13033 4868 13037 4924
rect 12973 4864 13037 4868
rect 13053 4924 13117 4928
rect 13053 4868 13057 4924
rect 13057 4868 13113 4924
rect 13113 4868 13117 4924
rect 13053 4864 13117 4868
rect 3917 4380 3981 4384
rect 3917 4324 3921 4380
rect 3921 4324 3977 4380
rect 3977 4324 3981 4380
rect 3917 4320 3981 4324
rect 3997 4380 4061 4384
rect 3997 4324 4001 4380
rect 4001 4324 4057 4380
rect 4057 4324 4061 4380
rect 3997 4320 4061 4324
rect 4077 4380 4141 4384
rect 4077 4324 4081 4380
rect 4081 4324 4137 4380
rect 4137 4324 4141 4380
rect 4077 4320 4141 4324
rect 4157 4380 4221 4384
rect 4157 4324 4161 4380
rect 4161 4324 4217 4380
rect 4217 4324 4221 4380
rect 4157 4320 4221 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 15778 4380 15842 4384
rect 15778 4324 15782 4380
rect 15782 4324 15838 4380
rect 15838 4324 15842 4380
rect 15778 4320 15842 4324
rect 15858 4380 15922 4384
rect 15858 4324 15862 4380
rect 15862 4324 15918 4380
rect 15918 4324 15922 4380
rect 15858 4320 15922 4324
rect 15938 4380 16002 4384
rect 15938 4324 15942 4380
rect 15942 4324 15998 4380
rect 15998 4324 16002 4380
rect 15938 4320 16002 4324
rect 16018 4380 16082 4384
rect 16018 4324 16022 4380
rect 16022 4324 16078 4380
rect 16078 4324 16082 4380
rect 16018 4320 16082 4324
rect 6882 3836 6946 3840
rect 6882 3780 6886 3836
rect 6886 3780 6942 3836
rect 6942 3780 6946 3836
rect 6882 3776 6946 3780
rect 6962 3836 7026 3840
rect 6962 3780 6966 3836
rect 6966 3780 7022 3836
rect 7022 3780 7026 3836
rect 6962 3776 7026 3780
rect 7042 3836 7106 3840
rect 7042 3780 7046 3836
rect 7046 3780 7102 3836
rect 7102 3780 7106 3836
rect 7042 3776 7106 3780
rect 7122 3836 7186 3840
rect 7122 3780 7126 3836
rect 7126 3780 7182 3836
rect 7182 3780 7186 3836
rect 7122 3776 7186 3780
rect 12813 3836 12877 3840
rect 12813 3780 12817 3836
rect 12817 3780 12873 3836
rect 12873 3780 12877 3836
rect 12813 3776 12877 3780
rect 12893 3836 12957 3840
rect 12893 3780 12897 3836
rect 12897 3780 12953 3836
rect 12953 3780 12957 3836
rect 12893 3776 12957 3780
rect 12973 3836 13037 3840
rect 12973 3780 12977 3836
rect 12977 3780 13033 3836
rect 13033 3780 13037 3836
rect 12973 3776 13037 3780
rect 13053 3836 13117 3840
rect 13053 3780 13057 3836
rect 13057 3780 13113 3836
rect 13113 3780 13117 3836
rect 13053 3776 13117 3780
rect 3917 3292 3981 3296
rect 3917 3236 3921 3292
rect 3921 3236 3977 3292
rect 3977 3236 3981 3292
rect 3917 3232 3981 3236
rect 3997 3292 4061 3296
rect 3997 3236 4001 3292
rect 4001 3236 4057 3292
rect 4057 3236 4061 3292
rect 3997 3232 4061 3236
rect 4077 3292 4141 3296
rect 4077 3236 4081 3292
rect 4081 3236 4137 3292
rect 4137 3236 4141 3292
rect 4077 3232 4141 3236
rect 4157 3292 4221 3296
rect 4157 3236 4161 3292
rect 4161 3236 4217 3292
rect 4217 3236 4221 3292
rect 4157 3232 4221 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 15778 3292 15842 3296
rect 15778 3236 15782 3292
rect 15782 3236 15838 3292
rect 15838 3236 15842 3292
rect 15778 3232 15842 3236
rect 15858 3292 15922 3296
rect 15858 3236 15862 3292
rect 15862 3236 15918 3292
rect 15918 3236 15922 3292
rect 15858 3232 15922 3236
rect 15938 3292 16002 3296
rect 15938 3236 15942 3292
rect 15942 3236 15998 3292
rect 15998 3236 16002 3292
rect 15938 3232 16002 3236
rect 16018 3292 16082 3296
rect 16018 3236 16022 3292
rect 16022 3236 16078 3292
rect 16078 3236 16082 3292
rect 16018 3232 16082 3236
rect 6882 2748 6946 2752
rect 6882 2692 6886 2748
rect 6886 2692 6942 2748
rect 6942 2692 6946 2748
rect 6882 2688 6946 2692
rect 6962 2748 7026 2752
rect 6962 2692 6966 2748
rect 6966 2692 7022 2748
rect 7022 2692 7026 2748
rect 6962 2688 7026 2692
rect 7042 2748 7106 2752
rect 7042 2692 7046 2748
rect 7046 2692 7102 2748
rect 7102 2692 7106 2748
rect 7042 2688 7106 2692
rect 7122 2748 7186 2752
rect 7122 2692 7126 2748
rect 7126 2692 7182 2748
rect 7182 2692 7186 2748
rect 7122 2688 7186 2692
rect 12813 2748 12877 2752
rect 12813 2692 12817 2748
rect 12817 2692 12873 2748
rect 12873 2692 12877 2748
rect 12813 2688 12877 2692
rect 12893 2748 12957 2752
rect 12893 2692 12897 2748
rect 12897 2692 12953 2748
rect 12953 2692 12957 2748
rect 12893 2688 12957 2692
rect 12973 2748 13037 2752
rect 12973 2692 12977 2748
rect 12977 2692 13033 2748
rect 13033 2692 13037 2748
rect 12973 2688 13037 2692
rect 13053 2748 13117 2752
rect 13053 2692 13057 2748
rect 13057 2692 13113 2748
rect 13113 2692 13117 2748
rect 13053 2688 13117 2692
rect 3917 2204 3981 2208
rect 3917 2148 3921 2204
rect 3921 2148 3977 2204
rect 3977 2148 3981 2204
rect 3917 2144 3981 2148
rect 3997 2204 4061 2208
rect 3997 2148 4001 2204
rect 4001 2148 4057 2204
rect 4057 2148 4061 2204
rect 3997 2144 4061 2148
rect 4077 2204 4141 2208
rect 4077 2148 4081 2204
rect 4081 2148 4137 2204
rect 4137 2148 4141 2204
rect 4077 2144 4141 2148
rect 4157 2204 4221 2208
rect 4157 2148 4161 2204
rect 4161 2148 4217 2204
rect 4217 2148 4221 2204
rect 4157 2144 4221 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 15778 2204 15842 2208
rect 15778 2148 15782 2204
rect 15782 2148 15838 2204
rect 15838 2148 15842 2204
rect 15778 2144 15842 2148
rect 15858 2204 15922 2208
rect 15858 2148 15862 2204
rect 15862 2148 15918 2204
rect 15918 2148 15922 2204
rect 15858 2144 15922 2148
rect 15938 2204 16002 2208
rect 15938 2148 15942 2204
rect 15942 2148 15998 2204
rect 15998 2148 16002 2204
rect 15938 2144 16002 2148
rect 16018 2204 16082 2208
rect 16018 2148 16022 2204
rect 16022 2148 16078 2204
rect 16078 2148 16082 2204
rect 16018 2144 16082 2148
<< metal4 >>
rect 4659 16284 4725 16285
rect 4659 16220 4660 16284
rect 4724 16220 4725 16284
rect 4659 16219 4725 16220
rect 3909 14176 4229 14736
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 13088 4229 14112
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 12000 4229 13024
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 10912 4229 11936
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 9824 4229 10848
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 8736 4229 9760
rect 4662 9757 4722 16219
rect 6874 14720 7195 14736
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7195 14720
rect 6874 13632 7195 14656
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7195 13632
rect 6874 12544 7195 13568
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7195 12544
rect 6874 11456 7195 12480
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7195 11456
rect 6874 10368 7195 11392
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9627 11252 9693 11253
rect 9627 11188 9628 11252
rect 9692 11188 9693 11252
rect 9627 11187 9693 11188
rect 9630 10573 9690 11187
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9627 10572 9693 10573
rect 9627 10508 9628 10572
rect 9692 10508 9693 10572
rect 9627 10507 9693 10508
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7195 10368
rect 4659 9756 4725 9757
rect 4659 9692 4660 9756
rect 4724 9692 4725 9756
rect 4659 9691 4725 9692
rect 6683 9484 6749 9485
rect 6683 9420 6684 9484
rect 6748 9420 6749 9484
rect 6683 9419 6749 9420
rect 4291 9076 4357 9077
rect 4291 9012 4292 9076
rect 4356 9012 4357 9076
rect 4291 9011 4357 9012
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 7648 4229 8672
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 6560 4229 7584
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 5472 4229 6496
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 4384 4229 5408
rect 4294 4997 4354 9011
rect 6686 7309 6746 9419
rect 6874 9280 7195 10304
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7195 9280
rect 6874 8192 7195 9216
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7195 8192
rect 6683 7308 6749 7309
rect 6683 7244 6684 7308
rect 6748 7244 6749 7308
rect 6683 7243 6749 7244
rect 6874 7104 7195 8128
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7195 7104
rect 6874 6016 7195 7040
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7195 6016
rect 4291 4996 4357 4997
rect 4291 4932 4292 4996
rect 4356 4932 4357 4996
rect 4291 4931 4357 4932
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 3296 4229 4320
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 2208 4229 3232
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2128 4229 2144
rect 6874 4928 7195 5952
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7195 4928
rect 6874 3840 7195 4864
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7195 3840
rect 6874 2752 7195 3776
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7195 2752
rect 6874 2128 7195 2688
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12805 14720 13125 14736
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 13632 13125 14656
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 12544 13125 13568
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 11456 13125 12480
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 10368 13125 11392
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 12805 9280 13125 10304
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 8192 13125 9216
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 7104 13125 8128
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 6016 13125 7040
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 4928 13125 5952
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 3840 13125 4864
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 2752 13125 3776
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2128 13125 2688
rect 15770 14176 16090 14736
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 15770 13088 16090 14112
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 12000 16090 13024
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 10912 16090 11936
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 9824 16090 10848
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15770 8736 16090 9760
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15770 7648 16090 8672
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 6560 16090 7584
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 5472 16090 6496
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 4384 16090 5408
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 15770 3296 16090 4320
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 2208 16090 3232
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 15770 2128 16090 2144
use sky130_fd_sc_hd__fill_2  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606256979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1606256979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1564 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _49_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1656 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_19
timestamp 1606256979
transform 1 0 2852 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_11
timestamp 1606256979
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18
timestamp 1606256979
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10
timestamp 1606256979
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2208 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2300 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 3128 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1606256979
transform 1 0 4416 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4508 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1606256979
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_31 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_46
timestamp 1606256979
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45
timestamp 1606256979
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 5428 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1606256979
transform 1 0 5520 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1606256979
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59
timestamp 1606256979
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53
timestamp 1606256979
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1606256979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1606256979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1606256979
transform 1 0 6164 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8096 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 7728 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1606256979
transform 1 0 8648 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69
timestamp 1606256979
transform 1 0 7452 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_78
timestamp 1606256979
transform 1 0 8280 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_74
timestamp 1606256979
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1606256979
transform 1 0 9108 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10120 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10212 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1606256979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1606256979
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1606256979
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 10120 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_85
timestamp 1606256979
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_96
timestamp 1606256979
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_107
timestamp 1606256979
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_108
timestamp 1606256979
transform 1 0 11040 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1606256979
transform 1 0 11224 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1606256979
transform 1 0 11132 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1606256979
transform 1 0 11960 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123
timestamp 1606256979
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119
timestamp 1606256979
transform 1 0 12052 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1606256979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1606256979
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1606256979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14076 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13340 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13984 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131
timestamp 1606256979
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_139
timestamp 1606256979
transform 1 0 13892 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_132 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 13248 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1606256979
transform 1 0 16192 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15456 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14720 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1606256979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_147
timestamp 1606256979
transform 1 0 14628 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_146
timestamp 1606256979
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1606256979
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_162
timestamp 1606256979
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_175
timestamp 1606256979
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_168
timestamp 1606256979
transform 1 0 16560 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_168
timestamp 1606256979
transform 1 0 16560 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606256979
transform 1 0 16836 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1606256979
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1606256979
transform 1 0 17756 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_176
timestamp 1606256979
transform 1 0 17296 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1606256979
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1606256979
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606256979
transform 1 0 17388 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606256979
transform 1 0 17388 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1606256979
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1606256979
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1606256979
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1606256979
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1606256979
transform 1 0 2300 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1564 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1606256979
transform 1 0 2944 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1606256979
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1606256979
transform 1 0 2116 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_17
timestamp 1606256979
transform 1 0 2668 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4416 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1606256979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1606256979
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1606256979
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5428 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_45
timestamp 1606256979
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7084 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 8740 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_63
timestamp 1606256979
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_81
timestamp 1606256979
transform 1 0 8556 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10672 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1606256979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1606256979
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_102
timestamp 1606256979
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1606256979
transform 1 0 11684 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12236 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_113
timestamp 1606256979
transform 1 0 11500 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_119
timestamp 1606256979
transform 1 0 12052 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13892 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_137
timestamp 1606256979
transform 1 0 13708 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1606256979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1606256979
transform 1 0 14720 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1606256979
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_160
timestamp 1606256979
transform 1 0 15824 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606256979
transform 1 0 17296 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1606256979
transform 1 0 17848 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1606256979
transform 1 0 16928 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_180
timestamp 1606256979
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_186
timestamp 1606256979
transform 1 0 18216 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 2668 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1606256979
transform 1 0 1656 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1606256979
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1606256979
transform 1 0 4324 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_33
timestamp 1606256979
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_39
timestamp 1606256979
transform 1 0 4692 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1606256979
transform 1 0 4968 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 5980 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 6808 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1606256979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_51
timestamp 1606256979
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606256979
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1606256979
transform 1 0 7636 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8648 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_3_68
timestamp 1606256979
transform 1 0 7360 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_80
timestamp 1606256979
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 10672 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1606256979
transform 1 0 9660 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_91
timestamp 1606256979
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_102
timestamp 1606256979
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1606256979
transform 1 0 12512 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1606256979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1606256979
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1606256979
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13616 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_3_133
timestamp 1606256979
transform 1 0 13340 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_152
timestamp 1606256979
transform 1 0 15088 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_164
timestamp 1606256979
transform 1 0 16192 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606256979
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606256979
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1606256979
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_176
timestamp 1606256979
transform 1 0 17296 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1606256979
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_188
timestamp 1606256979
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1606256979
transform 1 0 1472 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2024 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1606256979
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_8
timestamp 1606256979
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4048 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1606256979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_26
timestamp 1606256979
transform 1 0 3496 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1606256979
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1606256979
transform 1 0 6716 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1606256979
transform 1 0 5704 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_48
timestamp 1606256979
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1606256979
transform 1 0 6532 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7820 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_4_70
timestamp 1606256979
transform 1 0 7544 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 9752 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1606256979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1606256979
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1606256979
transform 1 0 9660 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1606256979
transform 1 0 11408 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_110
timestamp 1606256979
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_121
timestamp 1606256979
transform 1 0 12236 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_125
timestamp 1606256979
transform 1 0 12604 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13708 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1606256979
transform 1 0 12696 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_135
timestamp 1606256979
transform 1 0 13524 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1606256979
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1606256979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_146
timestamp 1606256979
transform 1 0 14536 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1606256979
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_163
timestamp 1606256979
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606256979
transform 1 0 17296 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1606256979
transform 1 0 17848 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_175
timestamp 1606256979
transform 1 0 17204 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_180
timestamp 1606256979
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_186
timestamp 1606256979
transform 1 0 18216 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 1380 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_19
timestamp 1606256979
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1606256979
transform 1 0 3036 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1606256979
transform 1 0 3956 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_25
timestamp 1606256979
transform 1 0 3404 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_40
timestamp 1606256979
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1606256979
transform 1 0 5980 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1606256979
transform 1 0 4968 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1606256979
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1606256979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_51
timestamp 1606256979
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1606256979
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1606256979
transform 1 0 7820 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1606256979
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_82
timestamp 1606256979
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8832 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1606256979
transform 1 0 9844 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_93
timestamp 1606256979
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_104
timestamp 1606256979
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _20_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 11868 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1606256979
transform 1 0 10856 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1606256979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_115
timestamp 1606256979
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1606256979
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 14076 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_139
timestamp 1606256979
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1606256979
transform 1 0 15732 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_157
timestamp 1606256979
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606256979
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606256979
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1606256979
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_168
timestamp 1606256979
transform 1 0 16560 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_176
timestamp 1606256979
transform 1 0 17296 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1606256979
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1606256979
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1606256979
transform 1 0 1656 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1564 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2208 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1606256979
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1606256979
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_10
timestamp 1606256979
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_26
timestamp 1606256979
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_21
timestamp 1606256979
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606256979
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_21
timestamp 1606256979
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1606256979
transform 1 0 3680 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1606256979
transform 1 0 3220 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1606256979
transform 1 0 3220 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_37
timestamp 1606256979
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606256979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4692 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_41
timestamp 1606256979
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 5428 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606256979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5060 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_46
timestamp 1606256979
transform 1 0 5336 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_48
timestamp 1606256979
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606256979
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1606256979
transform 1 0 8464 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1606256979
transform 1 0 7084 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7912 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 7636 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_63
timestamp 1606256979
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_69
timestamp 1606256979
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_78
timestamp 1606256979
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_83
timestamp 1606256979
transform 1 0 8740 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9108 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9936 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606256979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1606256979
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1606256979
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_103
timestamp 1606256979
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_108
timestamp 1606256979
transform 1 0 11040 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_112
timestamp 1606256979
transform 1 0 11408 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 10764 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1606256979
transform 1 0 11316 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_123
timestamp 1606256979
transform 1 0 12420 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1606256979
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_116
timestamp 1606256979
transform 1 0 11776 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 11868 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606256979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1606256979
transform 1 0 12512 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12144 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1606256979
transform 1 0 14168 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13524 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 13800 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_136
timestamp 1606256979
transform 1 0 13616 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 1606256979
transform 1 0 14076 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_133
timestamp 1606256979
transform 1 0 13340 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_144
timestamp 1606256979
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1606256979
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1606256979
transform 1 0 14536 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15548 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606256979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1606256979
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_157
timestamp 1606256979
transform 1 0 15548 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_155
timestamp 1606256979
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_166
timestamp 1606256979
transform 1 0 16376 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_169
timestamp 1606256979
transform 1 0 16652 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_174
timestamp 1606256979
transform 1 0 17112 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_180
timestamp 1606256979
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_175
timestamp 1606256979
transform 1 0 17204 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1606256979
transform 1 0 17296 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1606256979
transform 1 0 17388 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1606256979
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_186
timestamp 1606256979
transform 1 0 18216 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606256979
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1606256979
transform 1 0 17848 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1606256979
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_188
timestamp 1606256979
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1606256979
transform 1 0 1656 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2300 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1606256979
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_10
timestamp 1606256979
transform 1 0 2024 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4048 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1606256979
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1606256979
transform 1 0 5704 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 6348 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_48
timestamp 1606256979
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_54
timestamp 1606256979
transform 1 0 6072 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7360 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_66
timestamp 1606256979
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1606256979
transform 1 0 9016 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 9752 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1606256979
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1606256979
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_93
timestamp 1606256979
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12512 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1606256979
transform 1 0 11500 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_110
timestamp 1606256979
transform 1 0 11224 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_122
timestamp 1606256979
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13524 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_133
timestamp 1606256979
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1606256979
transform 1 0 16284 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1606256979
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1606256979
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1606256979
transform 1 0 17848 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_174
timestamp 1606256979
transform 1 0 17112 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_186
timestamp 1606256979
transform 1 0 18216 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 1564 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1606256979
transform 1 0 3220 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1606256979
transform 1 0 3680 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 4692 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_21
timestamp 1606256979
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_26
timestamp 1606256979
transform 1 0 3496 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_37
timestamp 1606256979
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4968 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1606256979
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_62
timestamp 1606256979
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 8464 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 7084 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_9_74
timestamp 1606256979
transform 1 0 7912 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 10304 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_96
timestamp 1606256979
transform 1 0 9936 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 11960 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_116
timestamp 1606256979
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1606256979
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1606256979
transform 1 0 13432 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1606256979
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_143
timestamp 1606256979
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1606256979
transform 1 0 14536 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1606256979
transform 1 0 15548 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_155
timestamp 1606256979
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1606256979
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1606256979
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1606256979
transform 1 0 16560 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_177
timestamp 1606256979
transform 1 0 17388 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1606256979
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 2852 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1606256979
transform 1 0 1840 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1606256979
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1606256979
transform 1 0 1748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_17
timestamp 1606256979
transform 1 0 2668 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1606256979
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_28
timestamp 1606256979
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1606256979
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1606256979
transform 1 0 6072 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5060 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_52
timestamp 1606256979
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1606256979
transform 1 0 8648 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1606256979
transform 1 0 7084 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1606256979
transform 1 0 7636 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_63
timestamp 1606256979
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_69
timestamp 1606256979
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_80
timestamp 1606256979
transform 1 0 8464 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1606256979
transform 1 0 10672 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1606256979
transform 1 0 8924 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1606256979
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1606256979
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 11316 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_107
timestamp 1606256979
transform 1 0 10948 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1606256979
transform 1 0 12972 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1606256979
transform 1 0 14168 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_127
timestamp 1606256979
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_138
timestamp 1606256979
transform 1 0 13800 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 15272 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1606256979
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1606256979
transform 1 0 17940 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16928 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_170
timestamp 1606256979
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_181
timestamp 1606256979
transform 1 0 17756 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_187
timestamp 1606256979
transform 1 0 18308 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1380 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_19
timestamp 1606256979
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1606256979
transform 1 0 4048 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4876 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 3036 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_30
timestamp 1606256979
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_36
timestamp 1606256979
transform 1 0 4416 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_40
timestamp 1606256979
transform 1 0 4784 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1606256979
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1606256979
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7544 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 6992 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_67
timestamp 1606256979
transform 1 0 7268 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 9200 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_11_86
timestamp 1606256979
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1606256979
transform 1 0 11132 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_108
timestamp 1606256979
transform 1 0 11040 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1606256979
transform 1 0 11960 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1606256979
transform 1 0 13524 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_132
timestamp 1606256979
transform 1 0 13248 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_144
timestamp 1606256979
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 15824 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1606256979
transform 1 0 14536 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_155
timestamp 1606256979
transform 1 0 15364 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_159
timestamp 1606256979
transform 1 0 15732 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1606256979
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_176
timestamp 1606256979
transform 1 0 17296 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1606256979
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_188
timestamp 1606256979
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1606256979
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 2944 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 1932 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1606256979
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_18
timestamp 1606256979
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4048 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1606256979
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5704 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_48
timestamp 1606256979
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7360 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_66
timestamp 1606256979
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1606256979
transform 1 0 10488 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_84
timestamp 1606256979
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12328 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1606256979
transform 1 0 11316 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_120
timestamp 1606256979
transform 1 0 12144 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1606256979
transform 1 0 13340 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1606256979
transform 1 0 14168 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_131
timestamp 1606256979
transform 1 0 13156 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_136
timestamp 1606256979
transform 1 0 13616 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1606256979
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16100 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1606256979
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_157
timestamp 1606256979
transform 1 0 15548 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_179
timestamp 1606256979
transform 1 0 17572 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_187
timestamp 1606256979
transform 1 0 18308 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_6
timestamp 1606256979
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_8
timestamp 1606256979
transform 1 0 1840 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1606256979
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1606256979
transform 1 0 1840 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1606256979
transform 1 0 1472 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1606256979
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_17
timestamp 1606256979
transform 1 0 2668 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 2944 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2024 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1606256979
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_26
timestamp 1606256979
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1606256979
transform 1 0 3680 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_36
timestamp 1606256979
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_37
timestamp 1606256979
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 4600 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1606256979
transform 1 0 4692 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1606256979
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4876 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 5888 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_48
timestamp 1606256979
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606256979
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_50
timestamp 1606256979
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1606256979
transform 1 0 8648 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1606256979
transform 1 0 7636 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1606256979
transform 1 0 7636 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1606256979
transform 1 0 8464 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_68
timestamp 1606256979
transform 1 0 7360 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_80
timestamp 1606256979
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1606256979
transform 1 0 9292 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10120 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1606256979
transform 1 0 8924 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1606256979
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1606256979
transform 1 0 12236 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1606256979
transform 1 0 11316 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 11960 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1606256979
transform 1 0 10948 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1606256979
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_109
timestamp 1606256979
transform 1 0 11132 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_117
timestamp 1606256979
transform 1 0 11868 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1606256979
transform 1 0 14260 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 14168 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1606256979
transform 1 0 13248 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_139
timestamp 1606256979
transform 1 0 13892 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_130
timestamp 1606256979
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1606256979
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_158
timestamp 1606256979
transform 1 0 15640 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_146
timestamp 1606256979
transform 1 0 14536 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1606256979
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_163
timestamp 1606256979
transform 1 0 16100 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16928 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_175
timestamp 1606256979
transform 1 0 17204 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_184
timestamp 1606256979
transform 1 0 18032 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_171
timestamp 1606256979
transform 1 0 16836 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_188
timestamp 1606256979
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 1380 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1606256979
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1606256979
transform 1 0 3036 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 3680 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4692 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_25
timestamp 1606256979
transform 1 0 3404 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_37
timestamp 1606256979
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1606256979
transform 1 0 5704 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1606256979
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1606256979
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_62
timestamp 1606256979
transform 1 0 6808 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 7728 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_70
timestamp 1606256979
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 10672 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1606256979
transform 1 0 9384 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_88
timestamp 1606256979
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_99
timestamp 1606256979
transform 1 0 10212 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_103
timestamp 1606256979
transform 1 0 10580 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1606256979
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13432 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1606256979
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 16284 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1606256979
transform 1 0 15272 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_150
timestamp 1606256979
transform 1 0 14904 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_163
timestamp 1606256979
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1606256979
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1606256979
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_187
timestamp 1606256979
transform 1 0 18308 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1606256979
transform 1 0 1656 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 2300 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1606256979
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_10
timestamp 1606256979
transform 1 0 2024 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4232 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1606256979
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_32
timestamp 1606256979
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1606256979
transform 1 0 6440 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 5888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_50
timestamp 1606256979
transform 1 0 5704 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_55
timestamp 1606256979
transform 1 0 6164 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7912 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 7452 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_67
timestamp 1606256979
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_72
timestamp 1606256979
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606256979
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 12236 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 11408 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_109
timestamp 1606256979
transform 1 0 11132 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_115
timestamp 1606256979
transform 1 0 11684 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1606256979
transform 1 0 13892 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_137
timestamp 1606256979
transform 1 0 13708 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 15272 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_148
timestamp 1606256979
transform 1 0 14720 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1606256979
transform 1 0 16928 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1606256979
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_181
timestamp 1606256979
transform 1 0 17756 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1606256979
transform 1 0 18492 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 2576 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 1564 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1606256979
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_14
timestamp 1606256979
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 3588 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_25
timestamp 1606256979
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1606256979
transform 1 0 5244 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 5704 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_43
timestamp 1606256979
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_48
timestamp 1606256979
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1606256979
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_62
timestamp 1606256979
transform 1 0 6808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 7544 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1606256979
transform 1 0 9200 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9660 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10672 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_86
timestamp 1606256979
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_91
timestamp 1606256979
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_102
timestamp 1606256979
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1606256979
transform 1 0 12512 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1606256979
transform 1 0 11500 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1606256979
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_123
timestamp 1606256979
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1606256979
transform 1 0 13800 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_133
timestamp 1606256979
transform 1 0 13340 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_137
timestamp 1606256979
transform 1 0 13708 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15272 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_17_147
timestamp 1606256979
transform 1 0 14628 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_153
timestamp 1606256979
transform 1 0 15180 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1606256979
transform 1 0 16928 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_170
timestamp 1606256979
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1606256979
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_184
timestamp 1606256979
transform 1 0 18032 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 2944 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 1932 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1606256979
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_18
timestamp 1606256979
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 4508 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1606256979
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1606256979
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_36
timestamp 1606256979
transform 1 0 4416 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 5520 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6532 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_46
timestamp 1606256979
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_57
timestamp 1606256979
transform 1 0 6348 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1606256979
transform 1 0 8556 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1606256979
transform 1 0 7544 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_68
timestamp 1606256979
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_79
timestamp 1606256979
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1606256979
transform 1 0 9936 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1606256979
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_93
timestamp 1606256979
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1606256979
transform 1 0 11960 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10948 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_105
timestamp 1606256979
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_116
timestamp 1606256979
transform 1 0 11776 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1606256979
transform 1 0 13432 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1606256979
transform 1 0 13892 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_18_127
timestamp 1606256979
transform 1 0 12788 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_133
timestamp 1606256979
transform 1 0 13340 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_137
timestamp 1606256979
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15640 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_148
timestamp 1606256979
transform 1 0 14720 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1606256979
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1606256979
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16652 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1606256979
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_185
timestamp 1606256979
transform 1 0 18124 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1606256979
transform 1 0 18492 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1606256979
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1606256979
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1606256979
transform 1 0 1472 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1606256979
transform 1 0 1748 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_13
timestamp 1606256979
transform 1 0 2300 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_16
timestamp 1606256979
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1606256979
transform 1 0 2484 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 2760 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4784 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1606256979
transform 1 0 4784 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_34
timestamp 1606256979
transform 1 0 4232 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_24
timestamp 1606256979
transform 1 0 3312 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1606256979
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_32
timestamp 1606256979
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5888 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_56
timestamp 1606256979
transform 1 0 6256 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1606256979
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_49
timestamp 1606256979
transform 1 0 5612 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_61
timestamp 1606256979
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6900 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1606256979
transform 1 0 8556 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_19_78
timestamp 1606256979
transform 1 0 8280 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_79
timestamp 1606256979
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10580 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 8832 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10672 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_100
timestamp 1606256979
transform 1 0 10304 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1606256979
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1606256979
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 11868 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 12420 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_119
timestamp 1606256979
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_113
timestamp 1606256979
transform 1 0 11500 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 14260 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1606256979
transform 1 0 13524 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_139
timestamp 1606256979
transform 1 0 13892 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_133
timestamp 1606256979
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_144
timestamp 1606256979
transform 1 0 14352 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1606256979
transform 1 0 16284 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1606256979
transform 1 0 15916 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_159
timestamp 1606256979
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1606256979
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1606256979
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1606256979
transform 1 0 17480 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1606256979
transform 1 0 16928 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_170
timestamp 1606256979
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1606256979
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_184
timestamp 1606256979
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_174
timestamp 1606256979
transform 1 0 17112 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_187
timestamp 1606256979
transform 1 0 18308 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 2852 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1606256979
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_15
timestamp 1606256979
transform 1 0 2484 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1606256979
transform 1 0 4876 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1606256979
transform 1 0 3864 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_28
timestamp 1606256979
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_39
timestamp 1606256979
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_50
timestamp 1606256979
transform 1 0 5704 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_58
timestamp 1606256979
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_71
timestamp 1606256979
transform 1 0 7636 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_83
timestamp 1606256979
transform 1 0 8740 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1606256979
transform 1 0 9108 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1606256979
transform 1 0 10212 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_96
timestamp 1606256979
transform 1 0 9936 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 11316 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_108
timestamp 1606256979
transform 1 0 11040 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_117
timestamp 1606256979
transform 1 0 11868 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1606256979
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1606256979
transform 1 0 13524 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_132
timestamp 1606256979
transform 1 0 13248 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_144
timestamp 1606256979
transform 1 0 14352 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 15824 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1606256979
transform 1 0 14812 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_148
timestamp 1606256979
transform 1 0 14720 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_158
timestamp 1606256979
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1606256979
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1606256979
transform 1 0 17204 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_173
timestamp 1606256979
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1606256979
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_188
timestamp 1606256979
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1606256979
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1606256979
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4140 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606256979
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_32
timestamp 1606256979
transform 1 0 4048 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_42
timestamp 1606256979
transform 1 0 4968 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_54
timestamp 1606256979
transform 1 0 6072 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_63
timestamp 1606256979
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_75
timestamp 1606256979
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9752 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_87
timestamp 1606256979
transform 1 0 9108 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_103
timestamp 1606256979
transform 1 0 10580 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_115
timestamp 1606256979
transform 1 0 11684 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_123
timestamp 1606256979
transform 1 0 12420 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1606256979
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1606256979
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606256979
transform 1 0 15640 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 15364 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_149
timestamp 1606256979
transform 1 0 14812 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_153
timestamp 1606256979
transform 1 0 15180 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_156
timestamp 1606256979
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1606256979
transform 1 0 17020 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_171
timestamp 1606256979
transform 1 0 16836 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_182
timestamp 1606256979
transform 1 0 17848 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_187
timestamp 1606256979
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
<< labels >>
rlabel metal2 s 1122 16520 1178 17000 6 IO_ISOL_N
port 0 nsew default input
rlabel metal2 s 17590 0 17646 480 6 SC_IN_BOT
port 1 nsew default input
rlabel metal2 s 3330 16520 3386 17000 6 SC_IN_TOP
port 2 nsew default input
rlabel metal2 s 18510 0 18566 480 6 SC_OUT_BOT
port 3 nsew default tristate
rlabel metal2 s 5538 16520 5594 17000 6 SC_OUT_TOP
port 4 nsew default tristate
rlabel metal2 s 1214 0 1270 480 6 bottom_grid_pin_0_
port 5 nsew default tristate
rlabel metal2 s 10322 0 10378 480 6 bottom_grid_pin_10_
port 6 nsew default tristate
rlabel metal2 s 11242 0 11298 480 6 bottom_grid_pin_11_
port 7 nsew default tristate
rlabel metal2 s 12162 0 12218 480 6 bottom_grid_pin_12_
port 8 nsew default tristate
rlabel metal2 s 13082 0 13138 480 6 bottom_grid_pin_13_
port 9 nsew default tristate
rlabel metal2 s 13910 0 13966 480 6 bottom_grid_pin_14_
port 10 nsew default tristate
rlabel metal2 s 14830 0 14886 480 6 bottom_grid_pin_15_
port 11 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 bottom_grid_pin_1_
port 12 nsew default tristate
rlabel metal2 s 3054 0 3110 480 6 bottom_grid_pin_2_
port 13 nsew default tristate
rlabel metal2 s 3974 0 4030 480 6 bottom_grid_pin_3_
port 14 nsew default tristate
rlabel metal2 s 4894 0 4950 480 6 bottom_grid_pin_4_
port 15 nsew default tristate
rlabel metal2 s 5814 0 5870 480 6 bottom_grid_pin_5_
port 16 nsew default tristate
rlabel metal2 s 6734 0 6790 480 6 bottom_grid_pin_6_
port 17 nsew default tristate
rlabel metal2 s 7562 0 7618 480 6 bottom_grid_pin_7_
port 18 nsew default tristate
rlabel metal2 s 8482 0 8538 480 6 bottom_grid_pin_8_
port 19 nsew default tristate
rlabel metal2 s 9402 0 9458 480 6 bottom_grid_pin_9_
port 20 nsew default tristate
rlabel metal2 s 15750 0 15806 480 6 bottom_width_0_height_0__pin_0_
port 21 nsew default input
rlabel metal2 s 16670 0 16726 480 6 bottom_width_0_height_0__pin_1_lower
port 22 nsew default tristate
rlabel metal2 s 386 0 442 480 6 bottom_width_0_height_0__pin_1_upper
port 23 nsew default tristate
rlabel metal2 s 7746 16520 7802 17000 6 ccff_head
port 24 nsew default input
rlabel metal2 s 9954 16520 10010 17000 6 ccff_tail
port 25 nsew default tristate
rlabel metal3 s 0 8848 480 8968 6 chanx_left_in[0]
port 26 nsew default input
rlabel metal3 s 0 12928 480 13048 6 chanx_left_in[10]
port 27 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[11]
port 28 nsew default input
rlabel metal3 s 0 13744 480 13864 6 chanx_left_in[12]
port 29 nsew default input
rlabel metal3 s 0 14152 480 14272 6 chanx_left_in[13]
port 30 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[14]
port 31 nsew default input
rlabel metal3 s 0 14968 480 15088 6 chanx_left_in[15]
port 32 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[16]
port 33 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[17]
port 34 nsew default input
rlabel metal3 s 0 16192 480 16312 6 chanx_left_in[18]
port 35 nsew default input
rlabel metal3 s 0 16600 480 16720 6 chanx_left_in[19]
port 36 nsew default input
rlabel metal3 s 0 9256 480 9376 6 chanx_left_in[1]
port 37 nsew default input
rlabel metal3 s 0 9664 480 9784 6 chanx_left_in[2]
port 38 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[3]
port 39 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[4]
port 40 nsew default input
rlabel metal3 s 0 10888 480 11008 6 chanx_left_in[5]
port 41 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[6]
port 42 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[7]
port 43 nsew default input
rlabel metal3 s 0 12112 480 12232 6 chanx_left_in[8]
port 44 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[9]
port 45 nsew default input
rlabel metal3 s 0 552 480 672 6 chanx_left_out[0]
port 46 nsew default tristate
rlabel metal3 s 0 4632 480 4752 6 chanx_left_out[10]
port 47 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[11]
port 48 nsew default tristate
rlabel metal3 s 0 5448 480 5568 6 chanx_left_out[12]
port 49 nsew default tristate
rlabel metal3 s 0 5856 480 5976 6 chanx_left_out[13]
port 50 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[14]
port 51 nsew default tristate
rlabel metal3 s 0 6672 480 6792 6 chanx_left_out[15]
port 52 nsew default tristate
rlabel metal3 s 0 7080 480 7200 6 chanx_left_out[16]
port 53 nsew default tristate
rlabel metal3 s 0 7488 480 7608 6 chanx_left_out[17]
port 54 nsew default tristate
rlabel metal3 s 0 7896 480 8016 6 chanx_left_out[18]
port 55 nsew default tristate
rlabel metal3 s 0 8304 480 8424 6 chanx_left_out[19]
port 56 nsew default tristate
rlabel metal3 s 0 960 480 1080 6 chanx_left_out[1]
port 57 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 58 nsew default tristate
rlabel metal3 s 0 1776 480 1896 6 chanx_left_out[3]
port 59 nsew default tristate
rlabel metal3 s 0 2184 480 2304 6 chanx_left_out[4]
port 60 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[5]
port 61 nsew default tristate
rlabel metal3 s 0 3000 480 3120 6 chanx_left_out[6]
port 62 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 chanx_left_out[7]
port 63 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[8]
port 64 nsew default tristate
rlabel metal3 s 0 4224 480 4344 6 chanx_left_out[9]
port 65 nsew default tristate
rlabel metal3 s 19520 8576 20000 8696 6 chanx_right_in[0]
port 66 nsew default input
rlabel metal3 s 19520 12792 20000 12912 6 chanx_right_in[10]
port 67 nsew default input
rlabel metal3 s 19520 13200 20000 13320 6 chanx_right_in[11]
port 68 nsew default input
rlabel metal3 s 19520 13744 20000 13864 6 chanx_right_in[12]
port 69 nsew default input
rlabel metal3 s 19520 14152 20000 14272 6 chanx_right_in[13]
port 70 nsew default input
rlabel metal3 s 19520 14560 20000 14680 6 chanx_right_in[14]
port 71 nsew default input
rlabel metal3 s 19520 14968 20000 15088 6 chanx_right_in[15]
port 72 nsew default input
rlabel metal3 s 19520 15376 20000 15496 6 chanx_right_in[16]
port 73 nsew default input
rlabel metal3 s 19520 15784 20000 15904 6 chanx_right_in[17]
port 74 nsew default input
rlabel metal3 s 19520 16192 20000 16312 6 chanx_right_in[18]
port 75 nsew default input
rlabel metal3 s 19520 16600 20000 16720 6 chanx_right_in[19]
port 76 nsew default input
rlabel metal3 s 19520 8984 20000 9104 6 chanx_right_in[1]
port 77 nsew default input
rlabel metal3 s 19520 9392 20000 9512 6 chanx_right_in[2]
port 78 nsew default input
rlabel metal3 s 19520 9800 20000 9920 6 chanx_right_in[3]
port 79 nsew default input
rlabel metal3 s 19520 10344 20000 10464 6 chanx_right_in[4]
port 80 nsew default input
rlabel metal3 s 19520 10752 20000 10872 6 chanx_right_in[5]
port 81 nsew default input
rlabel metal3 s 19520 11160 20000 11280 6 chanx_right_in[6]
port 82 nsew default input
rlabel metal3 s 19520 11568 20000 11688 6 chanx_right_in[7]
port 83 nsew default input
rlabel metal3 s 19520 11976 20000 12096 6 chanx_right_in[8]
port 84 nsew default input
rlabel metal3 s 19520 12384 20000 12504 6 chanx_right_in[9]
port 85 nsew default input
rlabel metal3 s 19520 144 20000 264 6 chanx_right_out[0]
port 86 nsew default tristate
rlabel metal3 s 19520 4360 20000 4480 6 chanx_right_out[10]
port 87 nsew default tristate
rlabel metal3 s 19520 4768 20000 4888 6 chanx_right_out[11]
port 88 nsew default tristate
rlabel metal3 s 19520 5176 20000 5296 6 chanx_right_out[12]
port 89 nsew default tristate
rlabel metal3 s 19520 5584 20000 5704 6 chanx_right_out[13]
port 90 nsew default tristate
rlabel metal3 s 19520 5992 20000 6112 6 chanx_right_out[14]
port 91 nsew default tristate
rlabel metal3 s 19520 6400 20000 6520 6 chanx_right_out[15]
port 92 nsew default tristate
rlabel metal3 s 19520 6944 20000 7064 6 chanx_right_out[16]
port 93 nsew default tristate
rlabel metal3 s 19520 7352 20000 7472 6 chanx_right_out[17]
port 94 nsew default tristate
rlabel metal3 s 19520 7760 20000 7880 6 chanx_right_out[18]
port 95 nsew default tristate
rlabel metal3 s 19520 8168 20000 8288 6 chanx_right_out[19]
port 96 nsew default tristate
rlabel metal3 s 19520 552 20000 672 6 chanx_right_out[1]
port 97 nsew default tristate
rlabel metal3 s 19520 960 20000 1080 6 chanx_right_out[2]
port 98 nsew default tristate
rlabel metal3 s 19520 1368 20000 1488 6 chanx_right_out[3]
port 99 nsew default tristate
rlabel metal3 s 19520 1776 20000 1896 6 chanx_right_out[4]
port 100 nsew default tristate
rlabel metal3 s 19520 2184 20000 2304 6 chanx_right_out[5]
port 101 nsew default tristate
rlabel metal3 s 19520 2592 20000 2712 6 chanx_right_out[6]
port 102 nsew default tristate
rlabel metal3 s 19520 3000 20000 3120 6 chanx_right_out[7]
port 103 nsew default tristate
rlabel metal3 s 19520 3544 20000 3664 6 chanx_right_out[8]
port 104 nsew default tristate
rlabel metal3 s 19520 3952 20000 4072 6 chanx_right_out[9]
port 105 nsew default tristate
rlabel metal2 s 14370 16520 14426 17000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 106 nsew default tristate
rlabel metal2 s 16578 16520 16634 17000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 107 nsew default input
rlabel metal2 s 18786 16520 18842 17000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 108 nsew default tristate
rlabel metal2 s 19430 0 19486 480 6 prog_clk_0_S_in
port 109 nsew default input
rlabel metal3 s 0 144 480 264 6 prog_clk_0_W_out
port 110 nsew default tristate
rlabel metal2 s 12162 16520 12218 17000 6 top_grid_pin_0_
port 111 nsew default tristate
rlabel metal4 s 3909 2128 4229 14736 6 VPWR
port 112 nsew default input
rlabel metal4 s 6875 2128 7195 14736 6 VGND
port 113 nsew default input
<< properties >>
string FIXED_BBOX 0 0 20000 17000
<< end >>
