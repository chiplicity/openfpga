magic
tech sky130A
magscale 1 2
timestamp 1605110485
<< locali >>
rect 8401 13923 8435 14025
rect 24501 9435 24535 9605
rect 6561 2431 6595 2601
<< viali >>
rect 17049 20893 17083 20927
rect 8401 20757 8435 20791
rect 13553 20757 13587 20791
rect 23673 20757 23707 20791
rect 7113 20553 7147 20587
rect 21925 20553 21959 20587
rect 20637 20485 20671 20519
rect 16957 20417 16991 20451
rect 3525 20349 3559 20383
rect 8309 20349 8343 20383
rect 13553 20349 13587 20383
rect 16681 20349 16715 20383
rect 17417 20349 17451 20383
rect 19257 20349 19291 20383
rect 21741 20349 21775 20383
rect 22293 20349 22327 20383
rect 23673 20349 23707 20383
rect 26157 20349 26191 20383
rect 3433 20281 3467 20315
rect 3770 20281 3804 20315
rect 8554 20281 8588 20315
rect 13798 20281 13832 20315
rect 19165 20281 19199 20315
rect 19502 20281 19536 20315
rect 23489 20281 23523 20315
rect 23940 20281 23974 20315
rect 4905 20213 4939 20247
rect 8125 20213 8159 20247
rect 9689 20213 9723 20247
rect 13461 20213 13495 20247
rect 14933 20213 14967 20247
rect 25053 20213 25087 20247
rect 26341 20213 26375 20247
rect 26801 20213 26835 20247
rect 3525 20009 3559 20043
rect 6653 20009 6687 20043
rect 13737 20009 13771 20043
rect 15761 20009 15795 20043
rect 17693 20009 17727 20043
rect 19257 20009 19291 20043
rect 26709 20009 26743 20043
rect 17785 19941 17819 19975
rect 21802 19941 21836 19975
rect 5273 19873 5307 19907
rect 5540 19873 5574 19907
rect 8125 19873 8159 19907
rect 10800 19873 10834 19907
rect 11060 19873 11094 19907
rect 16129 19873 16163 19907
rect 26525 19873 26559 19907
rect 8217 19805 8251 19839
rect 8309 19805 8343 19839
rect 13829 19805 13863 19839
rect 14013 19805 14047 19839
rect 16221 19805 16255 19839
rect 16313 19805 16347 19839
rect 17877 19805 17911 19839
rect 21557 19805 21591 19839
rect 7573 19737 7607 19771
rect 7757 19737 7791 19771
rect 17325 19737 17359 19771
rect 3157 19669 3191 19703
rect 7205 19669 7239 19703
rect 8861 19669 8895 19703
rect 12173 19669 12207 19703
rect 13369 19669 13403 19703
rect 14473 19669 14507 19703
rect 22937 19669 22971 19703
rect 23765 19669 23799 19703
rect 25329 19669 25363 19703
rect 5641 19465 5675 19499
rect 8125 19465 8159 19499
rect 13093 19465 13127 19499
rect 13737 19465 13771 19499
rect 17693 19465 17727 19499
rect 21189 19465 21223 19499
rect 23489 19465 23523 19499
rect 2605 19397 2639 19431
rect 13461 19397 13495 19431
rect 17049 19397 17083 19431
rect 23673 19397 23707 19431
rect 24777 19397 24811 19431
rect 3709 19329 3743 19363
rect 7757 19329 7791 19363
rect 8769 19329 8803 19363
rect 9505 19329 9539 19363
rect 22661 19329 22695 19363
rect 24133 19329 24167 19363
rect 24317 19329 24351 19363
rect 25881 19329 25915 19363
rect 3433 19261 3467 19295
rect 4629 19261 4663 19295
rect 5365 19261 5399 19295
rect 6285 19261 6319 19295
rect 9229 19261 9263 19295
rect 10885 19261 10919 19295
rect 14381 19261 14415 19295
rect 21833 19261 21867 19295
rect 22385 19261 22419 19295
rect 25145 19261 25179 19295
rect 25605 19261 25639 19295
rect 26801 19261 26835 19295
rect 2973 19193 3007 19227
rect 7573 19193 7607 19227
rect 14197 19193 14231 19227
rect 14648 19193 14682 19227
rect 23121 19193 23155 19227
rect 24041 19193 24075 19227
rect 25697 19193 25731 19227
rect 3065 19125 3099 19159
rect 3525 19125 3559 19159
rect 6561 19125 6595 19159
rect 7113 19125 7147 19159
rect 7481 19125 7515 19159
rect 8861 19125 8895 19159
rect 9321 19125 9355 19159
rect 11161 19125 11195 19159
rect 15761 19125 15795 19159
rect 16313 19125 16347 19159
rect 17325 19125 17359 19159
rect 21557 19125 21591 19159
rect 22017 19125 22051 19159
rect 22477 19125 22511 19159
rect 25237 19125 25271 19159
rect 26617 19125 26651 19159
rect 3433 18921 3467 18955
rect 6193 18921 6227 18955
rect 7573 18921 7607 18955
rect 8309 18921 8343 18955
rect 13645 18921 13679 18955
rect 15853 18921 15887 18955
rect 16589 18921 16623 18955
rect 22109 18921 22143 18955
rect 22661 18921 22695 18955
rect 24409 18921 24443 18955
rect 4445 18853 4479 18887
rect 6929 18853 6963 18887
rect 10876 18853 10910 18887
rect 14105 18853 14139 18887
rect 16221 18853 16255 18887
rect 16957 18853 16991 18887
rect 22477 18853 22511 18887
rect 1768 18785 1802 18819
rect 14013 18785 14047 18819
rect 17049 18785 17083 18819
rect 18337 18785 18371 18819
rect 18593 18785 18627 18819
rect 23029 18785 23063 18819
rect 24777 18785 24811 18819
rect 24869 18785 24903 18819
rect 1501 18717 1535 18751
rect 4537 18717 4571 18751
rect 4721 18717 4755 18751
rect 7665 18717 7699 18751
rect 7849 18717 7883 18751
rect 10609 18717 10643 18751
rect 14197 18717 14231 18751
rect 17141 18717 17175 18751
rect 20913 18717 20947 18751
rect 23121 18717 23155 18751
rect 23305 18717 23339 18751
rect 23765 18717 23799 18751
rect 24961 18717 24995 18751
rect 2881 18581 2915 18615
rect 4077 18581 4111 18615
rect 7205 18581 7239 18615
rect 8953 18581 8987 18615
rect 9965 18581 9999 18615
rect 11989 18581 12023 18615
rect 19717 18581 19751 18615
rect 21373 18581 21407 18615
rect 1685 18377 1719 18411
rect 4537 18377 4571 18411
rect 6837 18377 6871 18411
rect 7849 18377 7883 18411
rect 9781 18377 9815 18411
rect 10885 18377 10919 18411
rect 13277 18377 13311 18411
rect 16589 18377 16623 18411
rect 17049 18377 17083 18411
rect 17325 18377 17359 18411
rect 17877 18377 17911 18411
rect 19349 18377 19383 18411
rect 21189 18377 21223 18411
rect 22753 18377 22787 18411
rect 27537 18377 27571 18411
rect 1961 18309 1995 18343
rect 2973 18309 3007 18343
rect 4169 18309 4203 18343
rect 6653 18309 6687 18343
rect 14105 18309 14139 18343
rect 19625 18309 19659 18343
rect 21373 18309 21407 18343
rect 23673 18309 23707 18343
rect 25145 18309 25179 18343
rect 2605 18241 2639 18275
rect 3525 18241 3559 18275
rect 3709 18241 3743 18275
rect 6285 18241 6319 18275
rect 7389 18241 7423 18275
rect 9689 18241 9723 18275
rect 10425 18241 10459 18275
rect 13645 18241 13679 18275
rect 14749 18241 14783 18275
rect 20269 18241 20303 18275
rect 20361 18241 20395 18275
rect 21925 18241 21959 18275
rect 24317 18241 24351 18275
rect 3433 18173 3467 18207
rect 7297 18173 7331 18207
rect 10149 18173 10183 18207
rect 20177 18173 20211 18207
rect 21741 18173 21775 18207
rect 24777 18173 24811 18207
rect 26157 18173 26191 18207
rect 7205 18105 7239 18139
rect 9321 18105 9355 18139
rect 10241 18105 10275 18139
rect 12909 18105 12943 18139
rect 21833 18105 21867 18139
rect 23121 18105 23155 18139
rect 24133 18105 24167 18139
rect 26402 18105 26436 18139
rect 3065 18037 3099 18071
rect 4813 18037 4847 18071
rect 11253 18037 11287 18071
rect 13921 18037 13955 18071
rect 14473 18037 14507 18071
rect 14565 18037 14599 18071
rect 15209 18037 15243 18071
rect 18429 18037 18463 18071
rect 18889 18037 18923 18071
rect 19809 18037 19843 18071
rect 23489 18037 23523 18071
rect 24041 18037 24075 18071
rect 25973 18037 26007 18071
rect 7573 17833 7607 17867
rect 8033 17833 8067 17867
rect 10333 17833 10367 17867
rect 13553 17833 13587 17867
rect 17601 17833 17635 17867
rect 19717 17833 19751 17867
rect 21373 17833 21407 17867
rect 23029 17833 23063 17867
rect 23397 17833 23431 17867
rect 24777 17833 24811 17867
rect 26249 17833 26283 17867
rect 7297 17765 7331 17799
rect 19625 17765 19659 17799
rect 22753 17765 22787 17799
rect 1409 17697 1443 17731
rect 5273 17697 5307 17731
rect 5529 17697 5563 17731
rect 8401 17697 8435 17731
rect 10701 17697 10735 17731
rect 14013 17697 14047 17731
rect 16221 17697 16255 17731
rect 16488 17697 16522 17731
rect 23765 17697 23799 17731
rect 23857 17697 23891 17731
rect 8493 17629 8527 17663
rect 8677 17629 8711 17663
rect 10793 17629 10827 17663
rect 10885 17629 10919 17663
rect 14105 17629 14139 17663
rect 14289 17629 14323 17663
rect 19809 17629 19843 17663
rect 23949 17629 23983 17663
rect 10057 17561 10091 17595
rect 13645 17561 13679 17595
rect 18245 17561 18279 17595
rect 1593 17493 1627 17527
rect 2881 17493 2915 17527
rect 3157 17493 3191 17527
rect 6653 17493 6687 17527
rect 16037 17493 16071 17527
rect 19257 17493 19291 17527
rect 24501 17493 24535 17527
rect 2053 17289 2087 17323
rect 5365 17289 5399 17323
rect 8769 17289 8803 17323
rect 9965 17289 9999 17323
rect 11345 17289 11379 17323
rect 12909 17289 12943 17323
rect 14473 17289 14507 17323
rect 17785 17289 17819 17323
rect 19717 17289 19751 17323
rect 20085 17289 20119 17323
rect 23121 17289 23155 17323
rect 2697 17221 2731 17255
rect 9505 17221 9539 17255
rect 13277 17221 13311 17255
rect 16037 17221 16071 17255
rect 17509 17221 17543 17255
rect 3249 17153 3283 17187
rect 3433 17153 3467 17187
rect 8493 17153 8527 17187
rect 10609 17153 10643 17187
rect 13553 17153 13587 17187
rect 15025 17153 15059 17187
rect 15485 17153 15519 17187
rect 16589 17153 16623 17187
rect 17049 17153 17083 17187
rect 18613 17153 18647 17187
rect 18797 17153 18831 17187
rect 19349 17153 19383 17187
rect 24685 17153 24719 17187
rect 1409 17085 1443 17119
rect 3157 17085 3191 17119
rect 5641 17085 5675 17119
rect 14841 17085 14875 17119
rect 16405 17085 16439 17119
rect 18521 17085 18555 17119
rect 23489 17085 23523 17119
rect 26433 17085 26467 17119
rect 26985 17085 27019 17119
rect 9873 17017 9907 17051
rect 10425 17017 10459 17051
rect 11069 17017 11103 17051
rect 15945 17017 15979 17051
rect 16497 17017 16531 17051
rect 22753 17017 22787 17051
rect 24501 17017 24535 17051
rect 1593 16949 1627 16983
rect 2789 16949 2823 16983
rect 8033 16949 8067 16983
rect 10333 16949 10367 16983
rect 13921 16949 13955 16983
rect 14381 16949 14415 16983
rect 14933 16949 14967 16983
rect 18153 16949 18187 16983
rect 23857 16949 23891 16983
rect 24041 16949 24075 16983
rect 24409 16949 24443 16983
rect 26617 16949 26651 16983
rect 1685 16745 1719 16779
rect 2421 16745 2455 16779
rect 4353 16745 4387 16779
rect 5273 16745 5307 16779
rect 5733 16745 5767 16779
rect 10333 16745 10367 16779
rect 13829 16745 13863 16779
rect 14565 16745 14599 16779
rect 15301 16745 15335 16779
rect 15761 16745 15795 16779
rect 16313 16745 16347 16779
rect 18613 16745 18647 16779
rect 19257 16745 19291 16779
rect 23489 16745 23523 16779
rect 2789 16677 2823 16711
rect 5641 16677 5675 16711
rect 10701 16677 10735 16711
rect 15669 16677 15703 16711
rect 6837 16609 6871 16643
rect 7104 16609 7138 16643
rect 10793 16609 10827 16643
rect 12705 16609 12739 16643
rect 21169 16609 21203 16643
rect 24409 16609 24443 16643
rect 2881 16541 2915 16575
rect 3065 16541 3099 16575
rect 5825 16541 5859 16575
rect 10885 16541 10919 16575
rect 12449 16541 12483 16575
rect 15853 16541 15887 16575
rect 18705 16541 18739 16575
rect 18797 16541 18831 16575
rect 20913 16541 20947 16575
rect 24501 16541 24535 16575
rect 24685 16541 24719 16575
rect 24041 16473 24075 16507
rect 8217 16405 8251 16439
rect 10057 16405 10091 16439
rect 18245 16405 18279 16439
rect 22293 16405 22327 16439
rect 3893 16201 3927 16235
rect 5365 16201 5399 16235
rect 7021 16201 7055 16235
rect 11161 16201 11195 16235
rect 15393 16201 15427 16235
rect 16037 16201 16071 16235
rect 17877 16201 17911 16235
rect 18705 16201 18739 16235
rect 21005 16201 21039 16235
rect 23949 16201 23983 16235
rect 25053 16201 25087 16235
rect 27261 16201 27295 16235
rect 2789 16133 2823 16167
rect 5733 16133 5767 16167
rect 7389 16133 7423 16167
rect 10241 16133 10275 16167
rect 15669 16133 15703 16167
rect 18337 16133 18371 16167
rect 19073 16133 19107 16167
rect 21281 16133 21315 16167
rect 3433 16065 3467 16099
rect 4537 16065 4571 16099
rect 6009 16065 6043 16099
rect 19625 16065 19659 16099
rect 19717 16065 19751 16099
rect 24593 16065 24627 16099
rect 1409 15997 1443 16031
rect 8861 15997 8895 16031
rect 19533 15997 19567 16031
rect 23121 15997 23155 16031
rect 24317 15997 24351 16031
rect 25881 15997 25915 16031
rect 1676 15929 1710 15963
rect 3801 15929 3835 15963
rect 4261 15929 4295 15963
rect 8769 15929 8803 15963
rect 9106 15929 9140 15963
rect 10885 15929 10919 15963
rect 26126 15929 26160 15963
rect 4353 15861 4387 15895
rect 4905 15861 4939 15895
rect 12633 15861 12667 15895
rect 13001 15861 13035 15895
rect 19165 15861 19199 15895
rect 23489 15861 23523 15895
rect 24409 15861 24443 15895
rect 25697 15861 25731 15895
rect 1961 15657 1995 15691
rect 2513 15657 2547 15691
rect 2881 15657 2915 15691
rect 4077 15657 4111 15691
rect 10425 15657 10459 15691
rect 17785 15657 17819 15691
rect 18061 15657 18095 15691
rect 19165 15657 19199 15691
rect 24133 15657 24167 15691
rect 24869 15657 24903 15691
rect 25973 15657 26007 15691
rect 4445 15589 4479 15623
rect 11590 15589 11624 15623
rect 21986 15589 22020 15623
rect 9413 15521 9447 15555
rect 15301 15521 15335 15555
rect 15557 15521 15591 15555
rect 17969 15521 18003 15555
rect 18429 15521 18463 15555
rect 21741 15521 21775 15555
rect 26525 15521 26559 15555
rect 4537 15453 4571 15487
rect 4721 15453 4755 15487
rect 11345 15453 11379 15487
rect 18521 15453 18555 15487
rect 18613 15453 18647 15487
rect 1685 15385 1719 15419
rect 7757 15317 7791 15351
rect 8861 15317 8895 15351
rect 9229 15317 9263 15351
rect 12725 15317 12759 15351
rect 16681 15317 16715 15351
rect 23121 15317 23155 15351
rect 24501 15317 24535 15351
rect 26709 15317 26743 15351
rect 1685 15113 1719 15147
rect 4445 15113 4479 15147
rect 6469 15113 6503 15147
rect 7113 15113 7147 15147
rect 9045 15113 9079 15147
rect 9689 15113 9723 15147
rect 11713 15113 11747 15147
rect 15393 15113 15427 15147
rect 15761 15113 15795 15147
rect 17509 15113 17543 15147
rect 18337 15113 18371 15147
rect 20361 15113 20395 15147
rect 21373 15113 21407 15147
rect 21465 15113 21499 15147
rect 21925 15113 21959 15147
rect 26525 15113 26559 15147
rect 17877 15045 17911 15079
rect 7665 14977 7699 15011
rect 24501 14977 24535 15011
rect 25237 14977 25271 15011
rect 6653 14909 6687 14943
rect 7932 14909 7966 14943
rect 18981 14909 19015 14943
rect 21649 14909 21683 14943
rect 22293 14909 22327 14943
rect 7573 14841 7607 14875
rect 19226 14841 19260 14875
rect 24133 14841 24167 14875
rect 24961 14841 24995 14875
rect 4169 14773 4203 14807
rect 4905 14773 4939 14807
rect 11345 14773 11379 14807
rect 18889 14773 18923 14807
rect 24593 14773 24627 14807
rect 25053 14773 25087 14807
rect 6561 14569 6595 14603
rect 18153 14569 18187 14603
rect 18337 14569 18371 14603
rect 19901 14569 19935 14603
rect 24685 14569 24719 14603
rect 1746 14501 1780 14535
rect 11161 14501 11195 14535
rect 11713 14501 11747 14535
rect 15568 14501 15602 14535
rect 19441 14501 19475 14535
rect 22109 14501 22143 14535
rect 22744 14501 22778 14535
rect 5181 14433 5215 14467
rect 5448 14433 5482 14467
rect 8033 14433 8067 14467
rect 11621 14433 11655 14467
rect 15301 14433 15335 14467
rect 18705 14433 18739 14467
rect 20085 14433 20119 14467
rect 22477 14433 22511 14467
rect 1501 14365 1535 14399
rect 8125 14365 8159 14399
rect 8217 14365 8251 14399
rect 11805 14365 11839 14399
rect 12541 14365 12575 14399
rect 12817 14365 12851 14399
rect 18797 14365 18831 14399
rect 18889 14365 18923 14399
rect 10793 14297 10827 14331
rect 11253 14297 11287 14331
rect 2881 14229 2915 14263
rect 4353 14229 4387 14263
rect 7573 14229 7607 14263
rect 7665 14229 7699 14263
rect 9229 14229 9263 14263
rect 14289 14229 14323 14263
rect 16681 14229 16715 14263
rect 23857 14229 23891 14263
rect 4077 14025 4111 14059
rect 5641 14025 5675 14059
rect 8401 14025 8435 14059
rect 8677 14025 8711 14059
rect 10701 14025 10735 14059
rect 12449 14025 12483 14059
rect 15393 14025 15427 14059
rect 17785 14025 17819 14059
rect 19625 14025 19659 14059
rect 21925 14025 21959 14059
rect 23121 14025 23155 14059
rect 27537 14025 27571 14059
rect 5365 13957 5399 13991
rect 7573 13957 7607 13991
rect 9137 13957 9171 13991
rect 10241 13957 10275 13991
rect 12265 13957 12299 13991
rect 14289 13957 14323 13991
rect 15669 13957 15703 13991
rect 22017 13957 22051 13991
rect 2329 13889 2363 13923
rect 3249 13889 3283 13923
rect 3801 13889 3835 13923
rect 4813 13889 4847 13923
rect 7481 13889 7515 13923
rect 8033 13889 8067 13923
rect 8217 13889 8251 13923
rect 8401 13889 8435 13923
rect 9597 13889 9631 13923
rect 9689 13889 9723 13923
rect 11253 13889 11287 13923
rect 11437 13889 11471 13923
rect 12909 13889 12943 13923
rect 13001 13889 13035 13923
rect 14197 13889 14231 13923
rect 14933 13889 14967 13923
rect 18245 13889 18279 13923
rect 22477 13889 22511 13923
rect 22661 13889 22695 13923
rect 24225 13889 24259 13923
rect 1593 13821 1627 13855
rect 2237 13821 2271 13855
rect 4721 13821 4755 13855
rect 7113 13821 7147 13855
rect 9045 13821 9079 13855
rect 9505 13821 9539 13855
rect 11161 13821 11195 13855
rect 14749 13821 14783 13855
rect 20269 13821 20303 13855
rect 24133 13821 24167 13855
rect 26157 13821 26191 13855
rect 4629 13753 4663 13787
rect 11805 13753 11839 13787
rect 12817 13753 12851 13787
rect 13829 13753 13863 13787
rect 14657 13753 14691 13787
rect 17509 13753 17543 13787
rect 18490 13753 18524 13787
rect 26402 13753 26436 13787
rect 1777 13685 1811 13719
rect 2145 13685 2179 13719
rect 2789 13685 2823 13719
rect 4261 13685 4295 13719
rect 7941 13685 7975 13719
rect 10793 13685 10827 13719
rect 22385 13685 22419 13719
rect 23489 13685 23523 13719
rect 23673 13685 23707 13719
rect 24041 13685 24075 13719
rect 26065 13685 26099 13719
rect 1685 13481 1719 13515
rect 2237 13481 2271 13515
rect 2789 13481 2823 13515
rect 6837 13481 6871 13515
rect 7573 13481 7607 13515
rect 8033 13481 8067 13515
rect 9137 13481 9171 13515
rect 9689 13481 9723 13515
rect 10885 13481 10919 13515
rect 11345 13481 11379 13515
rect 11713 13481 11747 13515
rect 12173 13481 12207 13515
rect 13645 13481 13679 13515
rect 15301 13481 15335 13515
rect 15669 13481 15703 13515
rect 18797 13481 18831 13515
rect 22569 13481 22603 13515
rect 24041 13481 24075 13515
rect 24869 13481 24903 13515
rect 26249 13481 26283 13515
rect 4721 13413 4755 13447
rect 12081 13413 12115 13447
rect 14105 13413 14139 13447
rect 19073 13413 19107 13447
rect 25329 13413 25363 13447
rect 2145 13345 2179 13379
rect 4629 13345 4663 13379
rect 8401 13345 8435 13379
rect 10057 13345 10091 13379
rect 14013 13345 14047 13379
rect 25237 13345 25271 13379
rect 2421 13277 2455 13311
rect 4813 13277 4847 13311
rect 10149 13277 10183 13311
rect 10241 13277 10275 13311
rect 12265 13277 12299 13311
rect 14289 13277 14323 13311
rect 15761 13277 15795 13311
rect 15945 13277 15979 13311
rect 25513 13277 25547 13311
rect 8217 13209 8251 13243
rect 1777 13141 1811 13175
rect 3157 13141 3191 13175
rect 3709 13141 3743 13175
rect 4261 13141 4295 13175
rect 18429 13141 18463 13175
rect 22109 13141 22143 13175
rect 23765 13141 23799 13175
rect 3525 12937 3559 12971
rect 4721 12937 4755 12971
rect 8769 12937 8803 12971
rect 10425 12937 10459 12971
rect 11345 12937 11379 12971
rect 12173 12937 12207 12971
rect 13645 12937 13679 12971
rect 16037 12937 16071 12971
rect 17877 12937 17911 12971
rect 24225 12937 24259 12971
rect 25513 12937 25547 12971
rect 26525 12937 26559 12971
rect 5089 12869 5123 12903
rect 11805 12869 11839 12903
rect 14289 12869 14323 12903
rect 15761 12869 15795 12903
rect 24685 12869 24719 12903
rect 2697 12801 2731 12835
rect 3065 12801 3099 12835
rect 4169 12801 4203 12835
rect 6837 12801 6871 12835
rect 10149 12801 10183 12835
rect 14933 12801 14967 12835
rect 18613 12801 18647 12835
rect 20453 12801 20487 12835
rect 26065 12801 26099 12835
rect 2421 12733 2455 12767
rect 4077 12733 4111 12767
rect 13277 12733 13311 12767
rect 25053 12733 25087 12767
rect 25973 12733 26007 12767
rect 2513 12665 2547 12699
rect 3985 12665 4019 12699
rect 5365 12665 5399 12699
rect 6653 12665 6687 12699
rect 7082 12665 7116 12699
rect 17509 12665 17543 12699
rect 18521 12665 18555 12699
rect 20361 12665 20395 12699
rect 20720 12665 20754 12699
rect 25329 12665 25363 12699
rect 25881 12665 25915 12699
rect 1869 12597 1903 12631
rect 2053 12597 2087 12631
rect 3617 12597 3651 12631
rect 8217 12597 8251 12631
rect 9689 12597 9723 12631
rect 14197 12597 14231 12631
rect 14657 12597 14691 12631
rect 14749 12597 14783 12631
rect 15393 12597 15427 12631
rect 18061 12597 18095 12631
rect 18429 12597 18463 12631
rect 19165 12597 19199 12631
rect 21833 12597 21867 12631
rect 3065 12393 3099 12427
rect 13737 12393 13771 12427
rect 19165 12393 19199 12427
rect 20453 12393 20487 12427
rect 20913 12393 20947 12427
rect 26985 12393 27019 12427
rect 18030 12325 18064 12359
rect 2329 12257 2363 12291
rect 2421 12257 2455 12291
rect 4517 12257 4551 12291
rect 10609 12257 10643 12291
rect 15669 12257 15703 12291
rect 17785 12257 17819 12291
rect 21281 12257 21315 12291
rect 25237 12257 25271 12291
rect 25329 12257 25363 12291
rect 26893 12257 26927 12291
rect 1869 12189 1903 12223
rect 2605 12189 2639 12223
rect 3617 12189 3651 12223
rect 4261 12189 4295 12223
rect 10701 12189 10735 12223
rect 10793 12189 10827 12223
rect 15761 12189 15795 12223
rect 15945 12189 15979 12223
rect 21373 12189 21407 12223
rect 21557 12189 21591 12223
rect 22477 12189 22511 12223
rect 25513 12189 25547 12223
rect 27077 12189 27111 12223
rect 5641 12121 5675 12155
rect 14749 12121 14783 12155
rect 15301 12121 15335 12155
rect 24777 12121 24811 12155
rect 25973 12121 26007 12155
rect 1961 12053 1995 12087
rect 6929 12053 6963 12087
rect 10241 12053 10275 12087
rect 14289 12053 14323 12087
rect 16313 12053 16347 12087
rect 24225 12053 24259 12087
rect 24869 12053 24903 12087
rect 26525 12053 26559 12087
rect 27537 12053 27571 12087
rect 1685 11849 1719 11883
rect 3157 11849 3191 11883
rect 3985 11849 4019 11883
rect 4905 11849 4939 11883
rect 6561 11849 6595 11883
rect 10793 11849 10827 11883
rect 15117 11849 15151 11883
rect 16681 11849 16715 11883
rect 21465 11849 21499 11883
rect 24133 11849 24167 11883
rect 26709 11849 26743 11883
rect 4353 11781 4387 11815
rect 17509 11781 17543 11815
rect 20637 11781 20671 11815
rect 25605 11781 25639 11815
rect 26249 11781 26283 11815
rect 2421 11713 2455 11747
rect 4445 11713 4479 11747
rect 7297 11713 7331 11747
rect 7389 11713 7423 11747
rect 8493 11713 8527 11747
rect 10977 11713 11011 11747
rect 13645 11713 13679 11747
rect 16129 11713 16163 11747
rect 16313 11713 16347 11747
rect 17877 11713 17911 11747
rect 19073 11713 19107 11747
rect 21005 11713 21039 11747
rect 22109 11713 22143 11747
rect 27169 11713 27203 11747
rect 27353 11713 27387 11747
rect 27721 11713 27755 11747
rect 3341 11645 3375 11679
rect 13829 11645 13863 11679
rect 16037 11645 16071 11679
rect 17049 11645 17083 11679
rect 21281 11645 21315 11679
rect 21833 11645 21867 11679
rect 24225 11645 24259 11679
rect 24492 11645 24526 11679
rect 27077 11645 27111 11679
rect 6285 11577 6319 11611
rect 8738 11577 8772 11611
rect 18337 11577 18371 11611
rect 18797 11577 18831 11611
rect 20269 11577 20303 11611
rect 1777 11509 1811 11543
rect 2145 11509 2179 11543
rect 2237 11509 2271 11543
rect 2881 11509 2915 11543
rect 3525 11509 3559 11543
rect 6837 11509 6871 11543
rect 7205 11509 7239 11543
rect 8309 11509 8343 11543
rect 9873 11509 9907 11543
rect 10425 11509 10459 11543
rect 15669 11509 15703 11543
rect 18429 11509 18463 11543
rect 18889 11509 18923 11543
rect 19441 11509 19475 11543
rect 21925 11509 21959 11543
rect 26525 11509 26559 11543
rect 1961 11305 1995 11339
rect 3341 11305 3375 11339
rect 6561 11305 6595 11339
rect 8493 11305 8527 11339
rect 9689 11305 9723 11339
rect 16497 11305 16531 11339
rect 16773 11305 16807 11339
rect 17877 11305 17911 11339
rect 21189 11305 21223 11339
rect 21649 11305 21683 11339
rect 22017 11305 22051 11339
rect 24317 11305 24351 11339
rect 26709 11305 26743 11339
rect 27077 11305 27111 11339
rect 27445 11305 27479 11339
rect 27629 11305 27663 11339
rect 1685 11237 1719 11271
rect 3065 11237 3099 11271
rect 17141 11237 17175 11271
rect 24961 11237 24995 11271
rect 2329 11169 2363 11203
rect 6929 11169 6963 11203
rect 10057 11169 10091 11203
rect 12716 11169 12750 11203
rect 16129 11169 16163 11203
rect 18705 11169 18739 11203
rect 22109 11169 22143 11203
rect 25329 11169 25363 11203
rect 26525 11169 26559 11203
rect 2421 11101 2455 11135
rect 2513 11101 2547 11135
rect 7021 11101 7055 11135
rect 7113 11101 7147 11135
rect 10149 11101 10183 11135
rect 10241 11101 10275 11135
rect 12449 11101 12483 11135
rect 15301 11101 15335 11135
rect 17233 11101 17267 11135
rect 17417 11101 17451 11135
rect 18797 11101 18831 11135
rect 18889 11101 18923 11135
rect 22293 11101 22327 11135
rect 15853 11033 15887 11067
rect 18337 11033 18371 11067
rect 19441 11033 19475 11067
rect 21465 11033 21499 11067
rect 25513 11033 25547 11067
rect 7665 10965 7699 10999
rect 10701 10965 10735 10999
rect 13829 10965 13863 10999
rect 14473 10965 14507 10999
rect 2053 10761 2087 10795
rect 2421 10761 2455 10795
rect 7113 10761 7147 10795
rect 8861 10761 8895 10795
rect 10057 10761 10091 10795
rect 11069 10761 11103 10795
rect 12725 10761 12759 10795
rect 14197 10761 14231 10795
rect 15301 10761 15335 10795
rect 16957 10761 16991 10795
rect 17509 10761 17543 10795
rect 18889 10761 18923 10795
rect 21741 10761 21775 10795
rect 22109 10761 22143 10795
rect 25329 10761 25363 10795
rect 27353 10761 27387 10795
rect 2697 10693 2731 10727
rect 9137 10693 9171 10727
rect 14289 10693 14323 10727
rect 15853 10693 15887 10727
rect 7665 10625 7699 10659
rect 9505 10625 9539 10659
rect 10609 10625 10643 10659
rect 14933 10625 14967 10659
rect 16405 10625 16439 10659
rect 19441 10625 19475 10659
rect 1409 10557 1443 10591
rect 3065 10557 3099 10591
rect 3321 10557 3355 10591
rect 6653 10557 6687 10591
rect 7481 10557 7515 10591
rect 14657 10557 14691 10591
rect 16221 10557 16255 10591
rect 18429 10557 18463 10591
rect 26433 10557 26467 10591
rect 26985 10557 27019 10591
rect 27537 10557 27571 10591
rect 28089 10557 28123 10591
rect 5917 10489 5951 10523
rect 10517 10489 10551 10523
rect 13829 10489 13863 10523
rect 14749 10489 14783 10523
rect 15761 10489 15795 10523
rect 16313 10489 16347 10523
rect 17877 10489 17911 10523
rect 19257 10489 19291 10523
rect 1593 10421 1627 10455
rect 4445 10421 4479 10455
rect 6285 10421 6319 10455
rect 7573 10421 7607 10455
rect 9873 10421 9907 10455
rect 10425 10421 10459 10455
rect 13093 10421 13127 10455
rect 18705 10421 18739 10455
rect 19349 10421 19383 10455
rect 22477 10421 22511 10455
rect 23673 10421 23707 10455
rect 26617 10421 26651 10455
rect 27721 10421 27755 10455
rect 2053 10217 2087 10251
rect 2605 10217 2639 10251
rect 3157 10217 3191 10251
rect 6653 10217 6687 10251
rect 6929 10217 6963 10251
rect 7205 10217 7239 10251
rect 11897 10217 11931 10251
rect 15301 10217 15335 10251
rect 16313 10217 16347 10251
rect 16865 10217 16899 10251
rect 17233 10217 17267 10251
rect 18429 10217 18463 10251
rect 18797 10217 18831 10251
rect 19165 10217 19199 10251
rect 22753 10217 22787 10251
rect 24225 10217 24259 10251
rect 1961 10149 1995 10183
rect 3433 10149 3467 10183
rect 7573 10149 7607 10183
rect 9413 10149 9447 10183
rect 10762 10149 10796 10183
rect 13921 10149 13955 10183
rect 24317 10149 24351 10183
rect 8953 10081 8987 10115
rect 13829 10081 13863 10115
rect 15669 10081 15703 10115
rect 19257 10081 19291 10115
rect 20545 10081 20579 10115
rect 21629 10081 21663 10115
rect 26525 10081 26559 10115
rect 2237 10013 2271 10047
rect 7665 10013 7699 10047
rect 7757 10013 7791 10047
rect 10517 10013 10551 10047
rect 14013 10013 14047 10047
rect 15761 10013 15795 10047
rect 15945 10013 15979 10047
rect 19441 10013 19475 10047
rect 21373 10013 21407 10047
rect 24409 10013 24443 10047
rect 23857 9945 23891 9979
rect 1593 9877 1627 9911
rect 8309 9877 8343 9911
rect 8769 9877 8803 9911
rect 10057 9877 10091 9911
rect 13277 9877 13311 9911
rect 13461 9877 13495 9911
rect 20361 9877 20395 9911
rect 23765 9877 23799 9911
rect 26709 9877 26743 9911
rect 2329 9673 2363 9707
rect 3617 9673 3651 9707
rect 6561 9673 6595 9707
rect 7757 9673 7791 9707
rect 15393 9673 15427 9707
rect 16129 9673 16163 9707
rect 20453 9673 20487 9707
rect 24685 9673 24719 9707
rect 27537 9673 27571 9707
rect 3157 9605 3191 9639
rect 9321 9605 9355 9639
rect 12725 9605 12759 9639
rect 18797 9605 18831 9639
rect 23673 9605 23707 9639
rect 24501 9605 24535 9639
rect 26985 9605 27019 9639
rect 4077 9537 4111 9571
rect 7297 9537 7331 9571
rect 8309 9537 8343 9571
rect 9965 9537 9999 9571
rect 19441 9537 19475 9571
rect 22477 9537 22511 9571
rect 22569 9537 22603 9571
rect 23121 9537 23155 9571
rect 23489 9537 23523 9571
rect 24225 9537 24259 9571
rect 1409 9469 1443 9503
rect 2513 9469 2547 9503
rect 4169 9469 4203 9503
rect 4436 9469 4470 9503
rect 8217 9469 8251 9503
rect 9229 9469 9263 9503
rect 13185 9469 13219 9503
rect 19165 9469 19199 9503
rect 22385 9469 22419 9503
rect 24041 9469 24075 9503
rect 25605 9469 25639 9503
rect 2053 9401 2087 9435
rect 8769 9401 8803 9435
rect 10885 9401 10919 9435
rect 13452 9401 13486 9435
rect 19901 9401 19935 9435
rect 21925 9401 21959 9435
rect 24501 9401 24535 9435
rect 25145 9401 25179 9435
rect 25513 9401 25547 9435
rect 25872 9401 25906 9435
rect 1593 9333 1627 9367
rect 2697 9333 2731 9367
rect 5549 9333 5583 9367
rect 7573 9333 7607 9367
rect 8125 9333 8159 9367
rect 9689 9333 9723 9367
rect 9781 9333 9815 9367
rect 10609 9333 10643 9367
rect 13093 9333 13127 9367
rect 14565 9333 14599 9367
rect 15669 9333 15703 9367
rect 18245 9333 18279 9367
rect 18705 9333 18739 9367
rect 19257 9333 19291 9367
rect 21097 9333 21131 9367
rect 21465 9333 21499 9367
rect 22017 9333 22051 9367
rect 24133 9333 24167 9367
rect 1961 9129 1995 9163
rect 4537 9129 4571 9163
rect 7481 9129 7515 9163
rect 7757 9129 7791 9163
rect 8217 9129 8251 9163
rect 8861 9129 8895 9163
rect 13645 9129 13679 9163
rect 18889 9129 18923 9163
rect 19625 9129 19659 9163
rect 22201 9129 22235 9163
rect 22569 9129 22603 9163
rect 26709 9129 26743 9163
rect 2329 9061 2363 9095
rect 13277 9061 13311 9095
rect 1409 8993 1443 9027
rect 7113 8993 7147 9027
rect 8125 8993 8159 9027
rect 10609 8993 10643 9027
rect 17029 8993 17063 9027
rect 21833 8993 21867 9027
rect 23581 8993 23615 9027
rect 26525 8993 26559 9027
rect 8401 8925 8435 8959
rect 16773 8925 16807 8959
rect 23673 8925 23707 8959
rect 23857 8925 23891 8959
rect 9321 8857 9355 8891
rect 1593 8789 1627 8823
rect 6929 8789 6963 8823
rect 10425 8789 10459 8823
rect 14657 8789 14691 8823
rect 18153 8789 18187 8823
rect 19257 8789 19291 8823
rect 21649 8789 21683 8823
rect 23213 8789 23247 8823
rect 24225 8789 24259 8823
rect 25697 8789 25731 8823
rect 2053 8585 2087 8619
rect 4261 8585 4295 8619
rect 7113 8585 7147 8619
rect 7849 8585 7883 8619
rect 8585 8585 8619 8619
rect 11161 8585 11195 8619
rect 14473 8585 14507 8619
rect 16037 8585 16071 8619
rect 16865 8585 16899 8619
rect 19349 8585 19383 8619
rect 21465 8585 21499 8619
rect 22017 8585 22051 8619
rect 1593 8517 1627 8551
rect 17141 8517 17175 8551
rect 18797 8517 18831 8551
rect 23213 8517 23247 8551
rect 23673 8517 23707 8551
rect 2421 8449 2455 8483
rect 3985 8449 4019 8483
rect 5089 8449 5123 8483
rect 22937 8449 22971 8483
rect 24225 8449 24259 8483
rect 1409 8381 1443 8415
rect 4905 8381 4939 8415
rect 9781 8381 9815 8415
rect 14657 8381 14691 8415
rect 14913 8381 14947 8415
rect 18981 8381 19015 8415
rect 20085 8381 20119 8415
rect 4813 8313 4847 8347
rect 9689 8313 9723 8347
rect 10026 8313 10060 8347
rect 19993 8313 20027 8347
rect 20330 8313 20364 8347
rect 24041 8313 24075 8347
rect 25053 8313 25087 8347
rect 26525 8313 26559 8347
rect 4445 8245 4479 8279
rect 8125 8245 8159 8279
rect 9321 8245 9355 8279
rect 24133 8245 24167 8279
rect 24685 8245 24719 8279
rect 1593 8041 1627 8075
rect 4537 8041 4571 8075
rect 10517 8041 10551 8075
rect 21557 8041 21591 8075
rect 23305 8041 23339 8075
rect 24041 8041 24075 8075
rect 24409 8041 24443 8075
rect 26709 8041 26743 8075
rect 5978 7973 6012 8007
rect 23765 7973 23799 8007
rect 1409 7905 1443 7939
rect 4445 7905 4479 7939
rect 11693 7905 11727 7939
rect 16313 7905 16347 7939
rect 21649 7905 21683 7939
rect 26525 7905 26559 7939
rect 4629 7837 4663 7871
rect 5733 7837 5767 7871
rect 11437 7837 11471 7871
rect 16405 7837 16439 7871
rect 16589 7837 16623 7871
rect 21741 7837 21775 7871
rect 24501 7837 24535 7871
rect 24685 7837 24719 7871
rect 1961 7701 1995 7735
rect 4077 7701 4111 7735
rect 7113 7701 7147 7735
rect 12817 7701 12851 7735
rect 14565 7701 14599 7735
rect 15945 7701 15979 7735
rect 20177 7701 20211 7735
rect 21189 7701 21223 7735
rect 25053 7701 25087 7735
rect 26157 7701 26191 7735
rect 4169 7497 4203 7531
rect 4813 7497 4847 7531
rect 5733 7497 5767 7531
rect 10149 7497 10183 7531
rect 11529 7497 11563 7531
rect 21281 7497 21315 7531
rect 21833 7497 21867 7531
rect 24409 7497 24443 7531
rect 25513 7497 25547 7531
rect 27537 7497 27571 7531
rect 6837 7429 6871 7463
rect 14473 7429 14507 7463
rect 16129 7429 16163 7463
rect 17509 7429 17543 7463
rect 24225 7429 24259 7463
rect 7389 7361 7423 7395
rect 13553 7361 13587 7395
rect 15025 7361 15059 7395
rect 16773 7361 16807 7395
rect 19809 7361 19843 7395
rect 23489 7361 23523 7395
rect 25053 7361 25087 7395
rect 26157 7361 26191 7395
rect 1501 7293 1535 7327
rect 5365 7293 5399 7327
rect 6653 7293 6687 7327
rect 7297 7293 7331 7327
rect 8769 7293 8803 7327
rect 11805 7293 11839 7327
rect 17233 7293 17267 7327
rect 19901 7293 19935 7327
rect 20168 7293 20202 7327
rect 24869 7293 24903 7327
rect 25973 7293 26007 7327
rect 1768 7225 1802 7259
rect 4445 7225 4479 7259
rect 6193 7225 6227 7259
rect 8677 7225 8711 7259
rect 9014 7225 9048 7259
rect 12817 7225 12851 7259
rect 13277 7225 13311 7259
rect 14381 7225 14415 7259
rect 15945 7225 15979 7259
rect 24777 7225 24811 7259
rect 26424 7225 26458 7259
rect 2881 7157 2915 7191
rect 7205 7157 7239 7191
rect 12173 7157 12207 7191
rect 12909 7157 12943 7191
rect 13369 7157 13403 7191
rect 14841 7157 14875 7191
rect 14933 7157 14967 7191
rect 15577 7157 15611 7191
rect 16497 7157 16531 7191
rect 16589 7157 16623 7191
rect 18153 7157 18187 7191
rect 23949 7157 23983 7191
rect 1961 6953 1995 6987
rect 3341 6953 3375 6987
rect 6193 6953 6227 6987
rect 12633 6953 12667 6987
rect 13277 6953 13311 6987
rect 13737 6953 13771 6987
rect 14565 6953 14599 6987
rect 18981 6953 19015 6987
rect 19901 6953 19935 6987
rect 21281 6953 21315 6987
rect 22845 6953 22879 6987
rect 24133 6953 24167 6987
rect 24777 6953 24811 6987
rect 10057 6885 10091 6919
rect 21557 6885 21591 6919
rect 1409 6817 1443 6851
rect 4445 6817 4479 6851
rect 4537 6817 4571 6851
rect 6929 6817 6963 6851
rect 7389 6817 7423 6851
rect 12541 6817 12575 6851
rect 16589 6817 16623 6851
rect 16957 6817 16991 6851
rect 17417 6817 17451 6851
rect 19073 6817 19107 6851
rect 22937 6817 22971 6851
rect 24869 6817 24903 6851
rect 26525 6817 26559 6851
rect 4629 6749 4663 6783
rect 6285 6749 6319 6783
rect 6377 6749 6411 6783
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 12817 6749 12851 6783
rect 16129 6749 16163 6783
rect 17509 6749 17543 6783
rect 17601 6749 17635 6783
rect 18153 6749 18187 6783
rect 19165 6749 19199 6783
rect 23029 6749 23063 6783
rect 25053 6749 25087 6783
rect 1593 6681 1627 6715
rect 18613 6681 18647 6715
rect 22477 6681 22511 6715
rect 24409 6681 24443 6715
rect 26709 6681 26743 6715
rect 2421 6613 2455 6647
rect 4077 6613 4111 6647
rect 5181 6613 5215 6647
rect 5825 6613 5859 6647
rect 7297 6613 7331 6647
rect 8769 6613 8803 6647
rect 9689 6613 9723 6647
rect 12173 6613 12207 6647
rect 17049 6613 17083 6647
rect 20637 6613 20671 6647
rect 26249 6613 26283 6647
rect 2053 6409 2087 6443
rect 2329 6409 2363 6443
rect 6009 6409 6043 6443
rect 9045 6409 9079 6443
rect 9965 6409 9999 6443
rect 11069 6409 11103 6443
rect 12725 6409 12759 6443
rect 13093 6409 13127 6443
rect 17509 6409 17543 6443
rect 18061 6409 18095 6443
rect 19073 6409 19107 6443
rect 19441 6409 19475 6443
rect 20453 6409 20487 6443
rect 22569 6409 22603 6443
rect 22937 6409 22971 6443
rect 23213 6409 23247 6443
rect 24409 6409 24443 6443
rect 25237 6409 25271 6443
rect 26985 6409 27019 6443
rect 4997 6341 5031 6375
rect 9781 6341 9815 6375
rect 15761 6341 15795 6375
rect 17141 6341 17175 6375
rect 3709 6273 3743 6307
rect 3893 6273 3927 6307
rect 5457 6273 5491 6307
rect 5549 6273 5583 6307
rect 6653 6273 6687 6307
rect 7665 6273 7699 6307
rect 10517 6273 10551 6307
rect 12173 6273 12207 6307
rect 15393 6273 15427 6307
rect 16313 6273 16347 6307
rect 16497 6273 16531 6307
rect 18613 6273 18647 6307
rect 21097 6273 21131 6307
rect 26249 6273 26283 6307
rect 1409 6205 1443 6239
rect 2789 6205 2823 6239
rect 3617 6205 3651 6239
rect 7389 6205 7423 6239
rect 7481 6205 7515 6239
rect 17877 6205 17911 6239
rect 18429 6205 18463 6239
rect 21005 6205 21039 6239
rect 26433 6205 26467 6239
rect 3157 6137 3191 6171
rect 5365 6137 5399 6171
rect 9413 6137 9447 6171
rect 10425 6137 10459 6171
rect 15025 6137 15059 6171
rect 16221 6137 16255 6171
rect 1593 6069 1627 6103
rect 3249 6069 3283 6103
rect 4353 6069 4387 6103
rect 4721 6069 4755 6103
rect 7021 6069 7055 6103
rect 8033 6069 8067 6103
rect 10333 6069 10367 6103
rect 15853 6069 15887 6103
rect 18521 6069 18555 6103
rect 20545 6069 20579 6103
rect 20913 6069 20947 6103
rect 24777 6069 24811 6103
rect 26617 6069 26651 6103
rect 4353 5865 4387 5899
rect 5089 5865 5123 5899
rect 5457 5865 5491 5899
rect 5917 5865 5951 5899
rect 9965 5865 9999 5899
rect 10333 5865 10367 5899
rect 10609 5865 10643 5899
rect 11069 5865 11103 5899
rect 12173 5865 12207 5899
rect 12633 5865 12667 5899
rect 17233 5865 17267 5899
rect 18061 5865 18095 5899
rect 18613 5865 18647 5899
rect 19625 5865 19659 5899
rect 20637 5865 20671 5899
rect 20913 5865 20947 5899
rect 1768 5797 1802 5831
rect 6193 5797 6227 5831
rect 7389 5797 7423 5831
rect 12541 5797 12575 5831
rect 16120 5797 16154 5831
rect 1501 5729 1535 5763
rect 7481 5729 7515 5763
rect 10977 5729 11011 5763
rect 13645 5729 13679 5763
rect 15853 5729 15887 5763
rect 22641 5729 22675 5763
rect 26525 5729 26559 5763
rect 7665 5661 7699 5695
rect 11253 5661 11287 5695
rect 12817 5661 12851 5695
rect 19717 5661 19751 5695
rect 19809 5661 19843 5695
rect 22385 5661 22419 5695
rect 2881 5525 2915 5559
rect 7021 5525 7055 5559
rect 13369 5525 13403 5559
rect 19257 5525 19291 5559
rect 23765 5525 23799 5559
rect 25513 5525 25547 5559
rect 26709 5525 26743 5559
rect 1593 5321 1627 5355
rect 2789 5321 2823 5355
rect 3985 5321 4019 5355
rect 6653 5321 6687 5355
rect 7665 5321 7699 5355
rect 10793 5321 10827 5355
rect 12265 5321 12299 5355
rect 12633 5321 12667 5355
rect 14657 5321 14691 5355
rect 16037 5321 16071 5355
rect 17049 5321 17083 5355
rect 18981 5321 19015 5355
rect 19717 5321 19751 5355
rect 20545 5321 20579 5355
rect 27353 5321 27387 5355
rect 10701 5253 10735 5287
rect 15577 5253 15611 5287
rect 20085 5253 20119 5287
rect 22477 5253 22511 5287
rect 26801 5253 26835 5287
rect 2421 5185 2455 5219
rect 3341 5185 3375 5219
rect 3433 5185 3467 5219
rect 7113 5185 7147 5219
rect 10333 5185 10367 5219
rect 11437 5185 11471 5219
rect 13277 5185 13311 5219
rect 16681 5185 16715 5219
rect 20361 5185 20395 5219
rect 21189 5185 21223 5219
rect 1409 5117 1443 5151
rect 8125 5117 8159 5151
rect 15945 5117 15979 5151
rect 16405 5117 16439 5151
rect 20913 5117 20947 5151
rect 25421 5117 25455 5151
rect 3249 5049 3283 5083
rect 7941 5049 7975 5083
rect 8370 5049 8404 5083
rect 11161 5049 11195 5083
rect 13093 5049 13127 5083
rect 13544 5049 13578 5083
rect 17417 5049 17451 5083
rect 21005 5049 21039 5083
rect 25666 5049 25700 5083
rect 2053 4981 2087 5015
rect 2881 4981 2915 5015
rect 6193 4981 6227 5015
rect 9505 4981 9539 5015
rect 11253 4981 11287 5015
rect 11897 4981 11931 5015
rect 16497 4981 16531 5015
rect 19349 4981 19383 5015
rect 22753 4981 22787 5015
rect 25237 4981 25271 5015
rect 1593 4777 1627 4811
rect 3157 4777 3191 4811
rect 7573 4777 7607 4811
rect 8125 4777 8159 4811
rect 10517 4777 10551 4811
rect 11253 4777 11287 4811
rect 11437 4777 11471 4811
rect 11805 4777 11839 4811
rect 13001 4777 13035 4811
rect 13369 4777 13403 4811
rect 16129 4777 16163 4811
rect 19625 4777 19659 4811
rect 20545 4777 20579 4811
rect 10885 4709 10919 4743
rect 16488 4709 16522 4743
rect 1409 4641 1443 4675
rect 2053 4641 2087 4675
rect 2513 4641 2547 4675
rect 4896 4641 4930 4675
rect 7481 4641 7515 4675
rect 13461 4641 13495 4675
rect 16221 4641 16255 4675
rect 23581 4641 23615 4675
rect 23848 4641 23882 4675
rect 26525 4641 26559 4675
rect 2421 4573 2455 4607
rect 4629 4573 4663 4607
rect 7757 4573 7791 4607
rect 11897 4573 11931 4607
rect 12081 4573 12115 4607
rect 13645 4573 13679 4607
rect 19717 4573 19751 4607
rect 19901 4573 19935 4607
rect 24961 4505 24995 4539
rect 2697 4437 2731 4471
rect 6009 4437 6043 4471
rect 7113 4437 7147 4471
rect 17601 4437 17635 4471
rect 19257 4437 19291 4471
rect 21649 4437 21683 4471
rect 26709 4437 26743 4471
rect 2605 4233 2639 4267
rect 4169 4233 4203 4267
rect 4813 4233 4847 4267
rect 7205 4233 7239 4267
rect 7481 4233 7515 4267
rect 11529 4233 11563 4267
rect 12173 4233 12207 4267
rect 13461 4233 13495 4267
rect 13737 4233 13771 4267
rect 17049 4233 17083 4267
rect 19349 4233 19383 4267
rect 21097 4233 21131 4267
rect 24225 4233 24259 4267
rect 27169 4233 27203 4267
rect 5181 4165 5215 4199
rect 7849 4165 7883 4199
rect 11805 4165 11839 4199
rect 13093 4165 13127 4199
rect 15853 4165 15887 4199
rect 19993 4165 20027 4199
rect 5917 4097 5951 4131
rect 16405 4097 16439 4131
rect 16497 4097 16531 4131
rect 18981 4097 19015 4131
rect 20637 4097 20671 4131
rect 21373 4097 21407 4131
rect 22017 4097 22051 4131
rect 22109 4097 22143 4131
rect 26801 4097 26835 4131
rect 1409 4029 1443 4063
rect 2789 4029 2823 4063
rect 3045 4029 3079 4063
rect 5273 4029 5307 4063
rect 19901 4029 19935 4063
rect 21925 4029 21959 4063
rect 23857 4029 23891 4063
rect 26249 4029 26283 4063
rect 27353 4029 27387 4063
rect 27905 4029 27939 4063
rect 2053 3961 2087 3995
rect 15485 3961 15519 3995
rect 16313 3961 16347 3995
rect 20361 3961 20395 3995
rect 1593 3893 1627 3927
rect 5457 3893 5491 3927
rect 15945 3893 15979 3927
rect 20453 3893 20487 3927
rect 21557 3893 21591 3927
rect 26433 3893 26467 3927
rect 27537 3893 27571 3927
rect 1593 3689 1627 3723
rect 3065 3689 3099 3723
rect 4353 3689 4387 3723
rect 5457 3689 5491 3723
rect 6193 3689 6227 3723
rect 7389 3689 7423 3723
rect 12173 3689 12207 3723
rect 15945 3689 15979 3723
rect 19349 3689 19383 3723
rect 20085 3689 20119 3723
rect 20913 3689 20947 3723
rect 21281 3689 21315 3723
rect 3525 3621 3559 3655
rect 6469 3621 6503 3655
rect 16313 3621 16347 3655
rect 17478 3621 17512 3655
rect 20361 3621 20395 3655
rect 1409 3553 1443 3587
rect 2513 3553 2547 3587
rect 11060 3553 11094 3587
rect 17233 3553 17267 3587
rect 25329 3553 25363 3587
rect 26525 3553 26559 3587
rect 2053 3485 2087 3519
rect 5549 3485 5583 3519
rect 5733 3485 5767 3519
rect 7481 3485 7515 3519
rect 7573 3485 7607 3519
rect 10793 3485 10827 3519
rect 21373 3485 21407 3519
rect 21465 3485 21499 3519
rect 25513 3417 25547 3451
rect 2697 3349 2731 3383
rect 4905 3349 4939 3383
rect 5089 3349 5123 3383
rect 6929 3349 6963 3383
rect 7021 3349 7055 3383
rect 18613 3349 18647 3383
rect 26709 3349 26743 3383
rect 2605 3145 2639 3179
rect 3893 3145 3927 3179
rect 5181 3145 5215 3179
rect 10609 3145 10643 3179
rect 11161 3145 11195 3179
rect 13185 3145 13219 3179
rect 15209 3145 15243 3179
rect 16589 3145 16623 3179
rect 17509 3145 17543 3179
rect 17785 3145 17819 3179
rect 22109 3145 22143 3179
rect 24317 3145 24351 3179
rect 24685 3145 24719 3179
rect 27353 3145 27387 3179
rect 6561 3077 6595 3111
rect 7849 3077 7883 3111
rect 11529 3077 11563 3111
rect 21557 3077 21591 3111
rect 24961 3077 24995 3111
rect 4445 3009 4479 3043
rect 7389 3009 7423 3043
rect 9137 3009 9171 3043
rect 19993 3009 20027 3043
rect 25329 3009 25363 3043
rect 1409 2941 1443 2975
rect 2237 2941 2271 2975
rect 2697 2941 2731 2975
rect 3433 2941 3467 2975
rect 4261 2941 4295 2975
rect 5457 2941 5491 2975
rect 5733 2941 5767 2975
rect 7205 2941 7239 2975
rect 8585 2941 8619 2975
rect 9229 2941 9263 2975
rect 9496 2941 9530 2975
rect 12449 2941 12483 2975
rect 14381 2941 14415 2975
rect 16681 2941 16715 2975
rect 16957 2941 16991 2975
rect 18889 2941 18923 2975
rect 19625 2941 19659 2975
rect 20177 2941 20211 2975
rect 20433 2941 20467 2975
rect 23673 2941 23707 2975
rect 24777 2941 24811 2975
rect 26433 2941 26467 2975
rect 26985 2941 27019 2975
rect 27537 2941 27571 2975
rect 28089 2941 28123 2975
rect 1685 2873 1719 2907
rect 3801 2873 3835 2907
rect 4353 2873 4387 2907
rect 7297 2873 7331 2907
rect 8217 2873 8251 2907
rect 12725 2873 12759 2907
rect 14657 2873 14691 2907
rect 19165 2873 19199 2907
rect 2881 2805 2915 2839
rect 6193 2805 6227 2839
rect 6837 2805 6871 2839
rect 23857 2805 23891 2839
rect 26617 2805 26651 2839
rect 27721 2805 27755 2839
rect 2329 2601 2363 2635
rect 5181 2601 5215 2635
rect 6285 2601 6319 2635
rect 6561 2601 6595 2635
rect 6929 2601 6963 2635
rect 9229 2601 9263 2635
rect 13645 2601 13679 2635
rect 16405 2601 16439 2635
rect 18613 2601 18647 2635
rect 19441 2601 19475 2635
rect 19993 2601 20027 2635
rect 20545 2601 20579 2635
rect 20913 2601 20947 2635
rect 21373 2601 21407 2635
rect 5825 2533 5859 2567
rect 1409 2465 1443 2499
rect 1961 2465 1995 2499
rect 2513 2465 2547 2499
rect 3249 2465 3283 2499
rect 3893 2465 3927 2499
rect 4077 2465 4111 2499
rect 5549 2465 5583 2499
rect 18981 2533 19015 2567
rect 19901 2533 19935 2567
rect 7297 2465 7331 2499
rect 7941 2465 7975 2499
rect 9781 2465 9815 2499
rect 10517 2465 10551 2499
rect 11069 2465 11103 2499
rect 11805 2465 11839 2499
rect 12817 2465 12851 2499
rect 15669 2465 15703 2499
rect 16957 2465 16991 2499
rect 17785 2465 17819 2499
rect 22293 2465 22327 2499
rect 23029 2465 23063 2499
rect 24041 2465 24075 2499
rect 24777 2465 24811 2499
rect 25697 2465 25731 2499
rect 26249 2465 26283 2499
rect 2789 2397 2823 2431
rect 4353 2397 4387 2431
rect 6561 2397 6595 2431
rect 7389 2397 7423 2431
rect 7481 2397 7515 2431
rect 9965 2397 9999 2431
rect 11253 2397 11287 2431
rect 13093 2397 13127 2431
rect 15945 2397 15979 2431
rect 17233 2397 17267 2431
rect 20085 2397 20119 2431
rect 22569 2397 22603 2431
rect 24225 2397 24259 2431
rect 6745 2329 6779 2363
rect 19533 2329 19567 2363
rect 1593 2261 1627 2295
rect 25881 2261 25915 2295
rect 27077 2261 27111 2295
<< metal1 >>
rect 3326 22108 3332 22160
rect 3384 22148 3390 22160
rect 12066 22148 12072 22160
rect 3384 22120 12072 22148
rect 3384 22108 3390 22120
rect 12066 22108 12072 22120
rect 12124 22108 12130 22160
rect 21818 22108 21824 22160
rect 21876 22148 21882 22160
rect 24854 22148 24860 22160
rect 21876 22120 24860 22148
rect 21876 22108 21882 22120
rect 24854 22108 24860 22120
rect 24912 22108 24918 22160
rect 1670 22040 1676 22092
rect 1728 22080 1734 22092
rect 2130 22080 2136 22092
rect 1728 22052 2136 22080
rect 1728 22040 1734 22052
rect 2130 22040 2136 22052
rect 2188 22040 2194 22092
rect 1104 21786 28888 21808
rect 1104 21734 5982 21786
rect 6034 21734 6046 21786
rect 6098 21734 6110 21786
rect 6162 21734 6174 21786
rect 6226 21734 15982 21786
rect 16034 21734 16046 21786
rect 16098 21734 16110 21786
rect 16162 21734 16174 21786
rect 16226 21734 25982 21786
rect 26034 21734 26046 21786
rect 26098 21734 26110 21786
rect 26162 21734 26174 21786
rect 26226 21734 28888 21786
rect 1104 21712 28888 21734
rect 1104 21242 28888 21264
rect 1104 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 20982 21242
rect 21034 21190 21046 21242
rect 21098 21190 21110 21242
rect 21162 21190 21174 21242
rect 21226 21190 28888 21242
rect 1104 21168 28888 21190
rect 3970 21088 3976 21140
rect 4028 21128 4034 21140
rect 7282 21128 7288 21140
rect 4028 21100 7288 21128
rect 4028 21088 4034 21100
rect 7282 21088 7288 21100
rect 7340 21088 7346 21140
rect 17034 20924 17040 20936
rect 16995 20896 17040 20924
rect 17034 20884 17040 20896
rect 17092 20884 17098 20936
rect 4062 20748 4068 20800
rect 4120 20788 4126 20800
rect 7558 20788 7564 20800
rect 4120 20760 7564 20788
rect 4120 20748 4126 20760
rect 7558 20748 7564 20760
rect 7616 20748 7622 20800
rect 8386 20788 8392 20800
rect 8347 20760 8392 20788
rect 8386 20748 8392 20760
rect 8444 20748 8450 20800
rect 13538 20788 13544 20800
rect 13499 20760 13544 20788
rect 13538 20748 13544 20760
rect 13596 20748 13602 20800
rect 23658 20788 23664 20800
rect 23619 20760 23664 20788
rect 23658 20748 23664 20760
rect 23716 20748 23722 20800
rect 1104 20698 28888 20720
rect 1104 20646 5982 20698
rect 6034 20646 6046 20698
rect 6098 20646 6110 20698
rect 6162 20646 6174 20698
rect 6226 20646 15982 20698
rect 16034 20646 16046 20698
rect 16098 20646 16110 20698
rect 16162 20646 16174 20698
rect 16226 20646 25982 20698
rect 26034 20646 26046 20698
rect 26098 20646 26110 20698
rect 26162 20646 26174 20698
rect 26226 20646 28888 20698
rect 1104 20624 28888 20646
rect 7101 20587 7159 20593
rect 7101 20553 7113 20587
rect 7147 20584 7159 20587
rect 8202 20584 8208 20596
rect 7147 20556 8208 20584
rect 7147 20553 7159 20556
rect 7101 20547 7159 20553
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 21634 20544 21640 20596
rect 21692 20584 21698 20596
rect 21913 20587 21971 20593
rect 21913 20584 21925 20587
rect 21692 20556 21925 20584
rect 21692 20544 21698 20556
rect 21913 20553 21925 20556
rect 21959 20553 21971 20587
rect 21913 20547 21971 20553
rect 20622 20516 20628 20528
rect 20583 20488 20628 20516
rect 20622 20476 20628 20488
rect 20680 20476 20686 20528
rect 16945 20451 17003 20457
rect 16945 20417 16957 20451
rect 16991 20448 17003 20451
rect 18322 20448 18328 20460
rect 16991 20420 18328 20448
rect 16991 20417 17003 20420
rect 16945 20411 17003 20417
rect 18322 20408 18328 20420
rect 18380 20408 18386 20460
rect 3510 20380 3516 20392
rect 3471 20352 3516 20380
rect 3510 20340 3516 20352
rect 3568 20340 3574 20392
rect 8297 20383 8355 20389
rect 8297 20349 8309 20383
rect 8343 20380 8355 20383
rect 8386 20380 8392 20392
rect 8343 20352 8392 20380
rect 8343 20349 8355 20352
rect 8297 20343 8355 20349
rect 8386 20340 8392 20352
rect 8444 20340 8450 20392
rect 12434 20340 12440 20392
rect 12492 20380 12498 20392
rect 13538 20380 13544 20392
rect 12492 20352 13544 20380
rect 12492 20340 12498 20352
rect 13538 20340 13544 20352
rect 13596 20340 13602 20392
rect 16666 20380 16672 20392
rect 16627 20352 16672 20380
rect 16666 20340 16672 20352
rect 16724 20380 16730 20392
rect 17405 20383 17463 20389
rect 17405 20380 17417 20383
rect 16724 20352 17417 20380
rect 16724 20340 16730 20352
rect 17405 20349 17417 20352
rect 17451 20349 17463 20383
rect 19242 20380 19248 20392
rect 19203 20352 19248 20380
rect 17405 20343 17463 20349
rect 19242 20340 19248 20352
rect 19300 20340 19306 20392
rect 20640 20380 20668 20476
rect 21729 20383 21787 20389
rect 21729 20380 21741 20383
rect 20640 20352 21741 20380
rect 21729 20349 21741 20352
rect 21775 20380 21787 20383
rect 22281 20383 22339 20389
rect 22281 20380 22293 20383
rect 21775 20352 22293 20380
rect 21775 20349 21787 20352
rect 21729 20343 21787 20349
rect 22281 20349 22293 20352
rect 22327 20349 22339 20383
rect 23658 20380 23664 20392
rect 23619 20352 23664 20380
rect 22281 20343 22339 20349
rect 23658 20340 23664 20352
rect 23716 20340 23722 20392
rect 26145 20383 26203 20389
rect 26145 20349 26157 20383
rect 26191 20380 26203 20383
rect 26191 20352 26832 20380
rect 26191 20349 26203 20352
rect 26145 20343 26203 20349
rect 3421 20315 3479 20321
rect 3421 20281 3433 20315
rect 3467 20312 3479 20315
rect 3758 20315 3816 20321
rect 3758 20312 3770 20315
rect 3467 20284 3770 20312
rect 3467 20281 3479 20284
rect 3421 20275 3479 20281
rect 3758 20281 3770 20284
rect 3804 20312 3816 20315
rect 4062 20312 4068 20324
rect 3804 20284 4068 20312
rect 3804 20281 3816 20284
rect 3758 20275 3816 20281
rect 4062 20272 4068 20284
rect 4120 20272 4126 20324
rect 8542 20315 8600 20321
rect 8542 20312 8554 20315
rect 8128 20284 8554 20312
rect 4890 20244 4896 20256
rect 4851 20216 4896 20244
rect 4890 20204 4896 20216
rect 4948 20204 4954 20256
rect 7834 20204 7840 20256
rect 7892 20244 7898 20256
rect 8128 20253 8156 20284
rect 8542 20281 8554 20284
rect 8588 20281 8600 20315
rect 13786 20315 13844 20321
rect 13786 20312 13798 20315
rect 8542 20275 8600 20281
rect 13464 20284 13798 20312
rect 13464 20256 13492 20284
rect 13786 20281 13798 20284
rect 13832 20281 13844 20315
rect 13786 20275 13844 20281
rect 19153 20315 19211 20321
rect 19153 20281 19165 20315
rect 19199 20312 19211 20315
rect 19490 20315 19548 20321
rect 19490 20312 19502 20315
rect 19199 20284 19502 20312
rect 19199 20281 19211 20284
rect 19153 20275 19211 20281
rect 19490 20281 19502 20284
rect 19536 20312 19548 20315
rect 20714 20312 20720 20324
rect 19536 20284 20720 20312
rect 19536 20281 19548 20284
rect 19490 20275 19548 20281
rect 20714 20272 20720 20284
rect 20772 20272 20778 20324
rect 23477 20315 23535 20321
rect 23477 20281 23489 20315
rect 23523 20312 23535 20315
rect 23928 20315 23986 20321
rect 23928 20312 23940 20315
rect 23523 20284 23940 20312
rect 23523 20281 23535 20284
rect 23477 20275 23535 20281
rect 23928 20281 23940 20284
rect 23974 20312 23986 20315
rect 24670 20312 24676 20324
rect 23974 20284 24676 20312
rect 23974 20281 23986 20284
rect 23928 20275 23986 20281
rect 24670 20272 24676 20284
rect 24728 20272 24734 20324
rect 8113 20247 8171 20253
rect 8113 20244 8125 20247
rect 7892 20216 8125 20244
rect 7892 20204 7898 20216
rect 8113 20213 8125 20216
rect 8159 20213 8171 20247
rect 9674 20244 9680 20256
rect 9635 20216 9680 20244
rect 8113 20207 8171 20213
rect 9674 20204 9680 20216
rect 9732 20204 9738 20256
rect 13446 20244 13452 20256
rect 13407 20216 13452 20244
rect 13446 20204 13452 20216
rect 13504 20204 13510 20256
rect 14921 20247 14979 20253
rect 14921 20213 14933 20247
rect 14967 20244 14979 20247
rect 15102 20244 15108 20256
rect 14967 20216 15108 20244
rect 14967 20213 14979 20216
rect 14921 20207 14979 20213
rect 15102 20204 15108 20216
rect 15160 20204 15166 20256
rect 25038 20244 25044 20256
rect 24999 20216 25044 20244
rect 25038 20204 25044 20216
rect 25096 20204 25102 20256
rect 26326 20244 26332 20256
rect 26287 20216 26332 20244
rect 26326 20204 26332 20216
rect 26384 20204 26390 20256
rect 26804 20253 26832 20352
rect 26789 20247 26847 20253
rect 26789 20213 26801 20247
rect 26835 20244 26847 20247
rect 26878 20244 26884 20256
rect 26835 20216 26884 20244
rect 26835 20213 26847 20216
rect 26789 20207 26847 20213
rect 26878 20204 26884 20216
rect 26936 20204 26942 20256
rect 1104 20154 28888 20176
rect 1104 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 20982 20154
rect 21034 20102 21046 20154
rect 21098 20102 21110 20154
rect 21162 20102 21174 20154
rect 21226 20102 28888 20154
rect 1104 20080 28888 20102
rect 3510 20040 3516 20052
rect 3471 20012 3516 20040
rect 3510 20000 3516 20012
rect 3568 20000 3574 20052
rect 6638 20040 6644 20052
rect 6599 20012 6644 20040
rect 6638 20000 6644 20012
rect 6696 20000 6702 20052
rect 13078 20000 13084 20052
rect 13136 20040 13142 20052
rect 13725 20043 13783 20049
rect 13725 20040 13737 20043
rect 13136 20012 13737 20040
rect 13136 20000 13142 20012
rect 13725 20009 13737 20012
rect 13771 20040 13783 20043
rect 15749 20043 15807 20049
rect 15749 20040 15761 20043
rect 13771 20012 15761 20040
rect 13771 20009 13783 20012
rect 13725 20003 13783 20009
rect 15749 20009 15761 20012
rect 15795 20009 15807 20043
rect 15749 20003 15807 20009
rect 17034 20000 17040 20052
rect 17092 20040 17098 20052
rect 17678 20040 17684 20052
rect 17092 20012 17684 20040
rect 17092 20000 17098 20012
rect 17678 20000 17684 20012
rect 17736 20000 17742 20052
rect 19242 20040 19248 20052
rect 19203 20012 19248 20040
rect 19242 20000 19248 20012
rect 19300 20000 19306 20052
rect 26697 20043 26755 20049
rect 26697 20009 26709 20043
rect 26743 20040 26755 20043
rect 28258 20040 28264 20052
rect 26743 20012 28264 20040
rect 26743 20009 26755 20012
rect 26697 20003 26755 20009
rect 28258 20000 28264 20012
rect 28316 20000 28322 20052
rect 3528 19904 3556 20000
rect 6656 19972 6684 20000
rect 8018 19972 8024 19984
rect 6656 19944 8024 19972
rect 8018 19932 8024 19944
rect 8076 19972 8082 19984
rect 8076 19944 8248 19972
rect 8076 19932 8082 19944
rect 5258 19904 5264 19916
rect 3528 19876 5264 19904
rect 5258 19864 5264 19876
rect 5316 19864 5322 19916
rect 5534 19913 5540 19916
rect 5528 19904 5540 19913
rect 5447 19876 5540 19904
rect 5528 19867 5540 19876
rect 5592 19904 5598 19916
rect 6730 19904 6736 19916
rect 5592 19876 6736 19904
rect 5534 19864 5540 19867
rect 5592 19864 5598 19876
rect 6730 19864 6736 19876
rect 6788 19864 6794 19916
rect 8113 19907 8171 19913
rect 8113 19904 8125 19907
rect 7576 19876 8125 19904
rect 6914 19728 6920 19780
rect 6972 19768 6978 19780
rect 7576 19777 7604 19876
rect 8113 19873 8125 19876
rect 8159 19873 8171 19907
rect 8220 19904 8248 19944
rect 10704 19944 10916 19972
rect 10704 19916 10732 19944
rect 8220 19876 8340 19904
rect 8113 19867 8171 19873
rect 8202 19836 8208 19848
rect 8163 19808 8208 19836
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 8312 19845 8340 19876
rect 8386 19864 8392 19916
rect 8444 19904 8450 19916
rect 10686 19904 10692 19916
rect 8444 19876 10692 19904
rect 8444 19864 8450 19876
rect 10686 19864 10692 19876
rect 10744 19864 10750 19916
rect 10788 19907 10846 19913
rect 10788 19873 10800 19907
rect 10834 19904 10846 19907
rect 10888 19904 10916 19944
rect 10962 19932 10968 19984
rect 11020 19932 11026 19984
rect 17310 19932 17316 19984
rect 17368 19972 17374 19984
rect 17773 19975 17831 19981
rect 17773 19972 17785 19975
rect 17368 19944 17785 19972
rect 17368 19932 17374 19944
rect 17773 19941 17785 19944
rect 17819 19941 17831 19975
rect 17773 19935 17831 19941
rect 21542 19932 21548 19984
rect 21600 19972 21606 19984
rect 21790 19975 21848 19981
rect 21790 19972 21802 19975
rect 21600 19944 21802 19972
rect 21600 19932 21606 19944
rect 21790 19941 21802 19944
rect 21836 19941 21848 19975
rect 21790 19935 21848 19941
rect 10834 19876 10916 19904
rect 10980 19904 11008 19932
rect 11048 19907 11106 19913
rect 11048 19904 11060 19907
rect 10980 19876 11060 19904
rect 10834 19873 10846 19876
rect 10788 19867 10846 19873
rect 11048 19873 11060 19876
rect 11094 19904 11106 19907
rect 11606 19904 11612 19916
rect 11094 19876 11612 19904
rect 11094 19873 11106 19876
rect 11048 19867 11106 19873
rect 11606 19864 11612 19876
rect 11664 19864 11670 19916
rect 16117 19907 16175 19913
rect 16117 19873 16129 19907
rect 16163 19904 16175 19907
rect 16390 19904 16396 19916
rect 16163 19876 16396 19904
rect 16163 19873 16175 19876
rect 16117 19867 16175 19873
rect 16390 19864 16396 19876
rect 16448 19904 16454 19916
rect 16448 19876 17356 19904
rect 16448 19864 16454 19876
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19805 8355 19839
rect 13817 19839 13875 19845
rect 13817 19836 13829 19839
rect 8297 19799 8355 19805
rect 13740 19808 13829 19836
rect 13740 19780 13768 19808
rect 13817 19805 13829 19808
rect 13863 19805 13875 19839
rect 13998 19836 14004 19848
rect 13911 19808 14004 19836
rect 13817 19799 13875 19805
rect 13998 19796 14004 19808
rect 14056 19836 14062 19848
rect 15102 19836 15108 19848
rect 14056 19808 15108 19836
rect 14056 19796 14062 19808
rect 15102 19796 15108 19808
rect 15160 19796 15166 19848
rect 15838 19796 15844 19848
rect 15896 19836 15902 19848
rect 16209 19839 16267 19845
rect 16209 19836 16221 19839
rect 15896 19808 16221 19836
rect 15896 19796 15902 19808
rect 16209 19805 16221 19808
rect 16255 19805 16267 19839
rect 16209 19799 16267 19805
rect 16298 19796 16304 19848
rect 16356 19836 16362 19848
rect 16356 19808 16401 19836
rect 16356 19796 16362 19808
rect 7561 19771 7619 19777
rect 7561 19768 7573 19771
rect 6972 19740 7573 19768
rect 6972 19728 6978 19740
rect 7561 19737 7573 19740
rect 7607 19737 7619 19771
rect 7742 19768 7748 19780
rect 7703 19740 7748 19768
rect 7561 19731 7619 19737
rect 7742 19728 7748 19740
rect 7800 19728 7806 19780
rect 13722 19728 13728 19780
rect 13780 19728 13786 19780
rect 17328 19777 17356 19876
rect 21634 19864 21640 19916
rect 21692 19864 21698 19916
rect 26513 19907 26571 19913
rect 26513 19873 26525 19907
rect 26559 19904 26571 19907
rect 26786 19904 26792 19916
rect 26559 19876 26792 19904
rect 26559 19873 26571 19876
rect 26513 19867 26571 19873
rect 26786 19864 26792 19876
rect 26844 19864 26850 19916
rect 17862 19836 17868 19848
rect 17823 19808 17868 19836
rect 17862 19796 17868 19808
rect 17920 19796 17926 19848
rect 21545 19839 21603 19845
rect 21545 19805 21557 19839
rect 21591 19836 21603 19839
rect 21652 19836 21680 19864
rect 21591 19808 21680 19836
rect 21591 19805 21603 19808
rect 21545 19799 21603 19805
rect 17313 19771 17371 19777
rect 17313 19737 17325 19771
rect 17359 19737 17371 19771
rect 17313 19731 17371 19737
rect 3142 19700 3148 19712
rect 3103 19672 3148 19700
rect 3142 19660 3148 19672
rect 3200 19660 3206 19712
rect 7190 19700 7196 19712
rect 7151 19672 7196 19700
rect 7190 19660 7196 19672
rect 7248 19660 7254 19712
rect 8846 19700 8852 19712
rect 8807 19672 8852 19700
rect 8846 19660 8852 19672
rect 8904 19660 8910 19712
rect 11422 19660 11428 19712
rect 11480 19700 11486 19712
rect 12161 19703 12219 19709
rect 12161 19700 12173 19703
rect 11480 19672 12173 19700
rect 11480 19660 11486 19672
rect 12161 19669 12173 19672
rect 12207 19669 12219 19703
rect 12161 19663 12219 19669
rect 13170 19660 13176 19712
rect 13228 19700 13234 19712
rect 13357 19703 13415 19709
rect 13357 19700 13369 19703
rect 13228 19672 13369 19700
rect 13228 19660 13234 19672
rect 13357 19669 13369 19672
rect 13403 19669 13415 19703
rect 13357 19663 13415 19669
rect 14461 19703 14519 19709
rect 14461 19669 14473 19703
rect 14507 19700 14519 19703
rect 15102 19700 15108 19712
rect 14507 19672 15108 19700
rect 14507 19669 14519 19672
rect 14461 19663 14519 19669
rect 15102 19660 15108 19672
rect 15160 19660 15166 19712
rect 22922 19700 22928 19712
rect 22883 19672 22928 19700
rect 22922 19660 22928 19672
rect 22980 19660 22986 19712
rect 23750 19700 23756 19712
rect 23711 19672 23756 19700
rect 23750 19660 23756 19672
rect 23808 19660 23814 19712
rect 25317 19703 25375 19709
rect 25317 19669 25329 19703
rect 25363 19700 25375 19703
rect 25590 19700 25596 19712
rect 25363 19672 25596 19700
rect 25363 19669 25375 19672
rect 25317 19663 25375 19669
rect 25590 19660 25596 19672
rect 25648 19660 25654 19712
rect 1104 19610 28888 19632
rect 1104 19558 5982 19610
rect 6034 19558 6046 19610
rect 6098 19558 6110 19610
rect 6162 19558 6174 19610
rect 6226 19558 15982 19610
rect 16034 19558 16046 19610
rect 16098 19558 16110 19610
rect 16162 19558 16174 19610
rect 16226 19558 25982 19610
rect 26034 19558 26046 19610
rect 26098 19558 26110 19610
rect 26162 19558 26174 19610
rect 26226 19558 28888 19610
rect 1104 19536 28888 19558
rect 5258 19456 5264 19508
rect 5316 19496 5322 19508
rect 5629 19499 5687 19505
rect 5629 19496 5641 19499
rect 5316 19468 5641 19496
rect 5316 19456 5322 19468
rect 5629 19465 5641 19468
rect 5675 19465 5687 19499
rect 5629 19459 5687 19465
rect 8018 19456 8024 19508
rect 8076 19496 8082 19508
rect 8113 19499 8171 19505
rect 8113 19496 8125 19499
rect 8076 19468 8125 19496
rect 8076 19456 8082 19468
rect 8113 19465 8125 19468
rect 8159 19465 8171 19499
rect 13078 19496 13084 19508
rect 13039 19468 13084 19496
rect 8113 19459 8171 19465
rect 13078 19456 13084 19468
rect 13136 19456 13142 19508
rect 13722 19496 13728 19508
rect 13683 19468 13728 19496
rect 13722 19456 13728 19468
rect 13780 19456 13786 19508
rect 17678 19496 17684 19508
rect 17639 19468 17684 19496
rect 17678 19456 17684 19468
rect 17736 19456 17742 19508
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 21177 19499 21235 19505
rect 21177 19496 21189 19499
rect 20864 19468 21189 19496
rect 20864 19456 20870 19468
rect 21177 19465 21189 19468
rect 21223 19496 21235 19499
rect 21634 19496 21640 19508
rect 21223 19468 21640 19496
rect 21223 19465 21235 19468
rect 21177 19459 21235 19465
rect 21634 19456 21640 19468
rect 21692 19456 21698 19508
rect 23474 19496 23480 19508
rect 23387 19468 23480 19496
rect 23474 19456 23480 19468
rect 23532 19496 23538 19508
rect 23532 19468 24348 19496
rect 23532 19456 23538 19468
rect 2593 19431 2651 19437
rect 2593 19397 2605 19431
rect 2639 19428 2651 19431
rect 13449 19431 13507 19437
rect 2639 19400 3740 19428
rect 2639 19397 2651 19400
rect 2593 19391 2651 19397
rect 3712 19372 3740 19400
rect 13449 19397 13461 19431
rect 13495 19428 13507 19431
rect 13998 19428 14004 19440
rect 13495 19400 14004 19428
rect 13495 19397 13507 19400
rect 13449 19391 13507 19397
rect 13998 19388 14004 19400
rect 14056 19388 14062 19440
rect 17037 19431 17095 19437
rect 17037 19397 17049 19431
rect 17083 19428 17095 19431
rect 17126 19428 17132 19440
rect 17083 19400 17132 19428
rect 17083 19397 17095 19400
rect 17037 19391 17095 19397
rect 17126 19388 17132 19400
rect 17184 19428 17190 19440
rect 17862 19428 17868 19440
rect 17184 19400 17868 19428
rect 17184 19388 17190 19400
rect 17862 19388 17868 19400
rect 17920 19388 17926 19440
rect 23661 19431 23719 19437
rect 23661 19397 23673 19431
rect 23707 19397 23719 19431
rect 23661 19391 23719 19397
rect 3694 19360 3700 19372
rect 3655 19332 3700 19360
rect 3694 19320 3700 19332
rect 3752 19320 3758 19372
rect 5534 19360 5540 19372
rect 5460 19332 5540 19360
rect 3142 19252 3148 19304
rect 3200 19292 3206 19304
rect 3421 19295 3479 19301
rect 3421 19292 3433 19295
rect 3200 19264 3433 19292
rect 3200 19252 3206 19264
rect 3421 19261 3433 19264
rect 3467 19292 3479 19295
rect 4617 19295 4675 19301
rect 4617 19292 4629 19295
rect 3467 19264 4629 19292
rect 3467 19261 3479 19264
rect 3421 19255 3479 19261
rect 4617 19261 4629 19264
rect 4663 19261 4675 19295
rect 4617 19255 4675 19261
rect 5353 19295 5411 19301
rect 5353 19261 5365 19295
rect 5399 19292 5411 19295
rect 5460 19292 5488 19332
rect 5534 19320 5540 19332
rect 5592 19320 5598 19372
rect 7742 19360 7748 19372
rect 7703 19332 7748 19360
rect 7742 19320 7748 19332
rect 7800 19320 7806 19372
rect 8754 19360 8760 19372
rect 8667 19332 8760 19360
rect 8754 19320 8760 19332
rect 8812 19360 8818 19372
rect 9493 19363 9551 19369
rect 9493 19360 9505 19363
rect 8812 19332 9505 19360
rect 8812 19320 8818 19332
rect 9493 19329 9505 19332
rect 9539 19360 9551 19363
rect 9674 19360 9680 19372
rect 9539 19332 9680 19360
rect 9539 19329 9551 19332
rect 9493 19323 9551 19329
rect 9674 19320 9680 19332
rect 9732 19320 9738 19372
rect 11790 19320 11796 19372
rect 11848 19360 11854 19372
rect 13906 19360 13912 19372
rect 11848 19332 13912 19360
rect 11848 19320 11854 19332
rect 13906 19320 13912 19332
rect 13964 19320 13970 19372
rect 22649 19363 22707 19369
rect 22649 19360 22661 19363
rect 22112 19332 22661 19360
rect 5399 19264 5488 19292
rect 6273 19295 6331 19301
rect 5399 19261 5411 19264
rect 5353 19255 5411 19261
rect 6273 19261 6285 19295
rect 6319 19292 6331 19295
rect 7760 19292 7788 19320
rect 6319 19264 7788 19292
rect 6319 19261 6331 19264
rect 6273 19255 6331 19261
rect 8386 19252 8392 19304
rect 8444 19292 8450 19304
rect 8846 19292 8852 19304
rect 8444 19264 8852 19292
rect 8444 19252 8450 19264
rect 8846 19252 8852 19264
rect 8904 19292 8910 19304
rect 9217 19295 9275 19301
rect 9217 19292 9229 19295
rect 8904 19264 9229 19292
rect 8904 19252 8910 19264
rect 9217 19261 9229 19264
rect 9263 19261 9275 19295
rect 9217 19255 9275 19261
rect 10873 19295 10931 19301
rect 10873 19261 10885 19295
rect 10919 19292 10931 19295
rect 10962 19292 10968 19304
rect 10919 19264 10968 19292
rect 10919 19261 10931 19264
rect 10873 19255 10931 19261
rect 10962 19252 10968 19264
rect 11020 19252 11026 19304
rect 14369 19295 14427 19301
rect 14369 19261 14381 19295
rect 14415 19292 14427 19295
rect 15102 19292 15108 19304
rect 14415 19264 15108 19292
rect 14415 19261 14427 19264
rect 14369 19255 14427 19261
rect 15102 19252 15108 19264
rect 15160 19252 15166 19304
rect 20714 19252 20720 19304
rect 20772 19292 20778 19304
rect 21821 19295 21879 19301
rect 21821 19292 21833 19295
rect 20772 19264 21833 19292
rect 20772 19252 20778 19264
rect 21821 19261 21833 19264
rect 21867 19292 21879 19295
rect 22112 19292 22140 19332
rect 22649 19329 22661 19332
rect 22695 19360 22707 19363
rect 22922 19360 22928 19372
rect 22695 19332 22928 19360
rect 22695 19329 22707 19332
rect 22649 19323 22707 19329
rect 22922 19320 22928 19332
rect 22980 19320 22986 19372
rect 21867 19264 22140 19292
rect 22373 19295 22431 19301
rect 21867 19261 21879 19264
rect 21821 19255 21879 19261
rect 22373 19261 22385 19295
rect 22419 19292 22431 19295
rect 22462 19292 22468 19304
rect 22419 19264 22468 19292
rect 22419 19261 22431 19264
rect 22373 19255 22431 19261
rect 22462 19252 22468 19264
rect 22520 19292 22526 19304
rect 23676 19292 23704 19391
rect 23750 19320 23756 19372
rect 23808 19360 23814 19372
rect 24320 19369 24348 19468
rect 24670 19388 24676 19440
rect 24728 19428 24734 19440
rect 24765 19431 24823 19437
rect 24765 19428 24777 19431
rect 24728 19400 24777 19428
rect 24728 19388 24734 19400
rect 24765 19397 24777 19400
rect 24811 19428 24823 19431
rect 24811 19400 25912 19428
rect 24811 19397 24823 19400
rect 24765 19391 24823 19397
rect 24121 19363 24179 19369
rect 24121 19360 24133 19363
rect 23808 19332 24133 19360
rect 23808 19320 23814 19332
rect 24121 19329 24133 19332
rect 24167 19329 24179 19363
rect 24121 19323 24179 19329
rect 24305 19363 24363 19369
rect 24305 19329 24317 19363
rect 24351 19360 24363 19363
rect 25038 19360 25044 19372
rect 24351 19332 25044 19360
rect 24351 19329 24363 19332
rect 24305 19323 24363 19329
rect 25038 19320 25044 19332
rect 25096 19320 25102 19372
rect 25884 19369 25912 19400
rect 25869 19363 25927 19369
rect 25869 19329 25881 19363
rect 25915 19360 25927 19363
rect 26142 19360 26148 19372
rect 25915 19332 26148 19360
rect 25915 19329 25927 19332
rect 25869 19323 25927 19329
rect 26142 19320 26148 19332
rect 26200 19320 26206 19372
rect 22520 19264 23704 19292
rect 22520 19252 22526 19264
rect 24854 19252 24860 19304
rect 24912 19292 24918 19304
rect 25133 19295 25191 19301
rect 25133 19292 25145 19295
rect 24912 19264 25145 19292
rect 24912 19252 24918 19264
rect 25133 19261 25145 19264
rect 25179 19292 25191 19295
rect 25590 19292 25596 19304
rect 25179 19264 25360 19292
rect 25551 19264 25596 19292
rect 25179 19261 25191 19264
rect 25133 19255 25191 19261
rect 2961 19227 3019 19233
rect 2961 19193 2973 19227
rect 3007 19224 3019 19227
rect 7561 19227 7619 19233
rect 7561 19224 7573 19227
rect 3007 19196 3556 19224
rect 3007 19193 3019 19196
rect 2961 19187 3019 19193
rect 3050 19156 3056 19168
rect 3011 19128 3056 19156
rect 3050 19116 3056 19128
rect 3108 19116 3114 19168
rect 3528 19165 3556 19196
rect 6564 19196 7573 19224
rect 6564 19168 6592 19196
rect 7561 19193 7573 19196
rect 7607 19224 7619 19227
rect 8110 19224 8116 19236
rect 7607 19196 8116 19224
rect 7607 19193 7619 19196
rect 7561 19187 7619 19193
rect 8110 19184 8116 19196
rect 8168 19184 8174 19236
rect 8294 19184 8300 19236
rect 8352 19224 8358 19236
rect 14185 19227 14243 19233
rect 8352 19196 8892 19224
rect 8352 19184 8358 19196
rect 3513 19159 3571 19165
rect 3513 19125 3525 19159
rect 3559 19156 3571 19159
rect 3602 19156 3608 19168
rect 3559 19128 3608 19156
rect 3559 19125 3571 19128
rect 3513 19119 3571 19125
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 6546 19156 6552 19168
rect 6507 19128 6552 19156
rect 6546 19116 6552 19128
rect 6604 19116 6610 19168
rect 7098 19156 7104 19168
rect 7059 19128 7104 19156
rect 7098 19116 7104 19128
rect 7156 19116 7162 19168
rect 7190 19116 7196 19168
rect 7248 19156 7254 19168
rect 8864 19165 8892 19196
rect 14185 19193 14197 19227
rect 14231 19224 14243 19227
rect 14636 19227 14694 19233
rect 14636 19224 14648 19227
rect 14231 19196 14648 19224
rect 14231 19193 14243 19196
rect 14185 19187 14243 19193
rect 14636 19193 14648 19196
rect 14682 19224 14694 19227
rect 14734 19224 14740 19236
rect 14682 19196 14740 19224
rect 14682 19193 14694 19196
rect 14636 19187 14694 19193
rect 14734 19184 14740 19196
rect 14792 19184 14798 19236
rect 23109 19227 23167 19233
rect 23109 19193 23121 19227
rect 23155 19224 23167 19227
rect 24029 19227 24087 19233
rect 24029 19224 24041 19227
rect 23155 19196 24041 19224
rect 23155 19193 23167 19196
rect 23109 19187 23167 19193
rect 24029 19193 24041 19196
rect 24075 19224 24087 19227
rect 25332 19224 25360 19264
rect 25590 19252 25596 19264
rect 25648 19292 25654 19304
rect 26789 19295 26847 19301
rect 26789 19292 26801 19295
rect 25648 19264 26801 19292
rect 25648 19252 25654 19264
rect 26789 19261 26801 19264
rect 26835 19261 26847 19295
rect 26789 19255 26847 19261
rect 25685 19227 25743 19233
rect 25685 19224 25697 19227
rect 24075 19196 25268 19224
rect 25332 19196 25697 19224
rect 24075 19193 24087 19196
rect 24029 19187 24087 19193
rect 7469 19159 7527 19165
rect 7469 19156 7481 19159
rect 7248 19128 7481 19156
rect 7248 19116 7254 19128
rect 7469 19125 7481 19128
rect 7515 19125 7527 19159
rect 7469 19119 7527 19125
rect 8849 19159 8907 19165
rect 8849 19125 8861 19159
rect 8895 19125 8907 19159
rect 8849 19119 8907 19125
rect 9306 19116 9312 19168
rect 9364 19156 9370 19168
rect 9364 19128 9409 19156
rect 9364 19116 9370 19128
rect 10594 19116 10600 19168
rect 10652 19156 10658 19168
rect 10778 19156 10784 19168
rect 10652 19128 10784 19156
rect 10652 19116 10658 19128
rect 10778 19116 10784 19128
rect 10836 19156 10842 19168
rect 11149 19159 11207 19165
rect 11149 19156 11161 19159
rect 10836 19128 11161 19156
rect 10836 19116 10842 19128
rect 11149 19125 11161 19128
rect 11195 19125 11207 19159
rect 11149 19119 11207 19125
rect 14274 19116 14280 19168
rect 14332 19156 14338 19168
rect 15749 19159 15807 19165
rect 15749 19156 15761 19159
rect 14332 19128 15761 19156
rect 14332 19116 14338 19128
rect 15749 19125 15761 19128
rect 15795 19156 15807 19159
rect 16298 19156 16304 19168
rect 15795 19128 16304 19156
rect 15795 19125 15807 19128
rect 15749 19119 15807 19125
rect 16298 19116 16304 19128
rect 16356 19116 16362 19168
rect 17310 19156 17316 19168
rect 17271 19128 17316 19156
rect 17310 19116 17316 19128
rect 17368 19116 17374 19168
rect 21542 19156 21548 19168
rect 21503 19128 21548 19156
rect 21542 19116 21548 19128
rect 21600 19116 21606 19168
rect 21910 19116 21916 19168
rect 21968 19156 21974 19168
rect 22005 19159 22063 19165
rect 22005 19156 22017 19159
rect 21968 19128 22017 19156
rect 21968 19116 21974 19128
rect 22005 19125 22017 19128
rect 22051 19125 22063 19159
rect 22005 19119 22063 19125
rect 22465 19159 22523 19165
rect 22465 19125 22477 19159
rect 22511 19156 22523 19159
rect 22646 19156 22652 19168
rect 22511 19128 22652 19156
rect 22511 19125 22523 19128
rect 22465 19119 22523 19125
rect 22646 19116 22652 19128
rect 22704 19116 22710 19168
rect 25240 19165 25268 19196
rect 25685 19193 25697 19196
rect 25731 19224 25743 19227
rect 25866 19224 25872 19236
rect 25731 19196 25872 19224
rect 25731 19193 25743 19196
rect 25685 19187 25743 19193
rect 25866 19184 25872 19196
rect 25924 19184 25930 19236
rect 25225 19159 25283 19165
rect 25225 19125 25237 19159
rect 25271 19125 25283 19159
rect 25225 19119 25283 19125
rect 26605 19159 26663 19165
rect 26605 19125 26617 19159
rect 26651 19156 26663 19159
rect 26786 19156 26792 19168
rect 26651 19128 26792 19156
rect 26651 19125 26663 19128
rect 26605 19119 26663 19125
rect 26786 19116 26792 19128
rect 26844 19116 26850 19168
rect 1104 19066 28888 19088
rect 1104 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 20982 19066
rect 21034 19014 21046 19066
rect 21098 19014 21110 19066
rect 21162 19014 21174 19066
rect 21226 19014 28888 19066
rect 1104 18992 28888 19014
rect 3050 18912 3056 18964
rect 3108 18952 3114 18964
rect 3418 18952 3424 18964
rect 3108 18924 3424 18952
rect 3108 18912 3114 18924
rect 3418 18912 3424 18924
rect 3476 18912 3482 18964
rect 6181 18955 6239 18961
rect 6181 18921 6193 18955
rect 6227 18952 6239 18955
rect 7190 18952 7196 18964
rect 6227 18924 7196 18952
rect 6227 18921 6239 18924
rect 6181 18915 6239 18921
rect 7190 18912 7196 18924
rect 7248 18912 7254 18964
rect 7558 18952 7564 18964
rect 7519 18924 7564 18952
rect 7558 18912 7564 18924
rect 7616 18912 7622 18964
rect 8294 18952 8300 18964
rect 8255 18924 8300 18952
rect 8294 18912 8300 18924
rect 8352 18912 8358 18964
rect 13633 18955 13691 18961
rect 13633 18921 13645 18955
rect 13679 18952 13691 18955
rect 13722 18952 13728 18964
rect 13679 18924 13728 18952
rect 13679 18921 13691 18924
rect 13633 18915 13691 18921
rect 13722 18912 13728 18924
rect 13780 18912 13786 18964
rect 15838 18952 15844 18964
rect 15799 18924 15844 18952
rect 15838 18912 15844 18924
rect 15896 18952 15902 18964
rect 16577 18955 16635 18961
rect 16577 18952 16589 18955
rect 15896 18924 16589 18952
rect 15896 18912 15902 18924
rect 16577 18921 16589 18924
rect 16623 18921 16635 18955
rect 16577 18915 16635 18921
rect 22097 18955 22155 18961
rect 22097 18921 22109 18955
rect 22143 18952 22155 18955
rect 22646 18952 22652 18964
rect 22143 18924 22652 18952
rect 22143 18921 22155 18924
rect 22097 18915 22155 18921
rect 22646 18912 22652 18924
rect 22704 18912 22710 18964
rect 23750 18912 23756 18964
rect 23808 18952 23814 18964
rect 24397 18955 24455 18961
rect 24397 18952 24409 18955
rect 23808 18924 24409 18952
rect 23808 18912 23814 18924
rect 24397 18921 24409 18924
rect 24443 18921 24455 18955
rect 24397 18915 24455 18921
rect 4154 18844 4160 18896
rect 4212 18884 4218 18896
rect 4430 18884 4436 18896
rect 4212 18856 4436 18884
rect 4212 18844 4218 18856
rect 4430 18844 4436 18856
rect 4488 18844 4494 18896
rect 6730 18844 6736 18896
rect 6788 18884 6794 18896
rect 6917 18887 6975 18893
rect 6917 18884 6929 18887
rect 6788 18856 6929 18884
rect 6788 18844 6794 18856
rect 6917 18853 6929 18856
rect 6963 18884 6975 18887
rect 7374 18884 7380 18896
rect 6963 18856 7380 18884
rect 6963 18853 6975 18856
rect 6917 18847 6975 18853
rect 7374 18844 7380 18856
rect 7432 18884 7438 18896
rect 8754 18884 8760 18896
rect 7432 18856 8760 18884
rect 7432 18844 7438 18856
rect 8754 18844 8760 18856
rect 8812 18844 8818 18896
rect 10870 18893 10876 18896
rect 10864 18884 10876 18893
rect 10783 18856 10876 18884
rect 10864 18847 10876 18856
rect 10928 18884 10934 18896
rect 11422 18884 11428 18896
rect 10928 18856 11428 18884
rect 10870 18844 10876 18847
rect 10928 18844 10934 18856
rect 11422 18844 11428 18856
rect 11480 18844 11486 18896
rect 14093 18887 14151 18893
rect 14093 18884 14105 18887
rect 13648 18856 14105 18884
rect 13648 18828 13676 18856
rect 14093 18853 14105 18856
rect 14139 18853 14151 18887
rect 14093 18847 14151 18853
rect 16209 18887 16267 18893
rect 16209 18853 16221 18887
rect 16255 18884 16267 18887
rect 16390 18884 16396 18896
rect 16255 18856 16396 18884
rect 16255 18853 16267 18856
rect 16209 18847 16267 18853
rect 16390 18844 16396 18856
rect 16448 18844 16454 18896
rect 16945 18887 17003 18893
rect 16945 18884 16957 18887
rect 16868 18856 16957 18884
rect 1762 18825 1768 18828
rect 1756 18816 1768 18825
rect 1675 18788 1768 18816
rect 1756 18779 1768 18788
rect 1820 18816 1826 18828
rect 3694 18816 3700 18828
rect 1820 18788 3700 18816
rect 1762 18776 1768 18779
rect 1820 18776 1826 18788
rect 3694 18776 3700 18788
rect 3752 18816 3758 18828
rect 3752 18788 4752 18816
rect 3752 18776 3758 18788
rect 1486 18748 1492 18760
rect 1447 18720 1492 18748
rect 1486 18708 1492 18720
rect 1544 18708 1550 18760
rect 4522 18748 4528 18760
rect 4483 18720 4528 18748
rect 4522 18708 4528 18720
rect 4580 18708 4586 18760
rect 4724 18757 4752 18788
rect 13630 18776 13636 18828
rect 13688 18776 13694 18828
rect 13814 18776 13820 18828
rect 13872 18816 13878 18828
rect 14001 18819 14059 18825
rect 14001 18816 14013 18819
rect 13872 18788 14013 18816
rect 13872 18776 13878 18788
rect 14001 18785 14013 18788
rect 14047 18785 14059 18819
rect 14001 18779 14059 18785
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18748 4767 18751
rect 4798 18748 4804 18760
rect 4755 18720 4804 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 7650 18748 7656 18760
rect 7611 18720 7656 18748
rect 7650 18708 7656 18720
rect 7708 18708 7714 18760
rect 7742 18708 7748 18760
rect 7800 18748 7806 18760
rect 7837 18751 7895 18757
rect 7837 18748 7849 18751
rect 7800 18720 7849 18748
rect 7800 18708 7806 18720
rect 7837 18717 7849 18720
rect 7883 18748 7895 18751
rect 8570 18748 8576 18760
rect 7883 18720 8576 18748
rect 7883 18717 7895 18720
rect 7837 18711 7895 18717
rect 8570 18708 8576 18720
rect 8628 18708 8634 18760
rect 10594 18748 10600 18760
rect 10555 18720 10600 18748
rect 10594 18708 10600 18720
rect 10652 18708 10658 18760
rect 14182 18748 14188 18760
rect 14143 18720 14188 18748
rect 14182 18708 14188 18720
rect 14240 18708 14246 18760
rect 12342 18640 12348 18692
rect 12400 18680 12406 18692
rect 16574 18680 16580 18692
rect 12400 18652 16580 18680
rect 12400 18640 12406 18652
rect 16574 18640 16580 18652
rect 16632 18680 16638 18692
rect 16868 18680 16896 18856
rect 16945 18853 16957 18856
rect 16991 18853 17003 18887
rect 19242 18884 19248 18896
rect 16945 18847 17003 18853
rect 18340 18856 19248 18884
rect 17034 18816 17040 18828
rect 16995 18788 17040 18816
rect 17034 18776 17040 18788
rect 17092 18776 17098 18828
rect 17862 18776 17868 18828
rect 17920 18816 17926 18828
rect 18340 18825 18368 18856
rect 19242 18844 19248 18856
rect 19300 18844 19306 18896
rect 22462 18884 22468 18896
rect 22423 18856 22468 18884
rect 22462 18844 22468 18856
rect 22520 18844 22526 18896
rect 18325 18819 18383 18825
rect 18325 18816 18337 18819
rect 17920 18788 18337 18816
rect 17920 18776 17926 18788
rect 18325 18785 18337 18788
rect 18371 18785 18383 18819
rect 18325 18779 18383 18785
rect 18414 18776 18420 18828
rect 18472 18816 18478 18828
rect 18581 18819 18639 18825
rect 18581 18816 18593 18819
rect 18472 18788 18593 18816
rect 18472 18776 18478 18788
rect 18581 18785 18593 18788
rect 18627 18785 18639 18819
rect 23014 18816 23020 18828
rect 22975 18788 23020 18816
rect 18581 18779 18639 18785
rect 23014 18776 23020 18788
rect 23072 18776 23078 18828
rect 24762 18816 24768 18828
rect 24723 18788 24768 18816
rect 24762 18776 24768 18788
rect 24820 18776 24826 18828
rect 24857 18819 24915 18825
rect 24857 18785 24869 18819
rect 24903 18816 24915 18819
rect 25130 18816 25136 18828
rect 24903 18788 25136 18816
rect 24903 18785 24915 18788
rect 24857 18779 24915 18785
rect 25130 18776 25136 18788
rect 25188 18776 25194 18828
rect 17126 18748 17132 18760
rect 17087 18720 17132 18748
rect 17126 18708 17132 18720
rect 17184 18708 17190 18760
rect 20901 18751 20959 18757
rect 20901 18717 20913 18751
rect 20947 18748 20959 18751
rect 21358 18748 21364 18760
rect 20947 18720 21364 18748
rect 20947 18717 20959 18720
rect 20901 18711 20959 18717
rect 21358 18708 21364 18720
rect 21416 18708 21422 18760
rect 23106 18748 23112 18760
rect 23067 18720 23112 18748
rect 23106 18708 23112 18720
rect 23164 18708 23170 18760
rect 23293 18751 23351 18757
rect 23293 18717 23305 18751
rect 23339 18748 23351 18751
rect 23474 18748 23480 18760
rect 23339 18720 23480 18748
rect 23339 18717 23351 18720
rect 23293 18711 23351 18717
rect 23474 18708 23480 18720
rect 23532 18708 23538 18760
rect 23753 18751 23811 18757
rect 23753 18717 23765 18751
rect 23799 18748 23811 18751
rect 24670 18748 24676 18760
rect 23799 18720 24676 18748
rect 23799 18717 23811 18720
rect 23753 18711 23811 18717
rect 24670 18708 24676 18720
rect 24728 18748 24734 18760
rect 24949 18751 25007 18757
rect 24949 18748 24961 18751
rect 24728 18720 24961 18748
rect 24728 18708 24734 18720
rect 24949 18717 24961 18720
rect 24995 18717 25007 18751
rect 24949 18711 25007 18717
rect 16632 18652 16896 18680
rect 16632 18640 16638 18652
rect 2866 18612 2872 18624
rect 2827 18584 2872 18612
rect 2866 18572 2872 18584
rect 2924 18572 2930 18624
rect 3510 18572 3516 18624
rect 3568 18612 3574 18624
rect 4065 18615 4123 18621
rect 4065 18612 4077 18615
rect 3568 18584 4077 18612
rect 3568 18572 3574 18584
rect 4065 18581 4077 18584
rect 4111 18581 4123 18615
rect 7190 18612 7196 18624
rect 7151 18584 7196 18612
rect 4065 18575 4123 18581
rect 7190 18572 7196 18584
rect 7248 18572 7254 18624
rect 8941 18615 8999 18621
rect 8941 18581 8953 18615
rect 8987 18612 8999 18615
rect 9306 18612 9312 18624
rect 8987 18584 9312 18612
rect 8987 18581 8999 18584
rect 8941 18575 8999 18581
rect 9306 18572 9312 18584
rect 9364 18612 9370 18624
rect 9766 18612 9772 18624
rect 9364 18584 9772 18612
rect 9364 18572 9370 18584
rect 9766 18572 9772 18584
rect 9824 18572 9830 18624
rect 9950 18612 9956 18624
rect 9911 18584 9956 18612
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 10410 18572 10416 18624
rect 10468 18612 10474 18624
rect 11977 18615 12035 18621
rect 11977 18612 11989 18615
rect 10468 18584 11989 18612
rect 10468 18572 10474 18584
rect 11977 18581 11989 18584
rect 12023 18581 12035 18615
rect 19702 18612 19708 18624
rect 19663 18584 19708 18612
rect 11977 18575 12035 18581
rect 19702 18572 19708 18584
rect 19760 18572 19766 18624
rect 21266 18572 21272 18624
rect 21324 18612 21330 18624
rect 21361 18615 21419 18621
rect 21361 18612 21373 18615
rect 21324 18584 21373 18612
rect 21324 18572 21330 18584
rect 21361 18581 21373 18584
rect 21407 18581 21419 18615
rect 21361 18575 21419 18581
rect 1104 18522 28888 18544
rect 1104 18470 5982 18522
rect 6034 18470 6046 18522
rect 6098 18470 6110 18522
rect 6162 18470 6174 18522
rect 6226 18470 15982 18522
rect 16034 18470 16046 18522
rect 16098 18470 16110 18522
rect 16162 18470 16174 18522
rect 16226 18470 25982 18522
rect 26034 18470 26046 18522
rect 26098 18470 26110 18522
rect 26162 18470 26174 18522
rect 26226 18470 28888 18522
rect 1104 18448 28888 18470
rect 1673 18411 1731 18417
rect 1673 18377 1685 18411
rect 1719 18408 1731 18411
rect 1762 18408 1768 18420
rect 1719 18380 1768 18408
rect 1719 18377 1731 18380
rect 1673 18371 1731 18377
rect 1762 18368 1768 18380
rect 1820 18368 1826 18420
rect 4522 18408 4528 18420
rect 4483 18380 4528 18408
rect 4522 18368 4528 18380
rect 4580 18368 4586 18420
rect 6822 18408 6828 18420
rect 6783 18380 6828 18408
rect 6822 18368 6828 18380
rect 6880 18368 6886 18420
rect 7558 18368 7564 18420
rect 7616 18408 7622 18420
rect 7837 18411 7895 18417
rect 7837 18408 7849 18411
rect 7616 18380 7849 18408
rect 7616 18368 7622 18380
rect 7837 18377 7849 18380
rect 7883 18377 7895 18411
rect 9766 18408 9772 18420
rect 9727 18380 9772 18408
rect 7837 18371 7895 18377
rect 9766 18368 9772 18380
rect 9824 18368 9830 18420
rect 10870 18408 10876 18420
rect 10831 18380 10876 18408
rect 10870 18368 10876 18380
rect 10928 18368 10934 18420
rect 13265 18411 13323 18417
rect 13265 18377 13277 18411
rect 13311 18408 13323 18411
rect 13446 18408 13452 18420
rect 13311 18380 13452 18408
rect 13311 18377 13323 18380
rect 13265 18371 13323 18377
rect 13446 18368 13452 18380
rect 13504 18408 13510 18420
rect 14182 18408 14188 18420
rect 13504 18380 14188 18408
rect 13504 18368 13510 18380
rect 14182 18368 14188 18380
rect 14240 18368 14246 18420
rect 16574 18408 16580 18420
rect 16535 18380 16580 18408
rect 16574 18368 16580 18380
rect 16632 18368 16638 18420
rect 17034 18408 17040 18420
rect 16995 18380 17040 18408
rect 17034 18368 17040 18380
rect 17092 18368 17098 18420
rect 17126 18368 17132 18420
rect 17184 18408 17190 18420
rect 17313 18411 17371 18417
rect 17313 18408 17325 18411
rect 17184 18380 17325 18408
rect 17184 18368 17190 18380
rect 17313 18377 17325 18380
rect 17359 18377 17371 18411
rect 17862 18408 17868 18420
rect 17823 18380 17868 18408
rect 17313 18371 17371 18377
rect 17862 18368 17868 18380
rect 17920 18368 17926 18420
rect 19334 18408 19340 18420
rect 19295 18380 19340 18408
rect 19334 18368 19340 18380
rect 19392 18408 19398 18420
rect 21174 18408 21180 18420
rect 19392 18380 20300 18408
rect 21135 18380 21180 18408
rect 19392 18368 19398 18380
rect 1486 18300 1492 18352
rect 1544 18340 1550 18352
rect 1949 18343 2007 18349
rect 1949 18340 1961 18343
rect 1544 18312 1961 18340
rect 1544 18300 1550 18312
rect 1949 18309 1961 18312
rect 1995 18309 2007 18343
rect 1949 18303 2007 18309
rect 2866 18300 2872 18352
rect 2924 18340 2930 18352
rect 2961 18343 3019 18349
rect 2961 18340 2973 18343
rect 2924 18312 2973 18340
rect 2924 18300 2930 18312
rect 2961 18309 2973 18312
rect 3007 18340 3019 18343
rect 4157 18343 4215 18349
rect 3007 18312 3740 18340
rect 3007 18309 3019 18312
rect 2961 18303 3019 18309
rect 3712 18284 3740 18312
rect 4157 18309 4169 18343
rect 4203 18340 4215 18343
rect 4430 18340 4436 18352
rect 4203 18312 4436 18340
rect 4203 18309 4215 18312
rect 4157 18303 4215 18309
rect 4430 18300 4436 18312
rect 4488 18300 4494 18352
rect 6641 18343 6699 18349
rect 6641 18309 6653 18343
rect 6687 18340 6699 18343
rect 7742 18340 7748 18352
rect 6687 18312 7748 18340
rect 6687 18309 6699 18312
rect 6641 18303 6699 18309
rect 7742 18300 7748 18312
rect 7800 18300 7806 18352
rect 13814 18300 13820 18352
rect 13872 18340 13878 18352
rect 14093 18343 14151 18349
rect 14093 18340 14105 18343
rect 13872 18312 14105 18340
rect 13872 18300 13878 18312
rect 14093 18309 14105 18312
rect 14139 18309 14151 18343
rect 16592 18340 16620 18368
rect 19613 18343 19671 18349
rect 19613 18340 19625 18343
rect 16592 18312 19625 18340
rect 14093 18303 14151 18309
rect 19613 18309 19625 18312
rect 19659 18340 19671 18343
rect 19659 18312 20208 18340
rect 19659 18309 19671 18312
rect 19613 18303 19671 18309
rect 2593 18275 2651 18281
rect 2593 18241 2605 18275
rect 2639 18272 2651 18275
rect 3510 18272 3516 18284
rect 2639 18244 3516 18272
rect 2639 18241 2651 18244
rect 2593 18235 2651 18241
rect 3510 18232 3516 18244
rect 3568 18232 3574 18284
rect 3694 18272 3700 18284
rect 3655 18244 3700 18272
rect 3694 18232 3700 18244
rect 3752 18232 3758 18284
rect 6273 18275 6331 18281
rect 6273 18241 6285 18275
rect 6319 18272 6331 18275
rect 7190 18272 7196 18284
rect 6319 18244 7196 18272
rect 6319 18241 6331 18244
rect 6273 18235 6331 18241
rect 7190 18232 7196 18244
rect 7248 18232 7254 18284
rect 7374 18272 7380 18284
rect 7335 18244 7380 18272
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 9582 18232 9588 18284
rect 9640 18272 9646 18284
rect 9677 18275 9735 18281
rect 9677 18272 9689 18275
rect 9640 18244 9689 18272
rect 9640 18232 9646 18244
rect 9677 18241 9689 18244
rect 9723 18272 9735 18275
rect 10410 18272 10416 18284
rect 9723 18244 10416 18272
rect 9723 18241 9735 18244
rect 9677 18235 9735 18241
rect 10410 18232 10416 18244
rect 10468 18232 10474 18284
rect 13538 18232 13544 18284
rect 13596 18272 13602 18284
rect 13633 18275 13691 18281
rect 13633 18272 13645 18275
rect 13596 18244 13645 18272
rect 13596 18232 13602 18244
rect 13633 18241 13645 18244
rect 13679 18272 13691 18275
rect 14734 18272 14740 18284
rect 13679 18244 14740 18272
rect 13679 18241 13691 18244
rect 13633 18235 13691 18241
rect 14734 18232 14740 18244
rect 14792 18232 14798 18284
rect 3418 18204 3424 18216
rect 3379 18176 3424 18204
rect 3418 18164 3424 18176
rect 3476 18164 3482 18216
rect 7208 18204 7236 18232
rect 20180 18216 20208 18312
rect 20272 18281 20300 18380
rect 21174 18368 21180 18380
rect 21232 18368 21238 18420
rect 21542 18368 21548 18420
rect 21600 18408 21606 18420
rect 22741 18411 22799 18417
rect 22741 18408 22753 18411
rect 21600 18380 22753 18408
rect 21600 18368 21606 18380
rect 22741 18377 22753 18380
rect 22787 18408 22799 18411
rect 23474 18408 23480 18420
rect 22787 18380 23480 18408
rect 22787 18377 22799 18380
rect 22741 18371 22799 18377
rect 23474 18368 23480 18380
rect 23532 18368 23538 18420
rect 26326 18368 26332 18420
rect 26384 18408 26390 18420
rect 27525 18411 27583 18417
rect 27525 18408 27537 18411
rect 26384 18380 27537 18408
rect 26384 18368 26390 18380
rect 27525 18377 27537 18380
rect 27571 18377 27583 18411
rect 27525 18371 27583 18377
rect 20714 18300 20720 18352
rect 20772 18340 20778 18352
rect 21361 18343 21419 18349
rect 21361 18340 21373 18343
rect 20772 18312 21373 18340
rect 20772 18300 20778 18312
rect 21361 18309 21373 18312
rect 21407 18309 21419 18343
rect 21361 18303 21419 18309
rect 23014 18300 23020 18352
rect 23072 18340 23078 18352
rect 23661 18343 23719 18349
rect 23661 18340 23673 18343
rect 23072 18312 23673 18340
rect 23072 18300 23078 18312
rect 23661 18309 23673 18312
rect 23707 18309 23719 18343
rect 25130 18340 25136 18352
rect 25091 18312 25136 18340
rect 23661 18303 23719 18309
rect 25130 18300 25136 18312
rect 25188 18300 25194 18352
rect 20257 18275 20315 18281
rect 20257 18241 20269 18275
rect 20303 18241 20315 18275
rect 20257 18235 20315 18241
rect 20349 18275 20407 18281
rect 20349 18241 20361 18275
rect 20395 18272 20407 18275
rect 21266 18272 21272 18284
rect 20395 18244 21272 18272
rect 20395 18241 20407 18244
rect 20349 18235 20407 18241
rect 7285 18207 7343 18213
rect 7285 18204 7297 18207
rect 7208 18176 7297 18204
rect 7285 18173 7297 18176
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 9950 18164 9956 18216
rect 10008 18204 10014 18216
rect 10137 18207 10195 18213
rect 10137 18204 10149 18207
rect 10008 18176 10149 18204
rect 10008 18164 10014 18176
rect 10137 18173 10149 18176
rect 10183 18173 10195 18207
rect 20162 18204 20168 18216
rect 20075 18176 20168 18204
rect 10137 18167 10195 18173
rect 20162 18164 20168 18176
rect 20220 18164 20226 18216
rect 7098 18096 7104 18148
rect 7156 18136 7162 18148
rect 7193 18139 7251 18145
rect 7193 18136 7205 18139
rect 7156 18108 7205 18136
rect 7156 18096 7162 18108
rect 7193 18105 7205 18108
rect 7239 18105 7251 18139
rect 7193 18099 7251 18105
rect 9309 18139 9367 18145
rect 9309 18105 9321 18139
rect 9355 18136 9367 18139
rect 10229 18139 10287 18145
rect 10229 18136 10241 18139
rect 9355 18108 10241 18136
rect 9355 18105 9367 18108
rect 9309 18099 9367 18105
rect 10229 18105 10241 18108
rect 10275 18136 10287 18139
rect 10318 18136 10324 18148
rect 10275 18108 10324 18136
rect 10275 18105 10287 18108
rect 10229 18099 10287 18105
rect 10318 18096 10324 18108
rect 10376 18096 10382 18148
rect 12897 18139 12955 18145
rect 12897 18105 12909 18139
rect 12943 18136 12955 18139
rect 13630 18136 13636 18148
rect 12943 18108 13636 18136
rect 12943 18105 12955 18108
rect 12897 18099 12955 18105
rect 13630 18096 13636 18108
rect 13688 18096 13694 18148
rect 20364 18136 20392 18235
rect 21266 18232 21272 18244
rect 21324 18272 21330 18284
rect 21913 18275 21971 18281
rect 21913 18272 21925 18275
rect 21324 18244 21925 18272
rect 21324 18232 21330 18244
rect 21913 18241 21925 18244
rect 21959 18241 21971 18275
rect 21913 18235 21971 18241
rect 24305 18275 24363 18281
rect 24305 18241 24317 18275
rect 24351 18272 24363 18275
rect 24670 18272 24676 18284
rect 24351 18244 24676 18272
rect 24351 18241 24363 18244
rect 24305 18235 24363 18241
rect 24670 18232 24676 18244
rect 24728 18232 24734 18284
rect 21358 18164 21364 18216
rect 21416 18204 21422 18216
rect 21729 18207 21787 18213
rect 21729 18204 21741 18207
rect 21416 18176 21741 18204
rect 21416 18164 21422 18176
rect 21729 18173 21741 18176
rect 21775 18173 21787 18207
rect 21729 18167 21787 18173
rect 23566 18164 23572 18216
rect 23624 18204 23630 18216
rect 24762 18204 24768 18216
rect 23624 18176 24768 18204
rect 23624 18164 23630 18176
rect 24762 18164 24768 18176
rect 24820 18164 24826 18216
rect 26142 18204 26148 18216
rect 26103 18176 26148 18204
rect 26142 18164 26148 18176
rect 26200 18164 26206 18216
rect 18892 18108 20392 18136
rect 3050 18068 3056 18080
rect 3011 18040 3056 18068
rect 3050 18028 3056 18040
rect 3108 18028 3114 18080
rect 4798 18068 4804 18080
rect 4759 18040 4804 18068
rect 4798 18028 4804 18040
rect 4856 18028 4862 18080
rect 10594 18028 10600 18080
rect 10652 18068 10658 18080
rect 11241 18071 11299 18077
rect 11241 18068 11253 18071
rect 10652 18040 11253 18068
rect 10652 18028 10658 18040
rect 11241 18037 11253 18040
rect 11287 18068 11299 18071
rect 12342 18068 12348 18080
rect 11287 18040 12348 18068
rect 11287 18037 11299 18040
rect 11241 18031 11299 18037
rect 12342 18028 12348 18040
rect 12400 18028 12406 18080
rect 13814 18028 13820 18080
rect 13872 18068 13878 18080
rect 13909 18071 13967 18077
rect 13909 18068 13921 18071
rect 13872 18040 13921 18068
rect 13872 18028 13878 18040
rect 13909 18037 13921 18040
rect 13955 18068 13967 18071
rect 14461 18071 14519 18077
rect 14461 18068 14473 18071
rect 13955 18040 14473 18068
rect 13955 18037 13967 18040
rect 13909 18031 13967 18037
rect 14461 18037 14473 18040
rect 14507 18037 14519 18071
rect 14461 18031 14519 18037
rect 14553 18071 14611 18077
rect 14553 18037 14565 18071
rect 14599 18068 14611 18071
rect 15197 18071 15255 18077
rect 15197 18068 15209 18071
rect 14599 18040 15209 18068
rect 14599 18037 14611 18040
rect 14553 18031 14611 18037
rect 15197 18037 15209 18040
rect 15243 18068 15255 18071
rect 15286 18068 15292 18080
rect 15243 18040 15292 18068
rect 15243 18037 15255 18040
rect 15197 18031 15255 18037
rect 15286 18028 15292 18040
rect 15344 18028 15350 18080
rect 18414 18068 18420 18080
rect 18375 18040 18420 18068
rect 18414 18028 18420 18040
rect 18472 18068 18478 18080
rect 18892 18077 18920 18108
rect 21174 18096 21180 18148
rect 21232 18136 21238 18148
rect 21818 18136 21824 18148
rect 21232 18108 21824 18136
rect 21232 18096 21238 18108
rect 21818 18096 21824 18108
rect 21876 18096 21882 18148
rect 23109 18139 23167 18145
rect 23109 18105 23121 18139
rect 23155 18136 23167 18139
rect 23934 18136 23940 18148
rect 23155 18108 23940 18136
rect 23155 18105 23167 18108
rect 23109 18099 23167 18105
rect 23934 18096 23940 18108
rect 23992 18136 23998 18148
rect 24121 18139 24179 18145
rect 24121 18136 24133 18139
rect 23992 18108 24133 18136
rect 23992 18096 23998 18108
rect 24121 18105 24133 18108
rect 24167 18105 24179 18139
rect 26390 18139 26448 18145
rect 26390 18136 26402 18139
rect 24121 18099 24179 18105
rect 25976 18108 26402 18136
rect 18877 18071 18935 18077
rect 18877 18068 18889 18071
rect 18472 18040 18889 18068
rect 18472 18028 18478 18040
rect 18877 18037 18889 18040
rect 18923 18037 18935 18071
rect 19794 18068 19800 18080
rect 19755 18040 19800 18068
rect 18877 18031 18935 18037
rect 19794 18028 19800 18040
rect 19852 18028 19858 18080
rect 23474 18068 23480 18080
rect 23387 18040 23480 18068
rect 23474 18028 23480 18040
rect 23532 18068 23538 18080
rect 24026 18068 24032 18080
rect 23532 18040 24032 18068
rect 23532 18028 23538 18040
rect 24026 18028 24032 18040
rect 24084 18028 24090 18080
rect 24854 18028 24860 18080
rect 24912 18068 24918 18080
rect 25976 18077 26004 18108
rect 26390 18105 26402 18108
rect 26436 18105 26448 18139
rect 26390 18099 26448 18105
rect 25961 18071 26019 18077
rect 25961 18068 25973 18071
rect 24912 18040 25973 18068
rect 24912 18028 24918 18040
rect 25961 18037 25973 18040
rect 26007 18037 26019 18071
rect 25961 18031 26019 18037
rect 1104 17978 28888 18000
rect 1104 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 20982 17978
rect 21034 17926 21046 17978
rect 21098 17926 21110 17978
rect 21162 17926 21174 17978
rect 21226 17926 28888 17978
rect 1104 17904 28888 17926
rect 7098 17824 7104 17876
rect 7156 17864 7162 17876
rect 7561 17867 7619 17873
rect 7561 17864 7573 17867
rect 7156 17836 7573 17864
rect 7156 17824 7162 17836
rect 7561 17833 7573 17836
rect 7607 17833 7619 17867
rect 7561 17827 7619 17833
rect 8021 17867 8079 17873
rect 8021 17833 8033 17867
rect 8067 17864 8079 17867
rect 8202 17864 8208 17876
rect 8067 17836 8208 17864
rect 8067 17833 8079 17836
rect 8021 17827 8079 17833
rect 8202 17824 8208 17836
rect 8260 17824 8266 17876
rect 10318 17864 10324 17876
rect 10279 17836 10324 17864
rect 10318 17824 10324 17836
rect 10376 17824 10382 17876
rect 13541 17867 13599 17873
rect 13541 17833 13553 17867
rect 13587 17864 13599 17867
rect 13722 17864 13728 17876
rect 13587 17836 13728 17864
rect 13587 17833 13599 17836
rect 13541 17827 13599 17833
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 17126 17824 17132 17876
rect 17184 17864 17190 17876
rect 17589 17867 17647 17873
rect 17589 17864 17601 17867
rect 17184 17836 17601 17864
rect 17184 17824 17190 17836
rect 17589 17833 17601 17836
rect 17635 17833 17647 17867
rect 17589 17827 17647 17833
rect 19705 17867 19763 17873
rect 19705 17833 19717 17867
rect 19751 17864 19763 17867
rect 19794 17864 19800 17876
rect 19751 17836 19800 17864
rect 19751 17833 19763 17836
rect 19705 17827 19763 17833
rect 19794 17824 19800 17836
rect 19852 17824 19858 17876
rect 21358 17864 21364 17876
rect 21319 17836 21364 17864
rect 21358 17824 21364 17836
rect 21416 17824 21422 17876
rect 23014 17864 23020 17876
rect 22975 17836 23020 17864
rect 23014 17824 23020 17836
rect 23072 17824 23078 17876
rect 23106 17824 23112 17876
rect 23164 17864 23170 17876
rect 23385 17867 23443 17873
rect 23385 17864 23397 17867
rect 23164 17836 23397 17864
rect 23164 17824 23170 17836
rect 23385 17833 23397 17836
rect 23431 17833 23443 17867
rect 23385 17827 23443 17833
rect 24670 17824 24676 17876
rect 24728 17864 24734 17876
rect 24765 17867 24823 17873
rect 24765 17864 24777 17867
rect 24728 17836 24777 17864
rect 24728 17824 24734 17836
rect 24765 17833 24777 17836
rect 24811 17833 24823 17867
rect 26234 17864 26240 17876
rect 26195 17836 26240 17864
rect 24765 17827 24823 17833
rect 26234 17824 26240 17836
rect 26292 17824 26298 17876
rect 7285 17799 7343 17805
rect 7285 17765 7297 17799
rect 7331 17796 7343 17799
rect 7650 17796 7656 17808
rect 7331 17768 7656 17796
rect 7331 17765 7343 17768
rect 7285 17759 7343 17765
rect 7650 17756 7656 17768
rect 7708 17756 7714 17808
rect 15102 17756 15108 17808
rect 15160 17796 15166 17808
rect 16298 17796 16304 17808
rect 15160 17768 16304 17796
rect 15160 17756 15166 17768
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 1670 17728 1676 17740
rect 1443 17700 1676 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 1670 17688 1676 17700
rect 1728 17728 1734 17740
rect 3602 17728 3608 17740
rect 1728 17700 3608 17728
rect 1728 17688 1734 17700
rect 3602 17688 3608 17700
rect 3660 17688 3666 17740
rect 5258 17728 5264 17740
rect 5219 17700 5264 17728
rect 5258 17688 5264 17700
rect 5316 17688 5322 17740
rect 5350 17688 5356 17740
rect 5408 17728 5414 17740
rect 5517 17731 5575 17737
rect 5517 17728 5529 17731
rect 5408 17700 5529 17728
rect 5408 17688 5414 17700
rect 5517 17697 5529 17700
rect 5563 17697 5575 17731
rect 5517 17691 5575 17697
rect 8018 17688 8024 17740
rect 8076 17728 8082 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 8076 17700 8401 17728
rect 8076 17688 8082 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 10686 17728 10692 17740
rect 10647 17700 10692 17728
rect 8389 17691 8447 17697
rect 10686 17688 10692 17700
rect 10744 17688 10750 17740
rect 13998 17728 14004 17740
rect 13959 17700 14004 17728
rect 13998 17688 14004 17700
rect 14056 17688 14062 17740
rect 16224 17737 16252 17768
rect 16298 17756 16304 17768
rect 16356 17796 16362 17808
rect 17862 17796 17868 17808
rect 16356 17768 17868 17796
rect 16356 17756 16362 17768
rect 17862 17756 17868 17768
rect 17920 17756 17926 17808
rect 19613 17799 19671 17805
rect 19613 17765 19625 17799
rect 19659 17796 19671 17799
rect 20070 17796 20076 17808
rect 19659 17768 20076 17796
rect 19659 17765 19671 17768
rect 19613 17759 19671 17765
rect 20070 17756 20076 17768
rect 20128 17796 20134 17808
rect 20622 17796 20628 17808
rect 20128 17768 20628 17796
rect 20128 17756 20134 17768
rect 20622 17756 20628 17768
rect 20680 17756 20686 17808
rect 22741 17799 22799 17805
rect 22741 17765 22753 17799
rect 22787 17796 22799 17799
rect 23124 17796 23152 17824
rect 22787 17768 23152 17796
rect 22787 17765 22799 17768
rect 22741 17759 22799 17765
rect 16482 17737 16488 17740
rect 16209 17731 16267 17737
rect 16209 17697 16221 17731
rect 16255 17697 16267 17731
rect 16476 17728 16488 17737
rect 16443 17700 16488 17728
rect 16209 17691 16267 17697
rect 16476 17691 16488 17700
rect 16482 17688 16488 17691
rect 16540 17688 16546 17740
rect 23750 17728 23756 17740
rect 23711 17700 23756 17728
rect 23750 17688 23756 17700
rect 23808 17688 23814 17740
rect 23845 17731 23903 17737
rect 23845 17697 23857 17731
rect 23891 17728 23903 17731
rect 24026 17728 24032 17740
rect 23891 17700 24032 17728
rect 23891 17697 23903 17700
rect 23845 17691 23903 17697
rect 24026 17688 24032 17700
rect 24084 17688 24090 17740
rect 8478 17660 8484 17672
rect 8439 17632 8484 17660
rect 8478 17620 8484 17632
rect 8536 17620 8542 17672
rect 8570 17620 8576 17672
rect 8628 17660 8634 17672
rect 8665 17663 8723 17669
rect 8665 17660 8677 17663
rect 8628 17632 8677 17660
rect 8628 17620 8634 17632
rect 8665 17629 8677 17632
rect 8711 17660 8723 17663
rect 9582 17660 9588 17672
rect 8711 17632 9588 17660
rect 8711 17629 8723 17632
rect 8665 17623 8723 17629
rect 9582 17620 9588 17632
rect 9640 17620 9646 17672
rect 10778 17660 10784 17672
rect 10739 17632 10784 17660
rect 10778 17620 10784 17632
rect 10836 17620 10842 17672
rect 10870 17620 10876 17672
rect 10928 17660 10934 17672
rect 14090 17660 14096 17672
rect 10928 17632 10973 17660
rect 14051 17632 14096 17660
rect 10928 17620 10934 17632
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 14277 17663 14335 17669
rect 14277 17629 14289 17663
rect 14323 17660 14335 17663
rect 14734 17660 14740 17672
rect 14323 17632 14740 17660
rect 14323 17629 14335 17632
rect 14277 17623 14335 17629
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 19702 17620 19708 17672
rect 19760 17660 19766 17672
rect 19797 17663 19855 17669
rect 19797 17660 19809 17663
rect 19760 17632 19809 17660
rect 19760 17620 19766 17632
rect 19797 17629 19809 17632
rect 19843 17629 19855 17663
rect 19797 17623 19855 17629
rect 23106 17620 23112 17672
rect 23164 17660 23170 17672
rect 23937 17663 23995 17669
rect 23937 17660 23949 17663
rect 23164 17632 23949 17660
rect 23164 17620 23170 17632
rect 23937 17629 23949 17632
rect 23983 17660 23995 17663
rect 24688 17660 24716 17824
rect 23983 17632 24716 17660
rect 23983 17629 23995 17632
rect 23937 17623 23995 17629
rect 10045 17595 10103 17601
rect 10045 17561 10057 17595
rect 10091 17592 10103 17595
rect 10888 17592 10916 17620
rect 13630 17592 13636 17604
rect 10091 17564 10916 17592
rect 13591 17564 13636 17592
rect 10091 17561 10103 17564
rect 10045 17555 10103 17561
rect 13630 17552 13636 17564
rect 13688 17552 13694 17604
rect 18230 17592 18236 17604
rect 18191 17564 18236 17592
rect 18230 17552 18236 17564
rect 18288 17552 18294 17604
rect 1578 17524 1584 17536
rect 1539 17496 1584 17524
rect 1578 17484 1584 17496
rect 1636 17484 1642 17536
rect 2866 17524 2872 17536
rect 2827 17496 2872 17524
rect 2866 17484 2872 17496
rect 2924 17484 2930 17536
rect 3142 17524 3148 17536
rect 3103 17496 3148 17524
rect 3142 17484 3148 17496
rect 3200 17484 3206 17536
rect 6641 17527 6699 17533
rect 6641 17493 6653 17527
rect 6687 17524 6699 17527
rect 7098 17524 7104 17536
rect 6687 17496 7104 17524
rect 6687 17493 6699 17496
rect 6641 17487 6699 17493
rect 7098 17484 7104 17496
rect 7156 17484 7162 17536
rect 15746 17484 15752 17536
rect 15804 17524 15810 17536
rect 16025 17527 16083 17533
rect 16025 17524 16037 17527
rect 15804 17496 16037 17524
rect 15804 17484 15810 17496
rect 16025 17493 16037 17496
rect 16071 17524 16083 17527
rect 16390 17524 16396 17536
rect 16071 17496 16396 17524
rect 16071 17493 16083 17496
rect 16025 17487 16083 17493
rect 16390 17484 16396 17496
rect 16448 17484 16454 17536
rect 19242 17524 19248 17536
rect 19203 17496 19248 17524
rect 19242 17484 19248 17496
rect 19300 17484 19306 17536
rect 24489 17527 24547 17533
rect 24489 17493 24501 17527
rect 24535 17524 24547 17527
rect 24670 17524 24676 17536
rect 24535 17496 24676 17524
rect 24535 17493 24547 17496
rect 24489 17487 24547 17493
rect 24670 17484 24676 17496
rect 24728 17484 24734 17536
rect 1104 17434 28888 17456
rect 1104 17382 5982 17434
rect 6034 17382 6046 17434
rect 6098 17382 6110 17434
rect 6162 17382 6174 17434
rect 6226 17382 15982 17434
rect 16034 17382 16046 17434
rect 16098 17382 16110 17434
rect 16162 17382 16174 17434
rect 16226 17382 25982 17434
rect 26034 17382 26046 17434
rect 26098 17382 26110 17434
rect 26162 17382 26174 17434
rect 26226 17382 28888 17434
rect 1104 17360 28888 17382
rect 2038 17320 2044 17332
rect 1999 17292 2044 17320
rect 2038 17280 2044 17292
rect 2096 17280 2102 17332
rect 5350 17320 5356 17332
rect 5311 17292 5356 17320
rect 5350 17280 5356 17292
rect 5408 17280 5414 17332
rect 8478 17280 8484 17332
rect 8536 17320 8542 17332
rect 8757 17323 8815 17329
rect 8757 17320 8769 17323
rect 8536 17292 8769 17320
rect 8536 17280 8542 17292
rect 8757 17289 8769 17292
rect 8803 17320 8815 17323
rect 9953 17323 10011 17329
rect 9953 17320 9965 17323
rect 8803 17292 9965 17320
rect 8803 17289 8815 17292
rect 8757 17283 8815 17289
rect 9953 17289 9965 17292
rect 9999 17289 10011 17323
rect 9953 17283 10011 17289
rect 10870 17280 10876 17332
rect 10928 17320 10934 17332
rect 11333 17323 11391 17329
rect 11333 17320 11345 17323
rect 10928 17292 11345 17320
rect 10928 17280 10934 17292
rect 11333 17289 11345 17292
rect 11379 17289 11391 17323
rect 11333 17283 11391 17289
rect 12897 17323 12955 17329
rect 12897 17289 12909 17323
rect 12943 17320 12955 17323
rect 13998 17320 14004 17332
rect 12943 17292 14004 17320
rect 12943 17289 12955 17292
rect 12897 17283 12955 17289
rect 13998 17280 14004 17292
rect 14056 17320 14062 17332
rect 14461 17323 14519 17329
rect 14461 17320 14473 17323
rect 14056 17292 14473 17320
rect 14056 17280 14062 17292
rect 14461 17289 14473 17292
rect 14507 17289 14519 17323
rect 17770 17320 17776 17332
rect 17731 17292 17776 17320
rect 14461 17283 14519 17289
rect 17770 17280 17776 17292
rect 17828 17280 17834 17332
rect 19705 17323 19763 17329
rect 19705 17289 19717 17323
rect 19751 17320 19763 17323
rect 19794 17320 19800 17332
rect 19751 17292 19800 17320
rect 19751 17289 19763 17292
rect 19705 17283 19763 17289
rect 19794 17280 19800 17292
rect 19852 17280 19858 17332
rect 20070 17320 20076 17332
rect 20031 17292 20076 17320
rect 20070 17280 20076 17292
rect 20128 17280 20134 17332
rect 23106 17320 23112 17332
rect 23067 17292 23112 17320
rect 23106 17280 23112 17292
rect 23164 17280 23170 17332
rect 2685 17255 2743 17261
rect 2685 17221 2697 17255
rect 2731 17252 2743 17255
rect 2731 17224 3464 17252
rect 2731 17221 2743 17224
rect 2685 17215 2743 17221
rect 2866 17144 2872 17196
rect 2924 17184 2930 17196
rect 3234 17184 3240 17196
rect 2924 17156 3240 17184
rect 2924 17144 2930 17156
rect 3234 17144 3240 17156
rect 3292 17144 3298 17196
rect 3436 17193 3464 17224
rect 3421 17187 3479 17193
rect 3421 17153 3433 17187
rect 3467 17184 3479 17187
rect 3694 17184 3700 17196
rect 3467 17156 3700 17184
rect 3467 17153 3479 17156
rect 3421 17147 3479 17153
rect 3694 17144 3700 17156
rect 3752 17184 3758 17196
rect 5368 17184 5396 17280
rect 9490 17252 9496 17264
rect 9403 17224 9496 17252
rect 9490 17212 9496 17224
rect 9548 17252 9554 17264
rect 10686 17252 10692 17264
rect 9548 17224 10692 17252
rect 9548 17212 9554 17224
rect 10686 17212 10692 17224
rect 10744 17212 10750 17264
rect 3752 17156 5396 17184
rect 8481 17187 8539 17193
rect 3752 17144 3758 17156
rect 8481 17153 8493 17187
rect 8527 17184 8539 17187
rect 8570 17184 8576 17196
rect 8527 17156 8576 17184
rect 8527 17153 8539 17156
rect 8481 17147 8539 17153
rect 8570 17144 8576 17156
rect 8628 17144 8634 17196
rect 10597 17187 10655 17193
rect 10597 17153 10609 17187
rect 10643 17184 10655 17187
rect 10888 17184 10916 17280
rect 13265 17255 13323 17261
rect 13265 17221 13277 17255
rect 13311 17252 13323 17255
rect 14090 17252 14096 17264
rect 13311 17224 14096 17252
rect 13311 17221 13323 17224
rect 13265 17215 13323 17221
rect 14090 17212 14096 17224
rect 14148 17252 14154 17264
rect 16025 17255 16083 17261
rect 16025 17252 16037 17255
rect 14148 17224 16037 17252
rect 14148 17212 14154 17224
rect 16025 17221 16037 17224
rect 16071 17221 16083 17255
rect 16025 17215 16083 17221
rect 17497 17255 17555 17261
rect 17497 17221 17509 17255
rect 17543 17252 17555 17255
rect 18414 17252 18420 17264
rect 17543 17224 18420 17252
rect 17543 17221 17555 17224
rect 17497 17215 17555 17221
rect 18414 17212 18420 17224
rect 18472 17252 18478 17264
rect 18472 17224 18828 17252
rect 18472 17212 18478 17224
rect 13538 17184 13544 17196
rect 10643 17156 10916 17184
rect 13499 17156 13544 17184
rect 10643 17153 10655 17156
rect 10597 17147 10655 17153
rect 13538 17144 13544 17156
rect 13596 17144 13602 17196
rect 13906 17144 13912 17196
rect 13964 17184 13970 17196
rect 15013 17187 15071 17193
rect 15013 17184 15025 17187
rect 13964 17156 15025 17184
rect 13964 17144 13970 17156
rect 15013 17153 15025 17156
rect 15059 17184 15071 17187
rect 15473 17187 15531 17193
rect 15473 17184 15485 17187
rect 15059 17156 15485 17184
rect 15059 17153 15071 17156
rect 15013 17147 15071 17153
rect 15473 17153 15485 17156
rect 15519 17184 15531 17187
rect 15838 17184 15844 17196
rect 15519 17156 15844 17184
rect 15519 17153 15531 17156
rect 15473 17147 15531 17153
rect 15838 17144 15844 17156
rect 15896 17184 15902 17196
rect 16482 17184 16488 17196
rect 15896 17156 16488 17184
rect 15896 17144 15902 17156
rect 16482 17144 16488 17156
rect 16540 17184 16546 17196
rect 16577 17187 16635 17193
rect 16577 17184 16589 17187
rect 16540 17156 16589 17184
rect 16540 17144 16546 17156
rect 16577 17153 16589 17156
rect 16623 17184 16635 17187
rect 17037 17187 17095 17193
rect 17037 17184 17049 17187
rect 16623 17156 17049 17184
rect 16623 17153 16635 17156
rect 16577 17147 16635 17153
rect 17037 17153 17049 17156
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 18230 17144 18236 17196
rect 18288 17184 18294 17196
rect 18800 17193 18828 17224
rect 18601 17187 18659 17193
rect 18601 17184 18613 17187
rect 18288 17156 18613 17184
rect 18288 17144 18294 17156
rect 18601 17153 18613 17156
rect 18647 17153 18659 17187
rect 18601 17147 18659 17153
rect 18785 17187 18843 17193
rect 18785 17153 18797 17187
rect 18831 17184 18843 17187
rect 18874 17184 18880 17196
rect 18831 17156 18880 17184
rect 18831 17153 18843 17156
rect 18785 17147 18843 17153
rect 18874 17144 18880 17156
rect 18932 17144 18938 17196
rect 19337 17187 19395 17193
rect 19337 17153 19349 17187
rect 19383 17184 19395 17187
rect 19702 17184 19708 17196
rect 19383 17156 19708 17184
rect 19383 17153 19395 17156
rect 19337 17147 19395 17153
rect 19702 17144 19708 17156
rect 19760 17144 19766 17196
rect 24670 17184 24676 17196
rect 24631 17156 24676 17184
rect 24670 17144 24676 17156
rect 24728 17144 24734 17196
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 2038 17116 2044 17128
rect 1443 17088 2044 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 3142 17116 3148 17128
rect 3103 17088 3148 17116
rect 3142 17076 3148 17088
rect 3200 17076 3206 17128
rect 5258 17076 5264 17128
rect 5316 17116 5322 17128
rect 5629 17119 5687 17125
rect 5629 17116 5641 17119
rect 5316 17088 5641 17116
rect 5316 17076 5322 17088
rect 5629 17085 5641 17088
rect 5675 17085 5687 17119
rect 14826 17116 14832 17128
rect 14787 17088 14832 17116
rect 5629 17079 5687 17085
rect 14826 17076 14832 17088
rect 14884 17076 14890 17128
rect 16390 17116 16396 17128
rect 16351 17088 16396 17116
rect 16390 17076 16396 17088
rect 16448 17116 16454 17128
rect 16758 17116 16764 17128
rect 16448 17088 16764 17116
rect 16448 17076 16454 17088
rect 16758 17076 16764 17088
rect 16816 17076 16822 17128
rect 17770 17076 17776 17128
rect 17828 17116 17834 17128
rect 18506 17116 18512 17128
rect 17828 17088 18512 17116
rect 17828 17076 17834 17088
rect 18506 17076 18512 17088
rect 18564 17076 18570 17128
rect 23474 17116 23480 17128
rect 23387 17088 23480 17116
rect 23474 17076 23480 17088
rect 23532 17116 23538 17128
rect 26418 17116 26424 17128
rect 23532 17088 24624 17116
rect 26379 17088 26424 17116
rect 23532 17076 23538 17088
rect 9861 17051 9919 17057
rect 9861 17017 9873 17051
rect 9907 17048 9919 17051
rect 10226 17048 10232 17060
rect 9907 17020 10232 17048
rect 9907 17017 9919 17020
rect 9861 17011 9919 17017
rect 10226 17008 10232 17020
rect 10284 17048 10290 17060
rect 10413 17051 10471 17057
rect 10413 17048 10425 17051
rect 10284 17020 10425 17048
rect 10284 17008 10290 17020
rect 10413 17017 10425 17020
rect 10459 17017 10471 17051
rect 10413 17011 10471 17017
rect 10778 17008 10784 17060
rect 10836 17048 10842 17060
rect 11057 17051 11115 17057
rect 11057 17048 11069 17051
rect 10836 17020 11069 17048
rect 10836 17008 10842 17020
rect 11057 17017 11069 17020
rect 11103 17048 11115 17051
rect 15933 17051 15991 17057
rect 15933 17048 15945 17051
rect 11103 17020 15945 17048
rect 11103 17017 11115 17020
rect 11057 17011 11115 17017
rect 15933 17017 15945 17020
rect 15979 17048 15991 17051
rect 16485 17051 16543 17057
rect 16485 17048 16497 17051
rect 15979 17020 16497 17048
rect 15979 17017 15991 17020
rect 15933 17011 15991 17017
rect 16485 17017 16497 17020
rect 16531 17048 16543 17051
rect 18598 17048 18604 17060
rect 16531 17020 18604 17048
rect 16531 17017 16543 17020
rect 16485 17011 16543 17017
rect 18598 17008 18604 17020
rect 18656 17008 18662 17060
rect 22741 17051 22799 17057
rect 22741 17017 22753 17051
rect 22787 17048 22799 17051
rect 23750 17048 23756 17060
rect 22787 17020 23756 17048
rect 22787 17017 22799 17020
rect 22741 17011 22799 17017
rect 23750 17008 23756 17020
rect 23808 17008 23814 17060
rect 24489 17051 24547 17057
rect 24489 17048 24501 17051
rect 23860 17020 24501 17048
rect 23860 16992 23888 17020
rect 24489 17017 24501 17020
rect 24535 17017 24547 17051
rect 24489 17011 24547 17017
rect 24596 17048 24624 17088
rect 26418 17076 26424 17088
rect 26476 17116 26482 17128
rect 26973 17119 27031 17125
rect 26973 17116 26985 17119
rect 26476 17088 26985 17116
rect 26476 17076 26482 17088
rect 26973 17085 26985 17088
rect 27019 17085 27031 17119
rect 26973 17079 27031 17085
rect 27338 17048 27344 17060
rect 24596 17020 27344 17048
rect 1581 16983 1639 16989
rect 1581 16949 1593 16983
rect 1627 16980 1639 16983
rect 1854 16980 1860 16992
rect 1627 16952 1860 16980
rect 1627 16949 1639 16952
rect 1581 16943 1639 16949
rect 1854 16940 1860 16952
rect 1912 16940 1918 16992
rect 2777 16983 2835 16989
rect 2777 16949 2789 16983
rect 2823 16980 2835 16983
rect 4062 16980 4068 16992
rect 2823 16952 4068 16980
rect 2823 16949 2835 16952
rect 2777 16943 2835 16949
rect 4062 16940 4068 16952
rect 4120 16940 4126 16992
rect 8018 16980 8024 16992
rect 7979 16952 8024 16980
rect 8018 16940 8024 16952
rect 8076 16940 8082 16992
rect 10318 16980 10324 16992
rect 10279 16952 10324 16980
rect 10318 16940 10324 16952
rect 10376 16940 10382 16992
rect 13906 16980 13912 16992
rect 13867 16952 13912 16980
rect 13906 16940 13912 16952
rect 13964 16940 13970 16992
rect 14369 16983 14427 16989
rect 14369 16949 14381 16983
rect 14415 16980 14427 16983
rect 14918 16980 14924 16992
rect 14415 16952 14924 16980
rect 14415 16949 14427 16952
rect 14369 16943 14427 16949
rect 14918 16940 14924 16952
rect 14976 16940 14982 16992
rect 17954 16940 17960 16992
rect 18012 16980 18018 16992
rect 18141 16983 18199 16989
rect 18141 16980 18153 16983
rect 18012 16952 18153 16980
rect 18012 16940 18018 16952
rect 18141 16949 18153 16952
rect 18187 16949 18199 16983
rect 23842 16980 23848 16992
rect 23803 16952 23848 16980
rect 18141 16943 18199 16949
rect 23842 16940 23848 16952
rect 23900 16940 23906 16992
rect 24026 16980 24032 16992
rect 23987 16952 24032 16980
rect 24026 16940 24032 16952
rect 24084 16940 24090 16992
rect 24397 16983 24455 16989
rect 24397 16949 24409 16983
rect 24443 16980 24455 16983
rect 24596 16980 24624 17020
rect 27338 17008 27344 17020
rect 27396 17008 27402 17060
rect 24443 16952 24624 16980
rect 24443 16949 24455 16952
rect 24397 16943 24455 16949
rect 25866 16940 25872 16992
rect 25924 16980 25930 16992
rect 26605 16983 26663 16989
rect 26605 16980 26617 16983
rect 25924 16952 26617 16980
rect 25924 16940 25930 16952
rect 26605 16949 26617 16952
rect 26651 16949 26663 16983
rect 26605 16943 26663 16949
rect 1104 16890 28888 16912
rect 1104 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 20982 16890
rect 21034 16838 21046 16890
rect 21098 16838 21110 16890
rect 21162 16838 21174 16890
rect 21226 16838 28888 16890
rect 1104 16816 28888 16838
rect 1670 16776 1676 16788
rect 1631 16748 1676 16776
rect 1670 16736 1676 16748
rect 1728 16736 1734 16788
rect 2409 16779 2467 16785
rect 2409 16745 2421 16779
rect 2455 16776 2467 16779
rect 3142 16776 3148 16788
rect 2455 16748 3148 16776
rect 2455 16745 2467 16748
rect 2409 16739 2467 16745
rect 3142 16736 3148 16748
rect 3200 16736 3206 16788
rect 4341 16779 4399 16785
rect 4341 16745 4353 16779
rect 4387 16776 4399 16779
rect 4798 16776 4804 16788
rect 4387 16748 4804 16776
rect 4387 16745 4399 16748
rect 4341 16739 4399 16745
rect 4798 16736 4804 16748
rect 4856 16736 4862 16788
rect 4982 16736 4988 16788
rect 5040 16776 5046 16788
rect 5261 16779 5319 16785
rect 5261 16776 5273 16779
rect 5040 16748 5273 16776
rect 5040 16736 5046 16748
rect 5261 16745 5273 16748
rect 5307 16745 5319 16779
rect 5718 16776 5724 16788
rect 5679 16748 5724 16776
rect 5261 16739 5319 16745
rect 5718 16736 5724 16748
rect 5776 16736 5782 16788
rect 9950 16736 9956 16788
rect 10008 16776 10014 16788
rect 10321 16779 10379 16785
rect 10321 16776 10333 16779
rect 10008 16748 10333 16776
rect 10008 16736 10014 16748
rect 10321 16745 10333 16748
rect 10367 16745 10379 16779
rect 10321 16739 10379 16745
rect 13817 16779 13875 16785
rect 13817 16745 13829 16779
rect 13863 16776 13875 16779
rect 13906 16776 13912 16788
rect 13863 16748 13912 16776
rect 13863 16745 13875 16748
rect 13817 16739 13875 16745
rect 13906 16736 13912 16748
rect 13964 16736 13970 16788
rect 14553 16779 14611 16785
rect 14553 16745 14565 16779
rect 14599 16776 14611 16779
rect 14826 16776 14832 16788
rect 14599 16748 14832 16776
rect 14599 16745 14611 16748
rect 14553 16739 14611 16745
rect 14826 16736 14832 16748
rect 14884 16736 14890 16788
rect 15286 16776 15292 16788
rect 15247 16748 15292 16776
rect 15286 16736 15292 16748
rect 15344 16736 15350 16788
rect 15746 16776 15752 16788
rect 15707 16748 15752 16776
rect 15746 16736 15752 16748
rect 15804 16736 15810 16788
rect 16298 16776 16304 16788
rect 16259 16748 16304 16776
rect 16298 16736 16304 16748
rect 16356 16736 16362 16788
rect 17954 16736 17960 16788
rect 18012 16776 18018 16788
rect 18601 16779 18659 16785
rect 18601 16776 18613 16779
rect 18012 16748 18613 16776
rect 18012 16736 18018 16748
rect 18601 16745 18613 16748
rect 18647 16745 18659 16779
rect 19242 16776 19248 16788
rect 19203 16748 19248 16776
rect 18601 16739 18659 16745
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 23477 16779 23535 16785
rect 23477 16745 23489 16779
rect 23523 16776 23535 16779
rect 24026 16776 24032 16788
rect 23523 16748 24032 16776
rect 23523 16745 23535 16748
rect 23477 16739 23535 16745
rect 24026 16736 24032 16748
rect 24084 16736 24090 16788
rect 2682 16668 2688 16720
rect 2740 16708 2746 16720
rect 2777 16711 2835 16717
rect 2777 16708 2789 16711
rect 2740 16680 2789 16708
rect 2740 16668 2746 16680
rect 2777 16677 2789 16680
rect 2823 16677 2835 16711
rect 5626 16708 5632 16720
rect 5587 16680 5632 16708
rect 2777 16671 2835 16677
rect 5626 16668 5632 16680
rect 5684 16668 5690 16720
rect 9858 16668 9864 16720
rect 9916 16708 9922 16720
rect 10689 16711 10747 16717
rect 10689 16708 10701 16711
rect 9916 16680 10701 16708
rect 9916 16668 9922 16680
rect 10689 16677 10701 16680
rect 10735 16708 10747 16711
rect 11054 16708 11060 16720
rect 10735 16680 11060 16708
rect 10735 16677 10747 16680
rect 10689 16671 10747 16677
rect 11054 16668 11060 16680
rect 11112 16668 11118 16720
rect 15654 16708 15660 16720
rect 15615 16680 15660 16708
rect 15654 16668 15660 16680
rect 15712 16668 15718 16720
rect 5258 16600 5264 16652
rect 5316 16640 5322 16652
rect 6822 16640 6828 16652
rect 5316 16612 6828 16640
rect 5316 16600 5322 16612
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 7098 16649 7104 16652
rect 7092 16640 7104 16649
rect 7059 16612 7104 16640
rect 7092 16603 7104 16612
rect 7098 16600 7104 16603
rect 7156 16600 7162 16652
rect 10781 16643 10839 16649
rect 10781 16609 10793 16643
rect 10827 16640 10839 16643
rect 10962 16640 10968 16652
rect 10827 16612 10968 16640
rect 10827 16609 10839 16612
rect 10781 16603 10839 16609
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 12526 16600 12532 16652
rect 12584 16640 12590 16652
rect 12693 16643 12751 16649
rect 12693 16640 12705 16643
rect 12584 16612 12705 16640
rect 12584 16600 12590 16612
rect 12693 16609 12705 16612
rect 12739 16609 12751 16643
rect 19702 16640 19708 16652
rect 12693 16603 12751 16609
rect 19260 16612 19708 16640
rect 2866 16572 2872 16584
rect 2827 16544 2872 16572
rect 2866 16532 2872 16544
rect 2924 16532 2930 16584
rect 3050 16572 3056 16584
rect 3011 16544 3056 16572
rect 3050 16532 3056 16544
rect 3108 16532 3114 16584
rect 5810 16532 5816 16584
rect 5868 16572 5874 16584
rect 5868 16544 5913 16572
rect 5868 16532 5874 16544
rect 10870 16532 10876 16584
rect 10928 16572 10934 16584
rect 10928 16544 10973 16572
rect 10928 16532 10934 16544
rect 12342 16532 12348 16584
rect 12400 16572 12406 16584
rect 12437 16575 12495 16581
rect 12437 16572 12449 16575
rect 12400 16544 12449 16572
rect 12400 16532 12406 16544
rect 12437 16541 12449 16544
rect 12483 16541 12495 16575
rect 15838 16572 15844 16584
rect 15799 16544 15844 16572
rect 12437 16535 12495 16541
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 18690 16572 18696 16584
rect 18651 16544 18696 16572
rect 18690 16532 18696 16544
rect 18748 16532 18754 16584
rect 18782 16532 18788 16584
rect 18840 16572 18846 16584
rect 19260 16572 19288 16612
rect 19702 16600 19708 16612
rect 19760 16640 19766 16652
rect 20990 16640 20996 16652
rect 19760 16612 20996 16640
rect 19760 16600 19766 16612
rect 20990 16600 20996 16612
rect 21048 16640 21054 16652
rect 21157 16643 21215 16649
rect 21157 16640 21169 16643
rect 21048 16612 21169 16640
rect 21048 16600 21054 16612
rect 21157 16609 21169 16612
rect 21203 16609 21215 16643
rect 21157 16603 21215 16609
rect 23750 16600 23756 16652
rect 23808 16640 23814 16652
rect 23808 16612 24072 16640
rect 23808 16600 23814 16612
rect 18840 16544 19288 16572
rect 18840 16532 18846 16544
rect 20714 16532 20720 16584
rect 20772 16572 20778 16584
rect 20901 16575 20959 16581
rect 20901 16572 20913 16575
rect 20772 16544 20913 16572
rect 20772 16532 20778 16544
rect 20901 16541 20913 16544
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 24044 16513 24072 16612
rect 24302 16600 24308 16652
rect 24360 16640 24366 16652
rect 24397 16643 24455 16649
rect 24397 16640 24409 16643
rect 24360 16612 24409 16640
rect 24360 16600 24366 16612
rect 24397 16609 24409 16612
rect 24443 16609 24455 16643
rect 24397 16603 24455 16609
rect 24486 16572 24492 16584
rect 24447 16544 24492 16572
rect 24486 16532 24492 16544
rect 24544 16532 24550 16584
rect 24670 16572 24676 16584
rect 24583 16544 24676 16572
rect 24670 16532 24676 16544
rect 24728 16572 24734 16584
rect 24854 16572 24860 16584
rect 24728 16544 24860 16572
rect 24728 16532 24734 16544
rect 24854 16532 24860 16544
rect 24912 16532 24918 16584
rect 24029 16507 24087 16513
rect 24029 16473 24041 16507
rect 24075 16473 24087 16507
rect 24029 16467 24087 16473
rect 8202 16436 8208 16448
rect 8163 16408 8208 16436
rect 8202 16396 8208 16408
rect 8260 16396 8266 16448
rect 10045 16439 10103 16445
rect 10045 16405 10057 16439
rect 10091 16436 10103 16439
rect 10318 16436 10324 16448
rect 10091 16408 10324 16436
rect 10091 16405 10103 16408
rect 10045 16399 10103 16405
rect 10318 16396 10324 16408
rect 10376 16436 10382 16448
rect 12710 16436 12716 16448
rect 10376 16408 12716 16436
rect 10376 16396 10382 16408
rect 12710 16396 12716 16408
rect 12768 16396 12774 16448
rect 18233 16439 18291 16445
rect 18233 16405 18245 16439
rect 18279 16436 18291 16439
rect 19150 16436 19156 16448
rect 18279 16408 19156 16436
rect 18279 16405 18291 16408
rect 18233 16399 18291 16405
rect 19150 16396 19156 16408
rect 19208 16396 19214 16448
rect 21818 16396 21824 16448
rect 21876 16436 21882 16448
rect 22281 16439 22339 16445
rect 22281 16436 22293 16439
rect 21876 16408 22293 16436
rect 21876 16396 21882 16408
rect 22281 16405 22293 16408
rect 22327 16405 22339 16439
rect 22281 16399 22339 16405
rect 1104 16346 28888 16368
rect 1104 16294 5982 16346
rect 6034 16294 6046 16346
rect 6098 16294 6110 16346
rect 6162 16294 6174 16346
rect 6226 16294 15982 16346
rect 16034 16294 16046 16346
rect 16098 16294 16110 16346
rect 16162 16294 16174 16346
rect 16226 16294 25982 16346
rect 26034 16294 26046 16346
rect 26098 16294 26110 16346
rect 26162 16294 26174 16346
rect 26226 16294 28888 16346
rect 1104 16272 28888 16294
rect 3234 16192 3240 16244
rect 3292 16232 3298 16244
rect 3881 16235 3939 16241
rect 3881 16232 3893 16235
rect 3292 16204 3893 16232
rect 3292 16192 3298 16204
rect 3881 16201 3893 16204
rect 3927 16201 3939 16235
rect 3881 16195 3939 16201
rect 5353 16235 5411 16241
rect 5353 16201 5365 16235
rect 5399 16232 5411 16235
rect 5810 16232 5816 16244
rect 5399 16204 5816 16232
rect 5399 16201 5411 16204
rect 5353 16195 5411 16201
rect 5810 16192 5816 16204
rect 5868 16232 5874 16244
rect 7009 16235 7067 16241
rect 7009 16232 7021 16235
rect 5868 16204 7021 16232
rect 5868 16192 5874 16204
rect 7009 16201 7021 16204
rect 7055 16232 7067 16235
rect 7098 16232 7104 16244
rect 7055 16204 7104 16232
rect 7055 16201 7067 16204
rect 7009 16195 7067 16201
rect 7098 16192 7104 16204
rect 7156 16192 7162 16244
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 11149 16235 11207 16241
rect 11149 16232 11161 16235
rect 11112 16204 11161 16232
rect 11112 16192 11118 16204
rect 11149 16201 11161 16204
rect 11195 16201 11207 16235
rect 11149 16195 11207 16201
rect 15381 16235 15439 16241
rect 15381 16201 15393 16235
rect 15427 16232 15439 16235
rect 15470 16232 15476 16244
rect 15427 16204 15476 16232
rect 15427 16201 15439 16204
rect 15381 16195 15439 16201
rect 15470 16192 15476 16204
rect 15528 16232 15534 16244
rect 15746 16232 15752 16244
rect 15528 16204 15752 16232
rect 15528 16192 15534 16204
rect 15746 16192 15752 16204
rect 15804 16192 15810 16244
rect 15838 16192 15844 16244
rect 15896 16232 15902 16244
rect 16025 16235 16083 16241
rect 16025 16232 16037 16235
rect 15896 16204 16037 16232
rect 15896 16192 15902 16204
rect 16025 16201 16037 16204
rect 16071 16201 16083 16235
rect 17862 16232 17868 16244
rect 17823 16204 17868 16232
rect 16025 16195 16083 16201
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 18690 16232 18696 16244
rect 18651 16204 18696 16232
rect 18690 16192 18696 16204
rect 18748 16192 18754 16244
rect 20990 16232 20996 16244
rect 20951 16204 20996 16232
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 23934 16232 23940 16244
rect 23895 16204 23940 16232
rect 23934 16192 23940 16204
rect 23992 16192 23998 16244
rect 24854 16232 24860 16244
rect 24596 16204 24860 16232
rect 2777 16167 2835 16173
rect 2777 16133 2789 16167
rect 2823 16133 2835 16167
rect 5718 16164 5724 16176
rect 5679 16136 5724 16164
rect 2777 16127 2835 16133
rect 2792 16096 2820 16127
rect 5718 16124 5724 16136
rect 5776 16124 5782 16176
rect 6914 16124 6920 16176
rect 6972 16164 6978 16176
rect 7377 16167 7435 16173
rect 7377 16164 7389 16167
rect 6972 16136 7389 16164
rect 6972 16124 6978 16136
rect 7377 16133 7389 16136
rect 7423 16133 7435 16167
rect 7377 16127 7435 16133
rect 10229 16167 10287 16173
rect 10229 16133 10241 16167
rect 10275 16164 10287 16167
rect 11330 16164 11336 16176
rect 10275 16136 11336 16164
rect 10275 16133 10287 16136
rect 10229 16127 10287 16133
rect 11330 16124 11336 16136
rect 11388 16124 11394 16176
rect 15654 16164 15660 16176
rect 15615 16136 15660 16164
rect 15654 16124 15660 16136
rect 15712 16124 15718 16176
rect 18325 16167 18383 16173
rect 18325 16133 18337 16167
rect 18371 16164 18383 16167
rect 18782 16164 18788 16176
rect 18371 16136 18788 16164
rect 18371 16133 18383 16136
rect 18325 16127 18383 16133
rect 18782 16124 18788 16136
rect 18840 16124 18846 16176
rect 19061 16167 19119 16173
rect 19061 16133 19073 16167
rect 19107 16164 19119 16167
rect 19107 16136 19748 16164
rect 19107 16133 19119 16136
rect 19061 16127 19119 16133
rect 3050 16096 3056 16108
rect 2792 16068 3056 16096
rect 3050 16056 3056 16068
rect 3108 16096 3114 16108
rect 3421 16099 3479 16105
rect 3421 16096 3433 16099
rect 3108 16068 3433 16096
rect 3108 16056 3114 16068
rect 3421 16065 3433 16068
rect 3467 16096 3479 16099
rect 4525 16099 4583 16105
rect 4525 16096 4537 16099
rect 3467 16068 4537 16096
rect 3467 16065 3479 16068
rect 3421 16059 3479 16065
rect 4525 16065 4537 16068
rect 4571 16096 4583 16099
rect 4798 16096 4804 16108
rect 4571 16068 4804 16096
rect 4571 16065 4583 16068
rect 4525 16059 4583 16065
rect 4798 16056 4804 16068
rect 4856 16056 4862 16108
rect 5626 16056 5632 16108
rect 5684 16096 5690 16108
rect 5997 16099 6055 16105
rect 5997 16096 6009 16099
rect 5684 16068 6009 16096
rect 5684 16056 5690 16068
rect 5997 16065 6009 16068
rect 6043 16065 6055 16099
rect 5997 16059 6055 16065
rect 19150 16056 19156 16108
rect 19208 16096 19214 16108
rect 19720 16105 19748 16136
rect 20714 16124 20720 16176
rect 20772 16164 20778 16176
rect 21269 16167 21327 16173
rect 21269 16164 21281 16167
rect 20772 16136 21281 16164
rect 20772 16124 20778 16136
rect 21269 16133 21281 16136
rect 21315 16164 21327 16167
rect 21726 16164 21732 16176
rect 21315 16136 21732 16164
rect 21315 16133 21327 16136
rect 21269 16127 21327 16133
rect 21726 16124 21732 16136
rect 21784 16124 21790 16176
rect 19613 16099 19671 16105
rect 19613 16096 19625 16099
rect 19208 16068 19625 16096
rect 19208 16056 19214 16068
rect 19613 16065 19625 16068
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 19705 16099 19763 16105
rect 19705 16065 19717 16099
rect 19751 16096 19763 16099
rect 21818 16096 21824 16108
rect 19751 16068 21824 16096
rect 19751 16065 19763 16068
rect 19705 16059 19763 16065
rect 21818 16056 21824 16068
rect 21876 16056 21882 16108
rect 24596 16105 24624 16204
rect 24854 16192 24860 16204
rect 24912 16232 24918 16244
rect 25041 16235 25099 16241
rect 25041 16232 25053 16235
rect 24912 16204 25053 16232
rect 24912 16192 24918 16204
rect 25041 16201 25053 16204
rect 25087 16232 25099 16235
rect 27249 16235 27307 16241
rect 27249 16232 27261 16235
rect 25087 16204 27261 16232
rect 25087 16201 25099 16204
rect 25041 16195 25099 16201
rect 27249 16201 27261 16204
rect 27295 16201 27307 16235
rect 27249 16195 27307 16201
rect 24581 16099 24639 16105
rect 24581 16065 24593 16099
rect 24627 16065 24639 16099
rect 24581 16059 24639 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1486 16028 1492 16040
rect 1443 16000 1492 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1486 15988 1492 16000
rect 1544 15988 1550 16040
rect 8846 16028 8852 16040
rect 8807 16000 8852 16028
rect 8846 15988 8852 16000
rect 8904 15988 8910 16040
rect 19334 15988 19340 16040
rect 19392 16028 19398 16040
rect 19521 16031 19579 16037
rect 19521 16028 19533 16031
rect 19392 16000 19533 16028
rect 19392 15988 19398 16000
rect 19521 15997 19533 16000
rect 19567 15997 19579 16031
rect 23106 16028 23112 16040
rect 23019 16000 23112 16028
rect 19521 15991 19579 15997
rect 23106 15988 23112 16000
rect 23164 16028 23170 16040
rect 24305 16031 24363 16037
rect 24305 16028 24317 16031
rect 23164 16000 24317 16028
rect 23164 15988 23170 16000
rect 24305 15997 24317 16000
rect 24351 16028 24363 16031
rect 24394 16028 24400 16040
rect 24351 16000 24400 16028
rect 24351 15997 24363 16000
rect 24305 15991 24363 15997
rect 24394 15988 24400 16000
rect 24452 15988 24458 16040
rect 25869 16031 25927 16037
rect 25869 15997 25881 16031
rect 25915 16028 25927 16031
rect 25958 16028 25964 16040
rect 25915 16000 25964 16028
rect 25915 15997 25927 16000
rect 25869 15991 25927 15997
rect 25958 15988 25964 16000
rect 26016 15988 26022 16040
rect 1670 15969 1676 15972
rect 1664 15960 1676 15969
rect 1631 15932 1676 15960
rect 1664 15923 1676 15932
rect 1670 15920 1676 15923
rect 1728 15920 1734 15972
rect 3602 15920 3608 15972
rect 3660 15960 3666 15972
rect 3789 15963 3847 15969
rect 3789 15960 3801 15963
rect 3660 15932 3801 15960
rect 3660 15920 3666 15932
rect 3789 15929 3801 15932
rect 3835 15960 3847 15963
rect 4246 15960 4252 15972
rect 3835 15932 4252 15960
rect 3835 15929 3847 15932
rect 3789 15923 3847 15929
rect 4246 15920 4252 15932
rect 4304 15920 4310 15972
rect 8757 15963 8815 15969
rect 8757 15929 8769 15963
rect 8803 15960 8815 15963
rect 9030 15960 9036 15972
rect 8803 15932 9036 15960
rect 8803 15929 8815 15932
rect 8757 15923 8815 15929
rect 9030 15920 9036 15932
rect 9088 15969 9094 15972
rect 9088 15963 9152 15969
rect 9088 15929 9106 15963
rect 9140 15929 9152 15963
rect 9088 15923 9152 15929
rect 10873 15963 10931 15969
rect 10873 15929 10885 15963
rect 10919 15960 10931 15963
rect 10962 15960 10968 15972
rect 10919 15932 10968 15960
rect 10919 15929 10931 15932
rect 10873 15923 10931 15929
rect 9088 15920 9094 15923
rect 10962 15920 10968 15932
rect 11020 15920 11026 15972
rect 26114 15963 26172 15969
rect 26114 15960 26126 15963
rect 25700 15932 26126 15960
rect 4062 15852 4068 15904
rect 4120 15892 4126 15904
rect 4341 15895 4399 15901
rect 4341 15892 4353 15895
rect 4120 15864 4353 15892
rect 4120 15852 4126 15864
rect 4341 15861 4353 15864
rect 4387 15892 4399 15895
rect 4893 15895 4951 15901
rect 4893 15892 4905 15895
rect 4387 15864 4905 15892
rect 4387 15861 4399 15864
rect 4341 15855 4399 15861
rect 4893 15861 4905 15864
rect 4939 15861 4951 15895
rect 4893 15855 4951 15861
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 12621 15895 12679 15901
rect 12621 15892 12633 15895
rect 12492 15864 12633 15892
rect 12492 15852 12498 15864
rect 12621 15861 12633 15864
rect 12667 15861 12679 15895
rect 12986 15892 12992 15904
rect 12947 15864 12992 15892
rect 12621 15855 12679 15861
rect 12986 15852 12992 15864
rect 13044 15852 13050 15904
rect 19058 15852 19064 15904
rect 19116 15892 19122 15904
rect 19153 15895 19211 15901
rect 19153 15892 19165 15895
rect 19116 15864 19165 15892
rect 19116 15852 19122 15864
rect 19153 15861 19165 15864
rect 19199 15861 19211 15895
rect 19153 15855 19211 15861
rect 23477 15895 23535 15901
rect 23477 15861 23489 15895
rect 23523 15892 23535 15895
rect 23934 15892 23940 15904
rect 23523 15864 23940 15892
rect 23523 15861 23535 15864
rect 23477 15855 23535 15861
rect 23934 15852 23940 15864
rect 23992 15892 23998 15904
rect 24397 15895 24455 15901
rect 24397 15892 24409 15895
rect 23992 15864 24409 15892
rect 23992 15852 23998 15864
rect 24397 15861 24409 15864
rect 24443 15861 24455 15895
rect 24397 15855 24455 15861
rect 25222 15852 25228 15904
rect 25280 15892 25286 15904
rect 25700 15901 25728 15932
rect 26114 15929 26126 15932
rect 26160 15929 26172 15963
rect 26114 15923 26172 15929
rect 25685 15895 25743 15901
rect 25685 15892 25697 15895
rect 25280 15864 25697 15892
rect 25280 15852 25286 15864
rect 25685 15861 25697 15864
rect 25731 15861 25743 15895
rect 25685 15855 25743 15861
rect 1104 15802 28888 15824
rect 1104 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 20982 15802
rect 21034 15750 21046 15802
rect 21098 15750 21110 15802
rect 21162 15750 21174 15802
rect 21226 15750 28888 15802
rect 1104 15728 28888 15750
rect 1486 15648 1492 15700
rect 1544 15688 1550 15700
rect 1762 15688 1768 15700
rect 1544 15660 1768 15688
rect 1544 15648 1550 15660
rect 1762 15648 1768 15660
rect 1820 15688 1826 15700
rect 1949 15691 2007 15697
rect 1949 15688 1961 15691
rect 1820 15660 1961 15688
rect 1820 15648 1826 15660
rect 1949 15657 1961 15660
rect 1995 15657 2007 15691
rect 1949 15651 2007 15657
rect 2501 15691 2559 15697
rect 2501 15657 2513 15691
rect 2547 15688 2559 15691
rect 2682 15688 2688 15700
rect 2547 15660 2688 15688
rect 2547 15657 2559 15660
rect 2501 15651 2559 15657
rect 2682 15648 2688 15660
rect 2740 15648 2746 15700
rect 2866 15688 2872 15700
rect 2827 15660 2872 15688
rect 2866 15648 2872 15660
rect 2924 15648 2930 15700
rect 4062 15688 4068 15700
rect 4023 15660 4068 15688
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 10413 15691 10471 15697
rect 10413 15657 10425 15691
rect 10459 15688 10471 15691
rect 10870 15688 10876 15700
rect 10459 15660 10876 15688
rect 10459 15657 10471 15660
rect 10413 15651 10471 15657
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 16298 15688 16304 15700
rect 15304 15660 16304 15688
rect 4430 15620 4436 15632
rect 4391 15592 4436 15620
rect 4430 15580 4436 15592
rect 4488 15580 4494 15632
rect 11330 15580 11336 15632
rect 11388 15620 11394 15632
rect 11578 15623 11636 15629
rect 11578 15620 11590 15623
rect 11388 15592 11590 15620
rect 11388 15580 11394 15592
rect 11578 15589 11590 15592
rect 11624 15589 11636 15623
rect 11578 15583 11636 15589
rect 15304 15564 15332 15660
rect 16298 15648 16304 15660
rect 16356 15688 16362 15700
rect 17773 15691 17831 15697
rect 17773 15688 17785 15691
rect 16356 15660 17785 15688
rect 16356 15648 16362 15660
rect 17773 15657 17785 15660
rect 17819 15657 17831 15691
rect 17773 15651 17831 15657
rect 18049 15691 18107 15697
rect 18049 15657 18061 15691
rect 18095 15688 18107 15691
rect 18690 15688 18696 15700
rect 18095 15660 18696 15688
rect 18095 15657 18107 15660
rect 18049 15651 18107 15657
rect 18690 15648 18696 15660
rect 18748 15648 18754 15700
rect 19150 15688 19156 15700
rect 19111 15660 19156 15688
rect 19150 15648 19156 15660
rect 19208 15648 19214 15700
rect 24121 15691 24179 15697
rect 24121 15657 24133 15691
rect 24167 15688 24179 15691
rect 24486 15688 24492 15700
rect 24167 15660 24492 15688
rect 24167 15657 24179 15660
rect 24121 15651 24179 15657
rect 24486 15648 24492 15660
rect 24544 15648 24550 15700
rect 24854 15688 24860 15700
rect 24815 15660 24860 15688
rect 24854 15648 24860 15660
rect 24912 15648 24918 15700
rect 25958 15688 25964 15700
rect 25919 15660 25964 15688
rect 25958 15648 25964 15660
rect 26016 15648 26022 15700
rect 21818 15580 21824 15632
rect 21876 15620 21882 15632
rect 21974 15623 22032 15629
rect 21974 15620 21986 15623
rect 21876 15592 21986 15620
rect 21876 15580 21882 15592
rect 21974 15589 21986 15592
rect 22020 15589 22032 15623
rect 21974 15583 22032 15589
rect 8294 15512 8300 15564
rect 8352 15552 8358 15564
rect 9401 15555 9459 15561
rect 9401 15552 9413 15555
rect 8352 15524 9413 15552
rect 8352 15512 8358 15524
rect 9401 15521 9413 15524
rect 9447 15552 9459 15555
rect 9582 15552 9588 15564
rect 9447 15524 9588 15552
rect 9447 15521 9459 15524
rect 9401 15515 9459 15521
rect 9582 15512 9588 15524
rect 9640 15512 9646 15564
rect 15286 15552 15292 15564
rect 15199 15524 15292 15552
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 15378 15512 15384 15564
rect 15436 15552 15442 15564
rect 15545 15555 15603 15561
rect 15545 15552 15557 15555
rect 15436 15524 15557 15552
rect 15436 15512 15442 15524
rect 15545 15521 15557 15524
rect 15591 15521 15603 15555
rect 17954 15552 17960 15564
rect 17915 15524 17960 15552
rect 15545 15515 15603 15521
rect 17954 15512 17960 15524
rect 18012 15512 18018 15564
rect 18414 15552 18420 15564
rect 18375 15524 18420 15552
rect 18414 15512 18420 15524
rect 18472 15512 18478 15564
rect 21726 15552 21732 15564
rect 21687 15524 21732 15552
rect 21726 15512 21732 15524
rect 21784 15512 21790 15564
rect 26510 15552 26516 15564
rect 26471 15524 26516 15552
rect 26510 15512 26516 15524
rect 26568 15512 26574 15564
rect 4522 15484 4528 15496
rect 4483 15456 4528 15484
rect 4522 15444 4528 15456
rect 4580 15444 4586 15496
rect 4709 15487 4767 15493
rect 4709 15453 4721 15487
rect 4755 15484 4767 15487
rect 4890 15484 4896 15496
rect 4755 15456 4896 15484
rect 4755 15453 4767 15456
rect 4709 15447 4767 15453
rect 1670 15416 1676 15428
rect 1583 15388 1676 15416
rect 1670 15376 1676 15388
rect 1728 15416 1734 15428
rect 4724 15416 4752 15447
rect 4890 15444 4896 15456
rect 4948 15444 4954 15496
rect 11238 15484 11244 15496
rect 9232 15456 11244 15484
rect 1728 15388 4752 15416
rect 1728 15376 1734 15388
rect 7650 15308 7656 15360
rect 7708 15348 7714 15360
rect 7745 15351 7803 15357
rect 7745 15348 7757 15351
rect 7708 15320 7757 15348
rect 7708 15308 7714 15320
rect 7745 15317 7757 15320
rect 7791 15348 7803 15351
rect 8478 15348 8484 15360
rect 7791 15320 8484 15348
rect 7791 15317 7803 15320
rect 7745 15311 7803 15317
rect 8478 15308 8484 15320
rect 8536 15348 8542 15360
rect 8846 15348 8852 15360
rect 8536 15320 8852 15348
rect 8536 15308 8542 15320
rect 8846 15308 8852 15320
rect 8904 15348 8910 15360
rect 9232 15357 9260 15456
rect 11238 15444 11244 15456
rect 11296 15484 11302 15496
rect 11333 15487 11391 15493
rect 11333 15484 11345 15487
rect 11296 15456 11345 15484
rect 11296 15444 11302 15456
rect 11333 15453 11345 15456
rect 11379 15453 11391 15487
rect 18506 15484 18512 15496
rect 18467 15456 18512 15484
rect 11333 15447 11391 15453
rect 18506 15444 18512 15456
rect 18564 15444 18570 15496
rect 18601 15487 18659 15493
rect 18601 15453 18613 15487
rect 18647 15453 18659 15487
rect 18601 15447 18659 15453
rect 18046 15376 18052 15428
rect 18104 15416 18110 15428
rect 18616 15416 18644 15447
rect 18874 15416 18880 15428
rect 18104 15388 18880 15416
rect 18104 15376 18110 15388
rect 18874 15376 18880 15388
rect 18932 15416 18938 15428
rect 19242 15416 19248 15428
rect 18932 15388 19248 15416
rect 18932 15376 18938 15388
rect 19242 15376 19248 15388
rect 19300 15376 19306 15428
rect 9217 15351 9275 15357
rect 9217 15348 9229 15351
rect 8904 15320 9229 15348
rect 8904 15308 8910 15320
rect 9217 15317 9229 15320
rect 9263 15317 9275 15351
rect 9217 15311 9275 15317
rect 12434 15308 12440 15360
rect 12492 15348 12498 15360
rect 12713 15351 12771 15357
rect 12713 15348 12725 15351
rect 12492 15320 12725 15348
rect 12492 15308 12498 15320
rect 12713 15317 12725 15320
rect 12759 15317 12771 15351
rect 16666 15348 16672 15360
rect 16627 15320 16672 15348
rect 12713 15311 12771 15317
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 23106 15348 23112 15360
rect 23067 15320 23112 15348
rect 23106 15308 23112 15320
rect 23164 15308 23170 15360
rect 24302 15308 24308 15360
rect 24360 15348 24366 15360
rect 24489 15351 24547 15357
rect 24489 15348 24501 15351
rect 24360 15320 24501 15348
rect 24360 15308 24366 15320
rect 24489 15317 24501 15320
rect 24535 15348 24547 15351
rect 24762 15348 24768 15360
rect 24535 15320 24768 15348
rect 24535 15317 24547 15320
rect 24489 15311 24547 15317
rect 24762 15308 24768 15320
rect 24820 15308 24826 15360
rect 26697 15351 26755 15357
rect 26697 15317 26709 15351
rect 26743 15348 26755 15351
rect 27246 15348 27252 15360
rect 26743 15320 27252 15348
rect 26743 15317 26755 15320
rect 26697 15311 26755 15317
rect 27246 15308 27252 15320
rect 27304 15308 27310 15360
rect 1104 15258 28888 15280
rect 1104 15206 5982 15258
rect 6034 15206 6046 15258
rect 6098 15206 6110 15258
rect 6162 15206 6174 15258
rect 6226 15206 15982 15258
rect 16034 15206 16046 15258
rect 16098 15206 16110 15258
rect 16162 15206 16174 15258
rect 16226 15206 25982 15258
rect 26034 15206 26046 15258
rect 26098 15206 26110 15258
rect 26162 15206 26174 15258
rect 26226 15206 28888 15258
rect 1104 15184 28888 15206
rect 1394 15104 1400 15156
rect 1452 15144 1458 15156
rect 1673 15147 1731 15153
rect 1673 15144 1685 15147
rect 1452 15116 1685 15144
rect 1452 15104 1458 15116
rect 1673 15113 1685 15116
rect 1719 15144 1731 15147
rect 1762 15144 1768 15156
rect 1719 15116 1768 15144
rect 1719 15113 1731 15116
rect 1673 15107 1731 15113
rect 1762 15104 1768 15116
rect 1820 15104 1826 15156
rect 4430 15144 4436 15156
rect 4391 15116 4436 15144
rect 4430 15104 4436 15116
rect 4488 15104 4494 15156
rect 5166 15104 5172 15156
rect 5224 15144 5230 15156
rect 6457 15147 6515 15153
rect 6457 15144 6469 15147
rect 5224 15116 6469 15144
rect 5224 15104 5230 15116
rect 6457 15113 6469 15116
rect 6503 15144 6515 15147
rect 6822 15144 6828 15156
rect 6503 15116 6828 15144
rect 6503 15113 6515 15116
rect 6457 15107 6515 15113
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 7101 15147 7159 15153
rect 7101 15113 7113 15147
rect 7147 15144 7159 15147
rect 7926 15144 7932 15156
rect 7147 15116 7932 15144
rect 7147 15113 7159 15116
rect 7101 15107 7159 15113
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14940 6699 14943
rect 7116 14940 7144 15107
rect 7926 15104 7932 15116
rect 7984 15144 7990 15156
rect 8294 15144 8300 15156
rect 7984 15116 8300 15144
rect 7984 15104 7990 15116
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 9030 15144 9036 15156
rect 8991 15116 9036 15144
rect 9030 15104 9036 15116
rect 9088 15104 9094 15156
rect 9674 15144 9680 15156
rect 9635 15116 9680 15144
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 11238 15104 11244 15156
rect 11296 15144 11302 15156
rect 11701 15147 11759 15153
rect 11701 15144 11713 15147
rect 11296 15116 11713 15144
rect 11296 15104 11302 15116
rect 11701 15113 11713 15116
rect 11747 15144 11759 15147
rect 12342 15144 12348 15156
rect 11747 15116 12348 15144
rect 11747 15113 11759 15116
rect 11701 15107 11759 15113
rect 12342 15104 12348 15116
rect 12400 15144 12406 15156
rect 12986 15144 12992 15156
rect 12400 15116 12992 15144
rect 12400 15104 12406 15116
rect 12986 15104 12992 15116
rect 13044 15104 13050 15156
rect 15378 15144 15384 15156
rect 15339 15116 15384 15144
rect 15378 15104 15384 15116
rect 15436 15104 15442 15156
rect 15749 15147 15807 15153
rect 15749 15113 15761 15147
rect 15795 15144 15807 15147
rect 16298 15144 16304 15156
rect 15795 15116 16304 15144
rect 15795 15113 15807 15116
rect 15749 15107 15807 15113
rect 16298 15104 16304 15116
rect 16356 15104 16362 15156
rect 17497 15147 17555 15153
rect 17497 15113 17509 15147
rect 17543 15144 17555 15147
rect 17954 15144 17960 15156
rect 17543 15116 17960 15144
rect 17543 15113 17555 15116
rect 17497 15107 17555 15113
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 18325 15147 18383 15153
rect 18325 15113 18337 15147
rect 18371 15144 18383 15147
rect 18414 15144 18420 15156
rect 18371 15116 18420 15144
rect 18371 15113 18383 15116
rect 18325 15107 18383 15113
rect 18414 15104 18420 15116
rect 18472 15104 18478 15156
rect 19334 15104 19340 15156
rect 19392 15144 19398 15156
rect 20349 15147 20407 15153
rect 20349 15144 20361 15147
rect 19392 15116 20361 15144
rect 19392 15104 19398 15116
rect 20349 15113 20361 15116
rect 20395 15113 20407 15147
rect 20349 15107 20407 15113
rect 21361 15147 21419 15153
rect 21361 15113 21373 15147
rect 21407 15144 21419 15147
rect 21453 15147 21511 15153
rect 21453 15144 21465 15147
rect 21407 15116 21465 15144
rect 21407 15113 21419 15116
rect 21361 15107 21419 15113
rect 21453 15113 21465 15116
rect 21499 15144 21511 15147
rect 21726 15144 21732 15156
rect 21499 15116 21732 15144
rect 21499 15113 21511 15116
rect 21453 15107 21511 15113
rect 21726 15104 21732 15116
rect 21784 15104 21790 15156
rect 21818 15104 21824 15156
rect 21876 15144 21882 15156
rect 21913 15147 21971 15153
rect 21913 15144 21925 15147
rect 21876 15116 21925 15144
rect 21876 15104 21882 15116
rect 21913 15113 21925 15116
rect 21959 15113 21971 15147
rect 26510 15144 26516 15156
rect 26471 15116 26516 15144
rect 21913 15107 21971 15113
rect 26510 15104 26516 15116
rect 26568 15104 26574 15156
rect 17865 15079 17923 15085
rect 17865 15045 17877 15079
rect 17911 15076 17923 15079
rect 18046 15076 18052 15088
rect 17911 15048 18052 15076
rect 17911 15045 17923 15048
rect 17865 15039 17923 15045
rect 18046 15036 18052 15048
rect 18104 15036 18110 15088
rect 7650 15008 7656 15020
rect 7611 14980 7656 15008
rect 7650 14968 7656 14980
rect 7708 14968 7714 15020
rect 24489 15011 24547 15017
rect 24489 14977 24501 15011
rect 24535 15008 24547 15011
rect 25222 15008 25228 15020
rect 24535 14980 25228 15008
rect 24535 14977 24547 14980
rect 24489 14971 24547 14977
rect 25222 14968 25228 14980
rect 25280 14968 25286 15020
rect 7920 14943 7978 14949
rect 7920 14940 7932 14943
rect 6687 14912 7144 14940
rect 7852 14912 7932 14940
rect 6687 14909 6699 14912
rect 6641 14903 6699 14909
rect 7561 14875 7619 14881
rect 7561 14841 7573 14875
rect 7607 14872 7619 14875
rect 7852 14872 7880 14912
rect 7920 14909 7932 14912
rect 7966 14940 7978 14943
rect 8202 14940 8208 14952
rect 7966 14912 8208 14940
rect 7966 14909 7978 14912
rect 7920 14903 7978 14909
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 18966 14940 18972 14952
rect 18927 14912 18972 14940
rect 18966 14900 18972 14912
rect 19024 14900 19030 14952
rect 21637 14943 21695 14949
rect 21637 14909 21649 14943
rect 21683 14940 21695 14943
rect 22281 14943 22339 14949
rect 22281 14940 22293 14943
rect 21683 14912 22293 14940
rect 21683 14909 21695 14912
rect 21637 14903 21695 14909
rect 22281 14909 22293 14912
rect 22327 14909 22339 14943
rect 22281 14903 22339 14909
rect 19214 14875 19272 14881
rect 19214 14872 19226 14875
rect 7607 14844 7880 14872
rect 18892 14844 19226 14872
rect 7607 14841 7619 14844
rect 7561 14835 7619 14841
rect 18892 14816 18920 14844
rect 19214 14841 19226 14844
rect 19260 14841 19272 14875
rect 19214 14835 19272 14841
rect 19886 14832 19892 14884
rect 19944 14872 19950 14884
rect 21652 14872 21680 14903
rect 19944 14844 21680 14872
rect 24121 14875 24179 14881
rect 19944 14832 19950 14844
rect 24121 14841 24133 14875
rect 24167 14872 24179 14875
rect 24949 14875 25007 14881
rect 24949 14872 24961 14875
rect 24167 14844 24961 14872
rect 24167 14841 24179 14844
rect 24121 14835 24179 14841
rect 24949 14841 24961 14844
rect 24995 14872 25007 14875
rect 26142 14872 26148 14884
rect 24995 14844 26148 14872
rect 24995 14841 25007 14844
rect 24949 14835 25007 14841
rect 26142 14832 26148 14844
rect 26200 14832 26206 14884
rect 4157 14807 4215 14813
rect 4157 14773 4169 14807
rect 4203 14804 4215 14807
rect 4522 14804 4528 14816
rect 4203 14776 4528 14804
rect 4203 14773 4215 14776
rect 4157 14767 4215 14773
rect 4522 14764 4528 14776
rect 4580 14764 4586 14816
rect 4890 14804 4896 14816
rect 4851 14776 4896 14804
rect 4890 14764 4896 14776
rect 4948 14764 4954 14816
rect 11330 14804 11336 14816
rect 11291 14776 11336 14804
rect 11330 14764 11336 14776
rect 11388 14764 11394 14816
rect 18874 14804 18880 14816
rect 18835 14776 18880 14804
rect 18874 14764 18880 14776
rect 18932 14764 18938 14816
rect 24486 14764 24492 14816
rect 24544 14804 24550 14816
rect 24581 14807 24639 14813
rect 24581 14804 24593 14807
rect 24544 14776 24593 14804
rect 24544 14764 24550 14776
rect 24581 14773 24593 14776
rect 24627 14773 24639 14807
rect 24581 14767 24639 14773
rect 25038 14764 25044 14816
rect 25096 14804 25102 14816
rect 25096 14776 25141 14804
rect 25096 14764 25102 14776
rect 1104 14714 28888 14736
rect 1104 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 20982 14714
rect 21034 14662 21046 14714
rect 21098 14662 21110 14714
rect 21162 14662 21174 14714
rect 21226 14662 28888 14714
rect 1104 14640 28888 14662
rect 1394 14560 1400 14612
rect 1452 14600 1458 14612
rect 1452 14572 2728 14600
rect 1452 14560 1458 14572
rect 1670 14492 1676 14544
rect 1728 14541 1734 14544
rect 1728 14535 1792 14541
rect 1728 14501 1746 14535
rect 1780 14501 1792 14535
rect 2700 14532 2728 14572
rect 4890 14560 4896 14612
rect 4948 14600 4954 14612
rect 6549 14603 6607 14609
rect 6549 14600 6561 14603
rect 4948 14572 6561 14600
rect 4948 14560 4954 14572
rect 6549 14569 6561 14572
rect 6595 14569 6607 14603
rect 6549 14563 6607 14569
rect 18141 14603 18199 14609
rect 18141 14569 18153 14603
rect 18187 14600 18199 14603
rect 18325 14603 18383 14609
rect 18325 14600 18337 14603
rect 18187 14572 18337 14600
rect 18187 14569 18199 14572
rect 18141 14563 18199 14569
rect 18325 14569 18337 14572
rect 18371 14600 18383 14603
rect 18506 14600 18512 14612
rect 18371 14572 18512 14600
rect 18371 14569 18383 14572
rect 18325 14563 18383 14569
rect 18506 14560 18512 14572
rect 18564 14560 18570 14612
rect 19886 14600 19892 14612
rect 19847 14572 19892 14600
rect 19886 14560 19892 14572
rect 19944 14560 19950 14612
rect 24673 14603 24731 14609
rect 24673 14569 24685 14603
rect 24719 14600 24731 14603
rect 25038 14600 25044 14612
rect 24719 14572 25044 14600
rect 24719 14569 24731 14572
rect 24673 14563 24731 14569
rect 25038 14560 25044 14572
rect 25096 14560 25102 14612
rect 4246 14532 4252 14544
rect 2700 14504 4252 14532
rect 1728 14495 1792 14501
rect 1728 14492 1734 14495
rect 4246 14492 4252 14504
rect 4304 14492 4310 14544
rect 11149 14535 11207 14541
rect 11149 14501 11161 14535
rect 11195 14532 11207 14535
rect 11698 14532 11704 14544
rect 11195 14504 11704 14532
rect 11195 14501 11207 14504
rect 11149 14495 11207 14501
rect 11698 14492 11704 14504
rect 11756 14492 11762 14544
rect 15378 14492 15384 14544
rect 15436 14532 15442 14544
rect 15556 14535 15614 14541
rect 15556 14532 15568 14535
rect 15436 14504 15568 14532
rect 15436 14492 15442 14504
rect 15556 14501 15568 14504
rect 15602 14532 15614 14535
rect 16666 14532 16672 14544
rect 15602 14504 16672 14532
rect 15602 14501 15614 14504
rect 15556 14495 15614 14501
rect 16666 14492 16672 14504
rect 16724 14492 16730 14544
rect 18966 14492 18972 14544
rect 19024 14532 19030 14544
rect 19429 14535 19487 14541
rect 19429 14532 19441 14535
rect 19024 14504 19441 14532
rect 19024 14492 19030 14504
rect 19429 14501 19441 14504
rect 19475 14532 19487 14535
rect 20438 14532 20444 14544
rect 19475 14504 20444 14532
rect 19475 14501 19487 14504
rect 19429 14495 19487 14501
rect 20438 14492 20444 14504
rect 20496 14532 20502 14544
rect 22097 14535 22155 14541
rect 20496 14504 21772 14532
rect 20496 14492 20502 14504
rect 21744 14476 21772 14504
rect 22097 14501 22109 14535
rect 22143 14532 22155 14535
rect 22732 14535 22790 14541
rect 22732 14532 22744 14535
rect 22143 14504 22744 14532
rect 22143 14501 22155 14504
rect 22097 14495 22155 14501
rect 22732 14501 22744 14504
rect 22778 14532 22790 14535
rect 23106 14532 23112 14544
rect 22778 14504 23112 14532
rect 22778 14501 22790 14504
rect 22732 14495 22790 14501
rect 23106 14492 23112 14504
rect 23164 14492 23170 14544
rect 24854 14492 24860 14544
rect 24912 14532 24918 14544
rect 25406 14532 25412 14544
rect 24912 14504 25412 14532
rect 24912 14492 24918 14504
rect 25406 14492 25412 14504
rect 25464 14492 25470 14544
rect 5166 14464 5172 14476
rect 5127 14436 5172 14464
rect 5166 14424 5172 14436
rect 5224 14424 5230 14476
rect 5442 14473 5448 14476
rect 5436 14427 5448 14473
rect 5500 14464 5506 14476
rect 5500 14436 5536 14464
rect 5442 14424 5448 14427
rect 5500 14424 5506 14436
rect 7834 14424 7840 14476
rect 7892 14464 7898 14476
rect 8021 14467 8079 14473
rect 8021 14464 8033 14467
rect 7892 14436 8033 14464
rect 7892 14424 7898 14436
rect 8021 14433 8033 14436
rect 8067 14433 8079 14467
rect 8021 14427 8079 14433
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 11606 14464 11612 14476
rect 11112 14436 11612 14464
rect 11112 14424 11118 14436
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 15286 14464 15292 14476
rect 15247 14436 15292 14464
rect 15286 14424 15292 14436
rect 15344 14424 15350 14476
rect 17770 14424 17776 14476
rect 17828 14464 17834 14476
rect 18690 14464 18696 14476
rect 17828 14436 18696 14464
rect 17828 14424 17834 14436
rect 18690 14424 18696 14436
rect 18748 14424 18754 14476
rect 20073 14467 20131 14473
rect 20073 14433 20085 14467
rect 20119 14464 20131 14467
rect 20530 14464 20536 14476
rect 20119 14436 20536 14464
rect 20119 14433 20131 14436
rect 20073 14427 20131 14433
rect 20530 14424 20536 14436
rect 20588 14424 20594 14476
rect 21726 14424 21732 14476
rect 21784 14464 21790 14476
rect 22465 14467 22523 14473
rect 22465 14464 22477 14467
rect 21784 14436 22477 14464
rect 21784 14424 21790 14436
rect 22465 14433 22477 14436
rect 22511 14464 22523 14467
rect 22554 14464 22560 14476
rect 22511 14436 22560 14464
rect 22511 14433 22523 14436
rect 22465 14427 22523 14433
rect 22554 14424 22560 14436
rect 22612 14424 22618 14476
rect 1394 14356 1400 14408
rect 1452 14396 1458 14408
rect 1489 14399 1547 14405
rect 1489 14396 1501 14399
rect 1452 14368 1501 14396
rect 1452 14356 1458 14368
rect 1489 14365 1501 14368
rect 1535 14365 1547 14399
rect 1489 14359 1547 14365
rect 7466 14356 7472 14408
rect 7524 14396 7530 14408
rect 8113 14399 8171 14405
rect 8113 14396 8125 14399
rect 7524 14368 8125 14396
rect 7524 14356 7530 14368
rect 8113 14365 8125 14368
rect 8159 14365 8171 14399
rect 8113 14359 8171 14365
rect 8202 14356 8208 14408
rect 8260 14396 8266 14408
rect 8260 14368 8305 14396
rect 8260 14356 8266 14368
rect 11330 14356 11336 14408
rect 11388 14396 11394 14408
rect 11793 14399 11851 14405
rect 11793 14396 11805 14399
rect 11388 14368 11805 14396
rect 11388 14356 11394 14368
rect 11793 14365 11805 14368
rect 11839 14365 11851 14399
rect 11793 14359 11851 14365
rect 12529 14399 12587 14405
rect 12529 14365 12541 14399
rect 12575 14396 12587 14399
rect 12802 14396 12808 14408
rect 12575 14368 12808 14396
rect 12575 14365 12587 14368
rect 12529 14359 12587 14365
rect 12802 14356 12808 14368
rect 12860 14356 12866 14408
rect 18506 14356 18512 14408
rect 18564 14396 18570 14408
rect 18785 14399 18843 14405
rect 18785 14396 18797 14399
rect 18564 14368 18797 14396
rect 18564 14356 18570 14368
rect 18785 14365 18797 14368
rect 18831 14365 18843 14399
rect 18785 14359 18843 14365
rect 18874 14356 18880 14408
rect 18932 14396 18938 14408
rect 18932 14368 18977 14396
rect 18932 14356 18938 14368
rect 10781 14331 10839 14337
rect 10781 14297 10793 14331
rect 10827 14328 10839 14331
rect 11146 14328 11152 14340
rect 10827 14300 11152 14328
rect 10827 14297 10839 14300
rect 10781 14291 10839 14297
rect 11146 14288 11152 14300
rect 11204 14328 11210 14340
rect 11241 14331 11299 14337
rect 11241 14328 11253 14331
rect 11204 14300 11253 14328
rect 11204 14288 11210 14300
rect 11241 14297 11253 14300
rect 11287 14297 11299 14331
rect 11241 14291 11299 14297
rect 2866 14260 2872 14272
rect 2827 14232 2872 14260
rect 2866 14220 2872 14232
rect 2924 14220 2930 14272
rect 4338 14260 4344 14272
rect 4299 14232 4344 14260
rect 4338 14220 4344 14232
rect 4396 14220 4402 14272
rect 7561 14263 7619 14269
rect 7561 14229 7573 14263
rect 7607 14260 7619 14263
rect 7653 14263 7711 14269
rect 7653 14260 7665 14263
rect 7607 14232 7665 14260
rect 7607 14229 7619 14232
rect 7561 14223 7619 14229
rect 7653 14229 7665 14232
rect 7699 14260 7711 14263
rect 8018 14260 8024 14272
rect 7699 14232 8024 14260
rect 7699 14229 7711 14232
rect 7653 14223 7711 14229
rect 8018 14220 8024 14232
rect 8076 14220 8082 14272
rect 9214 14260 9220 14272
rect 9175 14232 9220 14260
rect 9214 14220 9220 14232
rect 9272 14220 9278 14272
rect 14274 14260 14280 14272
rect 14235 14232 14280 14260
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 16666 14260 16672 14272
rect 16627 14232 16672 14260
rect 16666 14220 16672 14232
rect 16724 14220 16730 14272
rect 23842 14260 23848 14272
rect 23803 14232 23848 14260
rect 23842 14220 23848 14232
rect 23900 14220 23906 14272
rect 1104 14170 28888 14192
rect 1104 14118 5982 14170
rect 6034 14118 6046 14170
rect 6098 14118 6110 14170
rect 6162 14118 6174 14170
rect 6226 14118 15982 14170
rect 16034 14118 16046 14170
rect 16098 14118 16110 14170
rect 16162 14118 16174 14170
rect 16226 14118 25982 14170
rect 26034 14118 26046 14170
rect 26098 14118 26110 14170
rect 26162 14118 26174 14170
rect 26226 14118 28888 14170
rect 1104 14096 28888 14118
rect 4062 14056 4068 14068
rect 4023 14028 4068 14056
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 4246 14016 4252 14068
rect 4304 14056 4310 14068
rect 5166 14056 5172 14068
rect 4304 14028 5172 14056
rect 4304 14016 4310 14028
rect 5166 14016 5172 14028
rect 5224 14056 5230 14068
rect 5629 14059 5687 14065
rect 5629 14056 5641 14059
rect 5224 14028 5641 14056
rect 5224 14016 5230 14028
rect 5629 14025 5641 14028
rect 5675 14025 5687 14059
rect 5629 14019 5687 14025
rect 8389 14059 8447 14065
rect 8389 14025 8401 14059
rect 8435 14056 8447 14059
rect 8665 14059 8723 14065
rect 8665 14056 8677 14059
rect 8435 14028 8677 14056
rect 8435 14025 8447 14028
rect 8389 14019 8447 14025
rect 8665 14025 8677 14028
rect 8711 14056 8723 14059
rect 8938 14056 8944 14068
rect 8711 14028 8944 14056
rect 8711 14025 8723 14028
rect 8665 14019 8723 14025
rect 8938 14016 8944 14028
rect 8996 14056 9002 14068
rect 9582 14056 9588 14068
rect 8996 14028 9588 14056
rect 8996 14016 9002 14028
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 10689 14059 10747 14065
rect 10689 14025 10701 14059
rect 10735 14056 10747 14059
rect 10735 14028 11468 14056
rect 10735 14025 10747 14028
rect 10689 14019 10747 14025
rect 5353 13991 5411 13997
rect 5353 13957 5365 13991
rect 5399 13988 5411 13991
rect 5442 13988 5448 14000
rect 5399 13960 5448 13988
rect 5399 13957 5411 13960
rect 5353 13951 5411 13957
rect 5442 13948 5448 13960
rect 5500 13948 5506 14000
rect 7561 13991 7619 13997
rect 7561 13957 7573 13991
rect 7607 13988 7619 13991
rect 9030 13988 9036 14000
rect 7607 13960 9036 13988
rect 7607 13957 7619 13960
rect 7561 13951 7619 13957
rect 9030 13948 9036 13960
rect 9088 13948 9094 14000
rect 9125 13991 9183 13997
rect 9125 13957 9137 13991
rect 9171 13988 9183 13991
rect 10229 13991 10287 13997
rect 10229 13988 10241 13991
rect 9171 13960 10241 13988
rect 9171 13957 9183 13960
rect 9125 13951 9183 13957
rect 10229 13957 10241 13960
rect 10275 13988 10287 13991
rect 10275 13960 11284 13988
rect 10275 13957 10287 13960
rect 10229 13951 10287 13957
rect 2314 13880 2320 13932
rect 2372 13920 2378 13932
rect 3237 13923 3295 13929
rect 3237 13920 3249 13923
rect 2372 13892 3249 13920
rect 2372 13880 2378 13892
rect 3237 13889 3249 13892
rect 3283 13920 3295 13923
rect 3510 13920 3516 13932
rect 3283 13892 3516 13920
rect 3283 13889 3295 13892
rect 3237 13883 3295 13889
rect 3510 13880 3516 13892
rect 3568 13920 3574 13932
rect 3789 13923 3847 13929
rect 3789 13920 3801 13923
rect 3568 13892 3801 13920
rect 3568 13880 3574 13892
rect 3789 13889 3801 13892
rect 3835 13920 3847 13923
rect 4798 13920 4804 13932
rect 3835 13892 4804 13920
rect 3835 13889 3847 13892
rect 3789 13883 3847 13889
rect 4798 13880 4804 13892
rect 4856 13880 4862 13932
rect 7466 13920 7472 13932
rect 7427 13892 7472 13920
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 8018 13920 8024 13932
rect 7979 13892 8024 13920
rect 8018 13880 8024 13892
rect 8076 13880 8082 13932
rect 8205 13923 8263 13929
rect 8205 13889 8217 13923
rect 8251 13920 8263 13923
rect 8389 13923 8447 13929
rect 8389 13920 8401 13923
rect 8251 13892 8401 13920
rect 8251 13889 8263 13892
rect 8205 13883 8263 13889
rect 8389 13889 8401 13892
rect 8435 13889 8447 13923
rect 9048 13920 9076 13948
rect 9585 13923 9643 13929
rect 9585 13920 9597 13923
rect 9048 13892 9597 13920
rect 8389 13883 8447 13889
rect 9585 13889 9597 13892
rect 9631 13889 9643 13923
rect 9585 13883 9643 13889
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 11256 13929 11284 13960
rect 11440 13929 11468 14028
rect 11606 14016 11612 14068
rect 11664 14056 11670 14068
rect 12437 14059 12495 14065
rect 12437 14056 12449 14059
rect 11664 14028 12449 14056
rect 11664 14016 11670 14028
rect 12437 14025 12449 14028
rect 12483 14025 12495 14059
rect 15378 14056 15384 14068
rect 15339 14028 15384 14056
rect 12437 14019 12495 14025
rect 15378 14016 15384 14028
rect 15436 14016 15442 14068
rect 16758 14016 16764 14068
rect 16816 14056 16822 14068
rect 17770 14056 17776 14068
rect 16816 14028 17776 14056
rect 16816 14016 16822 14028
rect 17770 14016 17776 14028
rect 17828 14016 17834 14068
rect 18874 14016 18880 14068
rect 18932 14056 18938 14068
rect 19613 14059 19671 14065
rect 19613 14056 19625 14059
rect 18932 14028 19625 14056
rect 18932 14016 18938 14028
rect 19613 14025 19625 14028
rect 19659 14025 19671 14059
rect 19613 14019 19671 14025
rect 20714 14016 20720 14068
rect 20772 14056 20778 14068
rect 21913 14059 21971 14065
rect 21913 14056 21925 14059
rect 20772 14028 21925 14056
rect 20772 14016 20778 14028
rect 21913 14025 21925 14028
rect 21959 14056 21971 14059
rect 23106 14056 23112 14068
rect 21959 14028 22508 14056
rect 23067 14028 23112 14056
rect 21959 14025 21971 14028
rect 21913 14019 21971 14025
rect 12253 13991 12311 13997
rect 12253 13957 12265 13991
rect 12299 13988 12311 13991
rect 12526 13988 12532 14000
rect 12299 13960 12532 13988
rect 12299 13957 12311 13960
rect 12253 13951 12311 13957
rect 12526 13948 12532 13960
rect 12584 13988 12590 14000
rect 14277 13991 14335 13997
rect 12584 13960 12940 13988
rect 12584 13948 12590 13960
rect 11241 13923 11299 13929
rect 9732 13892 9825 13920
rect 9732 13880 9738 13892
rect 11241 13889 11253 13923
rect 11287 13889 11299 13923
rect 11241 13883 11299 13889
rect 11425 13923 11483 13929
rect 11425 13889 11437 13923
rect 11471 13920 11483 13923
rect 12434 13920 12440 13932
rect 11471 13892 12440 13920
rect 11471 13889 11483 13892
rect 11425 13883 11483 13889
rect 12434 13880 12440 13892
rect 12492 13880 12498 13932
rect 12912 13929 12940 13960
rect 14277 13957 14289 13991
rect 14323 13988 14335 13991
rect 15010 13988 15016 14000
rect 14323 13960 15016 13988
rect 14323 13957 14335 13960
rect 14277 13951 14335 13957
rect 15010 13948 15016 13960
rect 15068 13948 15074 14000
rect 15286 13948 15292 14000
rect 15344 13988 15350 14000
rect 15657 13991 15715 13997
rect 15657 13988 15669 13991
rect 15344 13960 15669 13988
rect 15344 13948 15350 13960
rect 15657 13957 15669 13960
rect 15703 13988 15715 13991
rect 22005 13991 22063 13997
rect 15703 13960 18276 13988
rect 15703 13957 15715 13960
rect 15657 13951 15715 13957
rect 18248 13932 18276 13960
rect 22005 13957 22017 13991
rect 22051 13957 22063 13991
rect 22005 13951 22063 13957
rect 12897 13923 12955 13929
rect 12897 13889 12909 13923
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 14185 13923 14243 13929
rect 13044 13892 13089 13920
rect 13044 13880 13050 13892
rect 14185 13889 14197 13923
rect 14231 13920 14243 13923
rect 14918 13920 14924 13932
rect 14231 13892 14924 13920
rect 14231 13889 14243 13892
rect 14185 13883 14243 13889
rect 14918 13880 14924 13892
rect 14976 13880 14982 13932
rect 18230 13920 18236 13932
rect 18143 13892 18236 13920
rect 18230 13880 18236 13892
rect 18288 13880 18294 13932
rect 750 13812 756 13864
rect 808 13852 814 13864
rect 1581 13855 1639 13861
rect 1581 13852 1593 13855
rect 808 13824 1593 13852
rect 808 13812 814 13824
rect 1581 13821 1593 13824
rect 1627 13852 1639 13855
rect 2225 13855 2283 13861
rect 2225 13852 2237 13855
rect 1627 13824 2237 13852
rect 1627 13821 1639 13824
rect 1581 13815 1639 13821
rect 2225 13821 2237 13824
rect 2271 13852 2283 13855
rect 2682 13852 2688 13864
rect 2271 13824 2688 13852
rect 2271 13821 2283 13824
rect 2225 13815 2283 13821
rect 2682 13812 2688 13824
rect 2740 13812 2746 13864
rect 4062 13812 4068 13864
rect 4120 13852 4126 13864
rect 4709 13855 4767 13861
rect 4709 13852 4721 13855
rect 4120 13824 4721 13852
rect 4120 13812 4126 13824
rect 4709 13821 4721 13824
rect 4755 13852 4767 13855
rect 5166 13852 5172 13864
rect 4755 13824 5172 13852
rect 4755 13821 4767 13824
rect 4709 13815 4767 13821
rect 5166 13812 5172 13824
rect 5224 13852 5230 13864
rect 7006 13852 7012 13864
rect 5224 13824 7012 13852
rect 5224 13812 5230 13824
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 7101 13855 7159 13861
rect 7101 13821 7113 13855
rect 7147 13852 7159 13855
rect 7834 13852 7840 13864
rect 7147 13824 7840 13852
rect 7147 13821 7159 13824
rect 7101 13815 7159 13821
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 9033 13855 9091 13861
rect 9033 13821 9045 13855
rect 9079 13852 9091 13855
rect 9079 13824 9168 13852
rect 9079 13821 9091 13824
rect 9033 13815 9091 13821
rect 1670 13744 1676 13796
rect 1728 13784 1734 13796
rect 2314 13784 2320 13796
rect 1728 13756 2320 13784
rect 1728 13744 1734 13756
rect 2314 13744 2320 13756
rect 2372 13744 2378 13796
rect 4338 13744 4344 13796
rect 4396 13784 4402 13796
rect 4617 13787 4675 13793
rect 4617 13784 4629 13787
rect 4396 13756 4629 13784
rect 4396 13744 4402 13756
rect 4617 13753 4629 13756
rect 4663 13784 4675 13787
rect 8570 13784 8576 13796
rect 4663 13756 8576 13784
rect 4663 13753 4675 13756
rect 4617 13747 4675 13753
rect 8570 13744 8576 13756
rect 8628 13744 8634 13796
rect 9140 13784 9168 13824
rect 9214 13812 9220 13864
rect 9272 13852 9278 13864
rect 9493 13855 9551 13861
rect 9493 13852 9505 13855
rect 9272 13824 9505 13852
rect 9272 13812 9278 13824
rect 9493 13821 9505 13824
rect 9539 13821 9551 13855
rect 9692 13852 9720 13880
rect 9493 13815 9551 13821
rect 9600 13824 9720 13852
rect 9600 13784 9628 13824
rect 9766 13812 9772 13864
rect 9824 13852 9830 13864
rect 11146 13852 11152 13864
rect 9824 13824 10824 13852
rect 11107 13824 11152 13852
rect 9824 13812 9830 13824
rect 9140 13756 9628 13784
rect 1765 13719 1823 13725
rect 1765 13685 1777 13719
rect 1811 13716 1823 13719
rect 2038 13716 2044 13728
rect 1811 13688 2044 13716
rect 1811 13685 1823 13688
rect 1765 13679 1823 13685
rect 2038 13676 2044 13688
rect 2096 13676 2102 13728
rect 2133 13719 2191 13725
rect 2133 13685 2145 13719
rect 2179 13716 2191 13719
rect 2498 13716 2504 13728
rect 2179 13688 2504 13716
rect 2179 13685 2191 13688
rect 2133 13679 2191 13685
rect 2498 13676 2504 13688
rect 2556 13716 2562 13728
rect 2777 13719 2835 13725
rect 2777 13716 2789 13719
rect 2556 13688 2789 13716
rect 2556 13676 2562 13688
rect 2777 13685 2789 13688
rect 2823 13685 2835 13719
rect 4246 13716 4252 13728
rect 4207 13688 4252 13716
rect 2777 13679 2835 13685
rect 4246 13676 4252 13688
rect 4304 13676 4310 13728
rect 7006 13676 7012 13728
rect 7064 13716 7070 13728
rect 7929 13719 7987 13725
rect 7929 13716 7941 13719
rect 7064 13688 7941 13716
rect 7064 13676 7070 13688
rect 7929 13685 7941 13688
rect 7975 13716 7987 13719
rect 8110 13716 8116 13728
rect 7975 13688 8116 13716
rect 7975 13685 7987 13688
rect 7929 13679 7987 13685
rect 8110 13676 8116 13688
rect 8168 13676 8174 13728
rect 10796 13725 10824 13824
rect 11146 13812 11152 13824
rect 11204 13812 11210 13864
rect 14274 13852 14280 13864
rect 13740 13824 14280 13852
rect 11606 13744 11612 13796
rect 11664 13784 11670 13796
rect 11793 13787 11851 13793
rect 11793 13784 11805 13787
rect 11664 13756 11805 13784
rect 11664 13744 11670 13756
rect 11793 13753 11805 13756
rect 11839 13753 11851 13787
rect 12802 13784 12808 13796
rect 12763 13756 12808 13784
rect 11793 13747 11851 13753
rect 12802 13744 12808 13756
rect 12860 13744 12866 13796
rect 13630 13744 13636 13796
rect 13688 13784 13694 13796
rect 13740 13784 13768 13824
rect 14274 13812 14280 13824
rect 14332 13852 14338 13864
rect 14737 13855 14795 13861
rect 14737 13852 14749 13855
rect 14332 13824 14749 13852
rect 14332 13812 14338 13824
rect 14737 13821 14749 13824
rect 14783 13821 14795 13855
rect 14737 13815 14795 13821
rect 20257 13855 20315 13861
rect 20257 13821 20269 13855
rect 20303 13852 20315 13855
rect 20530 13852 20536 13864
rect 20303 13824 20536 13852
rect 20303 13821 20315 13824
rect 20257 13815 20315 13821
rect 20530 13812 20536 13824
rect 20588 13812 20594 13864
rect 22020 13852 22048 13951
rect 22480 13929 22508 14028
rect 23106 14016 23112 14028
rect 23164 14016 23170 14068
rect 25222 14016 25228 14068
rect 25280 14056 25286 14068
rect 27525 14059 27583 14065
rect 27525 14056 27537 14059
rect 25280 14028 27537 14056
rect 25280 14016 25286 14028
rect 27525 14025 27537 14028
rect 27571 14025 27583 14059
rect 27525 14019 27583 14025
rect 22465 13923 22523 13929
rect 22465 13889 22477 13923
rect 22511 13889 22523 13923
rect 22465 13883 22523 13889
rect 22649 13923 22707 13929
rect 22649 13889 22661 13923
rect 22695 13920 22707 13923
rect 23124 13920 23152 14016
rect 22695 13892 23152 13920
rect 22695 13889 22707 13892
rect 22649 13883 22707 13889
rect 23842 13880 23848 13932
rect 23900 13920 23906 13932
rect 24213 13923 24271 13929
rect 24213 13920 24225 13923
rect 23900 13892 24225 13920
rect 23900 13880 23906 13892
rect 24213 13889 24225 13892
rect 24259 13889 24271 13923
rect 24213 13883 24271 13889
rect 24026 13852 24032 13864
rect 22020 13824 24032 13852
rect 24026 13812 24032 13824
rect 24084 13852 24090 13864
rect 24121 13855 24179 13861
rect 24121 13852 24133 13855
rect 24084 13824 24133 13852
rect 24084 13812 24090 13824
rect 24121 13821 24133 13824
rect 24167 13821 24179 13855
rect 26142 13852 26148 13864
rect 26103 13824 26148 13852
rect 24121 13815 24179 13821
rect 26142 13812 26148 13824
rect 26200 13812 26206 13864
rect 13688 13756 13768 13784
rect 13817 13787 13875 13793
rect 13688 13744 13694 13756
rect 13817 13753 13829 13787
rect 13863 13784 13875 13787
rect 14642 13784 14648 13796
rect 13863 13756 14648 13784
rect 13863 13753 13875 13756
rect 13817 13747 13875 13753
rect 14642 13744 14648 13756
rect 14700 13744 14706 13796
rect 17497 13787 17555 13793
rect 17497 13753 17509 13787
rect 17543 13784 17555 13787
rect 17862 13784 17868 13796
rect 17543 13756 17868 13784
rect 17543 13753 17555 13756
rect 17497 13747 17555 13753
rect 17862 13744 17868 13756
rect 17920 13784 17926 13796
rect 18478 13787 18536 13793
rect 18478 13784 18490 13787
rect 17920 13756 18490 13784
rect 17920 13744 17926 13756
rect 18478 13753 18490 13756
rect 18524 13753 18536 13787
rect 26390 13787 26448 13793
rect 26390 13784 26402 13787
rect 18478 13747 18536 13753
rect 23492 13756 24072 13784
rect 23492 13728 23520 13756
rect 10781 13719 10839 13725
rect 10781 13685 10793 13719
rect 10827 13685 10839 13719
rect 10781 13679 10839 13685
rect 22094 13676 22100 13728
rect 22152 13716 22158 13728
rect 22373 13719 22431 13725
rect 22373 13716 22385 13719
rect 22152 13688 22385 13716
rect 22152 13676 22158 13688
rect 22373 13685 22385 13688
rect 22419 13685 22431 13719
rect 23474 13716 23480 13728
rect 23435 13688 23480 13716
rect 22373 13679 22431 13685
rect 23474 13676 23480 13688
rect 23532 13676 23538 13728
rect 23658 13716 23664 13728
rect 23619 13688 23664 13716
rect 23658 13676 23664 13688
rect 23716 13676 23722 13728
rect 24044 13725 24072 13756
rect 26068 13756 26402 13784
rect 26068 13728 26096 13756
rect 26390 13753 26402 13756
rect 26436 13753 26448 13787
rect 26390 13747 26448 13753
rect 24029 13719 24087 13725
rect 24029 13685 24041 13719
rect 24075 13685 24087 13719
rect 26050 13716 26056 13728
rect 26011 13688 26056 13716
rect 24029 13679 24087 13685
rect 26050 13676 26056 13688
rect 26108 13676 26114 13728
rect 1104 13626 28888 13648
rect 1104 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 20982 13626
rect 21034 13574 21046 13626
rect 21098 13574 21110 13626
rect 21162 13574 21174 13626
rect 21226 13574 28888 13626
rect 1104 13552 28888 13574
rect 1670 13512 1676 13524
rect 1631 13484 1676 13512
rect 1670 13472 1676 13484
rect 1728 13472 1734 13524
rect 1854 13472 1860 13524
rect 1912 13472 1918 13524
rect 2038 13472 2044 13524
rect 2096 13512 2102 13524
rect 2225 13515 2283 13521
rect 2225 13512 2237 13515
rect 2096 13484 2237 13512
rect 2096 13472 2102 13484
rect 2225 13481 2237 13484
rect 2271 13512 2283 13515
rect 2777 13515 2835 13521
rect 2777 13512 2789 13515
rect 2271 13484 2789 13512
rect 2271 13481 2283 13484
rect 2225 13475 2283 13481
rect 2777 13481 2789 13484
rect 2823 13481 2835 13515
rect 6822 13512 6828 13524
rect 6783 13484 6828 13512
rect 2777 13475 2835 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 7006 13472 7012 13524
rect 7064 13512 7070 13524
rect 7561 13515 7619 13521
rect 7561 13512 7573 13515
rect 7064 13484 7573 13512
rect 7064 13472 7070 13484
rect 7561 13481 7573 13484
rect 7607 13481 7619 13515
rect 7561 13475 7619 13481
rect 8021 13515 8079 13521
rect 8021 13481 8033 13515
rect 8067 13512 8079 13515
rect 8202 13512 8208 13524
rect 8067 13484 8208 13512
rect 8067 13481 8079 13484
rect 8021 13475 8079 13481
rect 8202 13472 8208 13484
rect 8260 13472 8266 13524
rect 9030 13472 9036 13524
rect 9088 13512 9094 13524
rect 9125 13515 9183 13521
rect 9125 13512 9137 13515
rect 9088 13484 9137 13512
rect 9088 13472 9094 13484
rect 9125 13481 9137 13484
rect 9171 13481 9183 13515
rect 9125 13475 9183 13481
rect 9214 13472 9220 13524
rect 9272 13512 9278 13524
rect 9677 13515 9735 13521
rect 9677 13512 9689 13515
rect 9272 13484 9689 13512
rect 9272 13472 9278 13484
rect 9677 13481 9689 13484
rect 9723 13481 9735 13515
rect 10870 13512 10876 13524
rect 10831 13484 10876 13512
rect 9677 13475 9735 13481
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 11330 13512 11336 13524
rect 11291 13484 11336 13512
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 11698 13512 11704 13524
rect 11659 13484 11704 13512
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 12158 13512 12164 13524
rect 12119 13484 12164 13512
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 13630 13512 13636 13524
rect 13591 13484 13636 13512
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 14642 13472 14648 13524
rect 14700 13512 14706 13524
rect 15289 13515 15347 13521
rect 15289 13512 15301 13515
rect 14700 13484 15301 13512
rect 14700 13472 14706 13484
rect 15289 13481 15301 13484
rect 15335 13481 15347 13515
rect 15289 13475 15347 13481
rect 15657 13515 15715 13521
rect 15657 13481 15669 13515
rect 15703 13512 15715 13515
rect 16298 13512 16304 13524
rect 15703 13484 16304 13512
rect 15703 13481 15715 13484
rect 15657 13475 15715 13481
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 18785 13515 18843 13521
rect 18785 13481 18797 13515
rect 18831 13512 18843 13515
rect 18874 13512 18880 13524
rect 18831 13484 18880 13512
rect 18831 13481 18843 13484
rect 18785 13475 18843 13481
rect 18874 13472 18880 13484
rect 18932 13472 18938 13524
rect 22554 13512 22560 13524
rect 22515 13484 22560 13512
rect 22554 13472 22560 13484
rect 22612 13472 22618 13524
rect 24026 13512 24032 13524
rect 23987 13484 24032 13512
rect 24026 13472 24032 13484
rect 24084 13472 24090 13524
rect 24857 13515 24915 13521
rect 24857 13481 24869 13515
rect 24903 13512 24915 13515
rect 25038 13512 25044 13524
rect 24903 13484 25044 13512
rect 24903 13481 24915 13484
rect 24857 13475 24915 13481
rect 25038 13472 25044 13484
rect 25096 13472 25102 13524
rect 26234 13512 26240 13524
rect 26147 13484 26240 13512
rect 26234 13472 26240 13484
rect 26292 13512 26298 13524
rect 26418 13512 26424 13524
rect 26292 13484 26424 13512
rect 26292 13472 26298 13484
rect 26418 13472 26424 13484
rect 26476 13472 26482 13524
rect 1872 13444 1900 13472
rect 4706 13444 4712 13456
rect 1688 13416 1900 13444
rect 4667 13416 4712 13444
rect 1688 13388 1716 13416
rect 4706 13404 4712 13416
rect 4764 13404 4770 13456
rect 12066 13444 12072 13456
rect 12027 13416 12072 13444
rect 12066 13404 12072 13416
rect 12124 13404 12130 13456
rect 14093 13447 14151 13453
rect 14093 13444 14105 13447
rect 13648 13416 14105 13444
rect 13648 13388 13676 13416
rect 14093 13413 14105 13416
rect 14139 13413 14151 13447
rect 14093 13407 14151 13413
rect 15378 13404 15384 13456
rect 15436 13444 15442 13456
rect 15838 13444 15844 13456
rect 15436 13416 15844 13444
rect 15436 13404 15442 13416
rect 15838 13404 15844 13416
rect 15896 13444 15902 13456
rect 15896 13416 15976 13444
rect 15896 13404 15902 13416
rect 1670 13336 1676 13388
rect 1728 13336 1734 13388
rect 1854 13336 1860 13388
rect 1912 13376 1918 13388
rect 2133 13379 2191 13385
rect 2133 13376 2145 13379
rect 1912 13348 2145 13376
rect 1912 13336 1918 13348
rect 2133 13345 2145 13348
rect 2179 13345 2191 13379
rect 2133 13339 2191 13345
rect 4617 13379 4675 13385
rect 4617 13345 4629 13379
rect 4663 13376 4675 13379
rect 5074 13376 5080 13388
rect 4663 13348 5080 13376
rect 4663 13345 4675 13348
rect 4617 13339 4675 13345
rect 5074 13336 5080 13348
rect 5132 13336 5138 13388
rect 8386 13376 8392 13388
rect 8347 13348 8392 13376
rect 8386 13336 8392 13348
rect 8444 13336 8450 13388
rect 10045 13379 10103 13385
rect 10045 13345 10057 13379
rect 10091 13376 10103 13379
rect 10091 13348 10824 13376
rect 10091 13345 10103 13348
rect 10045 13339 10103 13345
rect 2409 13311 2467 13317
rect 2409 13277 2421 13311
rect 2455 13308 2467 13311
rect 2590 13308 2596 13320
rect 2455 13280 2596 13308
rect 2455 13277 2467 13280
rect 2409 13271 2467 13277
rect 2590 13268 2596 13280
rect 2648 13308 2654 13320
rect 2866 13308 2872 13320
rect 2648 13280 2872 13308
rect 2648 13268 2654 13280
rect 2866 13268 2872 13280
rect 2924 13268 2930 13320
rect 4798 13308 4804 13320
rect 4759 13280 4804 13308
rect 4798 13268 4804 13280
rect 4856 13268 4862 13320
rect 10134 13308 10140 13320
rect 10095 13280 10140 13308
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 7926 13200 7932 13252
rect 7984 13240 7990 13252
rect 8205 13243 8263 13249
rect 8205 13240 8217 13243
rect 7984 13212 8217 13240
rect 7984 13200 7990 13212
rect 8205 13209 8217 13212
rect 8251 13209 8263 13243
rect 8205 13203 8263 13209
rect 9674 13200 9680 13252
rect 9732 13240 9738 13252
rect 10244 13240 10272 13271
rect 10796 13252 10824 13348
rect 13630 13336 13636 13388
rect 13688 13336 13694 13388
rect 13998 13376 14004 13388
rect 13959 13348 14004 13376
rect 13998 13336 14004 13348
rect 14056 13336 14062 13388
rect 15396 13376 15424 13404
rect 14292 13348 15424 13376
rect 11606 13268 11612 13320
rect 11664 13308 11670 13320
rect 12253 13311 12311 13317
rect 12253 13308 12265 13311
rect 11664 13280 12265 13308
rect 11664 13268 11670 13280
rect 12253 13277 12265 13280
rect 12299 13308 12311 13311
rect 12986 13308 12992 13320
rect 12299 13280 12992 13308
rect 12299 13277 12311 13280
rect 12253 13271 12311 13277
rect 12986 13268 12992 13280
rect 13044 13268 13050 13320
rect 13722 13268 13728 13320
rect 13780 13308 13786 13320
rect 14292 13317 14320 13348
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 13780 13280 14289 13308
rect 13780 13268 13786 13280
rect 14277 13277 14289 13280
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 15194 13268 15200 13320
rect 15252 13308 15258 13320
rect 15948 13317 15976 13416
rect 17954 13404 17960 13456
rect 18012 13444 18018 13456
rect 18230 13444 18236 13456
rect 18012 13416 18236 13444
rect 18012 13404 18018 13416
rect 18230 13404 18236 13416
rect 18288 13444 18294 13456
rect 19061 13447 19119 13453
rect 19061 13444 19073 13447
rect 18288 13416 19073 13444
rect 18288 13404 18294 13416
rect 19061 13413 19073 13416
rect 19107 13413 19119 13447
rect 19061 13407 19119 13413
rect 23658 13404 23664 13456
rect 23716 13444 23722 13456
rect 25317 13447 25375 13453
rect 25317 13444 25329 13447
rect 23716 13416 25329 13444
rect 23716 13404 23722 13416
rect 25317 13413 25329 13416
rect 25363 13413 25375 13447
rect 25317 13407 25375 13413
rect 25222 13376 25228 13388
rect 25183 13348 25228 13376
rect 25222 13336 25228 13348
rect 25280 13336 25286 13388
rect 15749 13311 15807 13317
rect 15749 13308 15761 13311
rect 15252 13280 15761 13308
rect 15252 13268 15258 13280
rect 15749 13277 15761 13280
rect 15795 13277 15807 13311
rect 15749 13271 15807 13277
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13277 15991 13311
rect 15933 13271 15991 13277
rect 25314 13268 25320 13320
rect 25372 13308 25378 13320
rect 25501 13311 25559 13317
rect 25501 13308 25513 13311
rect 25372 13280 25513 13308
rect 25372 13268 25378 13280
rect 25501 13277 25513 13280
rect 25547 13308 25559 13311
rect 26050 13308 26056 13320
rect 25547 13280 26056 13308
rect 25547 13277 25559 13280
rect 25501 13271 25559 13277
rect 26050 13268 26056 13280
rect 26108 13308 26114 13320
rect 26510 13308 26516 13320
rect 26108 13280 26516 13308
rect 26108 13268 26114 13280
rect 26510 13268 26516 13280
rect 26568 13268 26574 13320
rect 10410 13240 10416 13252
rect 9732 13212 10416 13240
rect 9732 13200 9738 13212
rect 10410 13200 10416 13212
rect 10468 13200 10474 13252
rect 10778 13200 10784 13252
rect 10836 13240 10842 13252
rect 19150 13240 19156 13252
rect 10836 13212 19156 13240
rect 10836 13200 10842 13212
rect 19150 13200 19156 13212
rect 19208 13200 19214 13252
rect 1765 13175 1823 13181
rect 1765 13141 1777 13175
rect 1811 13172 1823 13175
rect 2406 13172 2412 13184
rect 1811 13144 2412 13172
rect 1811 13141 1823 13144
rect 1765 13135 1823 13141
rect 2406 13132 2412 13144
rect 2464 13172 2470 13184
rect 3145 13175 3203 13181
rect 3145 13172 3157 13175
rect 2464 13144 3157 13172
rect 2464 13132 2470 13144
rect 3145 13141 3157 13144
rect 3191 13141 3203 13175
rect 3145 13135 3203 13141
rect 3697 13175 3755 13181
rect 3697 13141 3709 13175
rect 3743 13172 3755 13175
rect 4062 13172 4068 13184
rect 3743 13144 4068 13172
rect 3743 13141 3755 13144
rect 3697 13135 3755 13141
rect 4062 13132 4068 13144
rect 4120 13172 4126 13184
rect 4249 13175 4307 13181
rect 4249 13172 4261 13175
rect 4120 13144 4261 13172
rect 4120 13132 4126 13144
rect 4249 13141 4261 13144
rect 4295 13141 4307 13175
rect 4249 13135 4307 13141
rect 4338 13132 4344 13184
rect 4396 13172 4402 13184
rect 4522 13172 4528 13184
rect 4396 13144 4528 13172
rect 4396 13132 4402 13144
rect 4522 13132 4528 13144
rect 4580 13132 4586 13184
rect 18417 13175 18475 13181
rect 18417 13141 18429 13175
rect 18463 13172 18475 13175
rect 18506 13172 18512 13184
rect 18463 13144 18512 13172
rect 18463 13141 18475 13144
rect 18417 13135 18475 13141
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 22094 13132 22100 13184
rect 22152 13172 22158 13184
rect 23753 13175 23811 13181
rect 22152 13144 22197 13172
rect 22152 13132 22158 13144
rect 23753 13141 23765 13175
rect 23799 13172 23811 13175
rect 23842 13172 23848 13184
rect 23799 13144 23848 13172
rect 23799 13141 23811 13144
rect 23753 13135 23811 13141
rect 23842 13132 23848 13144
rect 23900 13132 23906 13184
rect 24670 13132 24676 13184
rect 24728 13172 24734 13184
rect 25498 13172 25504 13184
rect 24728 13144 25504 13172
rect 24728 13132 24734 13144
rect 25498 13132 25504 13144
rect 25556 13132 25562 13184
rect 1104 13082 28888 13104
rect 1104 13030 5982 13082
rect 6034 13030 6046 13082
rect 6098 13030 6110 13082
rect 6162 13030 6174 13082
rect 6226 13030 15982 13082
rect 16034 13030 16046 13082
rect 16098 13030 16110 13082
rect 16162 13030 16174 13082
rect 16226 13030 25982 13082
rect 26034 13030 26046 13082
rect 26098 13030 26110 13082
rect 26162 13030 26174 13082
rect 26226 13030 28888 13082
rect 1104 13008 28888 13030
rect 3510 12968 3516 12980
rect 3471 12940 3516 12968
rect 3510 12928 3516 12940
rect 3568 12928 3574 12980
rect 4706 12968 4712 12980
rect 4667 12940 4712 12968
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 8386 12928 8392 12980
rect 8444 12968 8450 12980
rect 8757 12971 8815 12977
rect 8757 12968 8769 12971
rect 8444 12940 8769 12968
rect 8444 12928 8450 12940
rect 8757 12937 8769 12940
rect 8803 12968 8815 12971
rect 8846 12968 8852 12980
rect 8803 12940 8852 12968
rect 8803 12937 8815 12940
rect 8757 12931 8815 12937
rect 8846 12928 8852 12940
rect 8904 12928 8910 12980
rect 10410 12968 10416 12980
rect 10371 12940 10416 12968
rect 10410 12928 10416 12940
rect 10468 12968 10474 12980
rect 11333 12971 11391 12977
rect 11333 12968 11345 12971
rect 10468 12940 11345 12968
rect 10468 12928 10474 12940
rect 11333 12937 11345 12940
rect 11379 12968 11391 12971
rect 11606 12968 11612 12980
rect 11379 12940 11612 12968
rect 11379 12937 11391 12940
rect 11333 12931 11391 12937
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 12158 12968 12164 12980
rect 12119 12940 12164 12968
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 13630 12968 13636 12980
rect 13591 12940 13636 12968
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 15838 12928 15844 12980
rect 15896 12968 15902 12980
rect 16025 12971 16083 12977
rect 16025 12968 16037 12971
rect 15896 12940 16037 12968
rect 15896 12928 15902 12940
rect 16025 12937 16037 12940
rect 16071 12937 16083 12971
rect 17862 12968 17868 12980
rect 17823 12940 17868 12968
rect 16025 12931 16083 12937
rect 17862 12928 17868 12940
rect 17920 12928 17926 12980
rect 23658 12928 23664 12980
rect 23716 12968 23722 12980
rect 24213 12971 24271 12977
rect 24213 12968 24225 12971
rect 23716 12940 24225 12968
rect 23716 12928 23722 12940
rect 24213 12937 24225 12940
rect 24259 12937 24271 12971
rect 24213 12931 24271 12937
rect 25222 12928 25228 12980
rect 25280 12968 25286 12980
rect 25501 12971 25559 12977
rect 25501 12968 25513 12971
rect 25280 12940 25513 12968
rect 25280 12928 25286 12940
rect 25501 12937 25513 12940
rect 25547 12968 25559 12971
rect 26513 12971 26571 12977
rect 26513 12968 26525 12971
rect 25547 12940 26525 12968
rect 25547 12937 25559 12940
rect 25501 12931 25559 12937
rect 26513 12937 26525 12940
rect 26559 12937 26571 12971
rect 26513 12931 26571 12937
rect 5074 12900 5080 12912
rect 5035 12872 5080 12900
rect 5074 12860 5080 12872
rect 5132 12860 5138 12912
rect 11793 12903 11851 12909
rect 11793 12869 11805 12903
rect 11839 12900 11851 12903
rect 12066 12900 12072 12912
rect 11839 12872 12072 12900
rect 11839 12869 11851 12872
rect 11793 12863 11851 12869
rect 12066 12860 12072 12872
rect 12124 12860 12130 12912
rect 14274 12900 14280 12912
rect 14235 12872 14280 12900
rect 14274 12860 14280 12872
rect 14332 12860 14338 12912
rect 15749 12903 15807 12909
rect 15749 12900 15761 12903
rect 14384 12872 15761 12900
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12832 2743 12835
rect 3053 12835 3111 12841
rect 3053 12832 3065 12835
rect 2731 12804 3065 12832
rect 2731 12801 2743 12804
rect 2685 12795 2743 12801
rect 3053 12801 3065 12804
rect 3099 12832 3111 12835
rect 3142 12832 3148 12844
rect 3099 12804 3148 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 3510 12792 3516 12844
rect 3568 12832 3574 12844
rect 4157 12835 4215 12841
rect 4157 12832 4169 12835
rect 3568 12804 4169 12832
rect 3568 12792 3574 12804
rect 4157 12801 4169 12804
rect 4203 12801 4215 12835
rect 6822 12832 6828 12844
rect 6783 12804 6828 12832
rect 4157 12795 4215 12801
rect 6822 12792 6828 12804
rect 6880 12792 6886 12844
rect 10134 12832 10140 12844
rect 10047 12804 10140 12832
rect 10134 12792 10140 12804
rect 10192 12832 10198 12844
rect 14384 12832 14412 12872
rect 15749 12869 15761 12872
rect 15795 12900 15807 12903
rect 16298 12900 16304 12912
rect 15795 12872 16304 12900
rect 15795 12869 15807 12872
rect 15749 12863 15807 12869
rect 16298 12860 16304 12872
rect 16356 12860 16362 12912
rect 14918 12832 14924 12844
rect 10192 12804 14412 12832
rect 14879 12804 14924 12832
rect 10192 12792 10198 12804
rect 14918 12792 14924 12804
rect 14976 12792 14982 12844
rect 17880 12832 17908 12928
rect 24673 12903 24731 12909
rect 24673 12869 24685 12903
rect 24719 12900 24731 12903
rect 25314 12900 25320 12912
rect 24719 12872 25320 12900
rect 24719 12869 24731 12872
rect 24673 12863 24731 12869
rect 25314 12860 25320 12872
rect 25372 12860 25378 12912
rect 18598 12832 18604 12844
rect 17880 12804 18604 12832
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 20438 12832 20444 12844
rect 20399 12804 20444 12832
rect 20438 12792 20444 12804
rect 20496 12792 20502 12844
rect 26050 12832 26056 12844
rect 26011 12804 26056 12832
rect 26050 12792 26056 12804
rect 26108 12792 26114 12844
rect 2406 12764 2412 12776
rect 2367 12736 2412 12764
rect 2406 12724 2412 12736
rect 2464 12724 2470 12776
rect 4062 12764 4068 12776
rect 4023 12736 4068 12764
rect 4062 12724 4068 12736
rect 4120 12724 4126 12776
rect 10042 12724 10048 12776
rect 10100 12764 10106 12776
rect 13265 12767 13323 12773
rect 13265 12764 13277 12767
rect 10100 12736 13277 12764
rect 10100 12724 10106 12736
rect 13265 12733 13277 12736
rect 13311 12764 13323 12767
rect 13998 12764 14004 12776
rect 13311 12736 14004 12764
rect 13311 12733 13323 12736
rect 13265 12727 13323 12733
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 25038 12764 25044 12776
rect 24951 12736 25044 12764
rect 25038 12724 25044 12736
rect 25096 12764 25102 12776
rect 25774 12764 25780 12776
rect 25096 12736 25780 12764
rect 25096 12724 25102 12736
rect 25774 12724 25780 12736
rect 25832 12764 25838 12776
rect 25961 12767 26019 12773
rect 25961 12764 25973 12767
rect 25832 12736 25973 12764
rect 25832 12724 25838 12736
rect 25961 12733 25973 12736
rect 26007 12733 26019 12767
rect 25961 12727 26019 12733
rect 2501 12699 2559 12705
rect 2501 12665 2513 12699
rect 2547 12696 2559 12699
rect 3973 12699 4031 12705
rect 2547 12668 3648 12696
rect 2547 12665 2559 12668
rect 2501 12659 2559 12665
rect 3620 12640 3648 12668
rect 3973 12665 3985 12699
rect 4019 12696 4031 12699
rect 4246 12696 4252 12708
rect 4019 12668 4252 12696
rect 4019 12665 4031 12668
rect 3973 12659 4031 12665
rect 4246 12656 4252 12668
rect 4304 12696 4310 12708
rect 5353 12699 5411 12705
rect 5353 12696 5365 12699
rect 4304 12668 5365 12696
rect 4304 12656 4310 12668
rect 5353 12665 5365 12668
rect 5399 12665 5411 12699
rect 5353 12659 5411 12665
rect 6641 12699 6699 12705
rect 6641 12665 6653 12699
rect 6687 12696 6699 12699
rect 6730 12696 6736 12708
rect 6687 12668 6736 12696
rect 6687 12665 6699 12668
rect 6641 12659 6699 12665
rect 6730 12656 6736 12668
rect 6788 12696 6794 12708
rect 7070 12699 7128 12705
rect 7070 12696 7082 12699
rect 6788 12668 7082 12696
rect 6788 12656 6794 12668
rect 7070 12665 7082 12668
rect 7116 12665 7128 12699
rect 7070 12659 7128 12665
rect 16758 12656 16764 12708
rect 16816 12696 16822 12708
rect 17497 12699 17555 12705
rect 17497 12696 17509 12699
rect 16816 12668 17509 12696
rect 16816 12656 16822 12668
rect 17497 12665 17509 12668
rect 17543 12696 17555 12699
rect 18509 12699 18567 12705
rect 18509 12696 18521 12699
rect 17543 12668 18521 12696
rect 17543 12665 17555 12668
rect 17497 12659 17555 12665
rect 18509 12665 18521 12668
rect 18555 12665 18567 12699
rect 18509 12659 18567 12665
rect 20349 12699 20407 12705
rect 20349 12665 20361 12699
rect 20395 12696 20407 12699
rect 20708 12699 20766 12705
rect 20708 12696 20720 12699
rect 20395 12668 20720 12696
rect 20395 12665 20407 12668
rect 20349 12659 20407 12665
rect 20708 12665 20720 12668
rect 20754 12696 20766 12699
rect 20806 12696 20812 12708
rect 20754 12668 20812 12696
rect 20754 12665 20766 12668
rect 20708 12659 20766 12665
rect 20806 12656 20812 12668
rect 20864 12656 20870 12708
rect 21726 12656 21732 12708
rect 21784 12696 21790 12708
rect 25314 12696 25320 12708
rect 21784 12668 25320 12696
rect 21784 12656 21790 12668
rect 25314 12656 25320 12668
rect 25372 12696 25378 12708
rect 25869 12699 25927 12705
rect 25869 12696 25881 12699
rect 25372 12668 25881 12696
rect 25372 12656 25378 12668
rect 25869 12665 25881 12668
rect 25915 12665 25927 12699
rect 25869 12659 25927 12665
rect 1854 12628 1860 12640
rect 1815 12600 1860 12628
rect 1854 12588 1860 12600
rect 1912 12588 1918 12640
rect 2038 12628 2044 12640
rect 1999 12600 2044 12628
rect 2038 12588 2044 12600
rect 2096 12588 2102 12640
rect 3602 12628 3608 12640
rect 3563 12600 3608 12628
rect 3602 12588 3608 12600
rect 3660 12588 3666 12640
rect 8202 12628 8208 12640
rect 8163 12600 8208 12628
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 14185 12631 14243 12637
rect 9732 12600 9777 12628
rect 9732 12588 9738 12600
rect 14185 12597 14197 12631
rect 14231 12628 14243 12631
rect 14642 12628 14648 12640
rect 14231 12600 14648 12628
rect 14231 12597 14243 12600
rect 14185 12591 14243 12597
rect 14642 12588 14648 12600
rect 14700 12588 14706 12640
rect 14734 12588 14740 12640
rect 14792 12628 14798 12640
rect 14792 12600 14837 12628
rect 14792 12588 14798 12600
rect 15194 12588 15200 12640
rect 15252 12628 15258 12640
rect 15381 12631 15439 12637
rect 15381 12628 15393 12631
rect 15252 12600 15393 12628
rect 15252 12588 15258 12600
rect 15381 12597 15393 12600
rect 15427 12628 15439 12631
rect 15470 12628 15476 12640
rect 15427 12600 15476 12628
rect 15427 12597 15439 12600
rect 15381 12591 15439 12597
rect 15470 12588 15476 12600
rect 15528 12588 15534 12640
rect 18046 12628 18052 12640
rect 18007 12600 18052 12628
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 18417 12631 18475 12637
rect 18417 12597 18429 12631
rect 18463 12628 18475 12631
rect 19150 12628 19156 12640
rect 18463 12600 19156 12628
rect 18463 12597 18475 12600
rect 18417 12591 18475 12597
rect 19150 12588 19156 12600
rect 19208 12588 19214 12640
rect 21542 12588 21548 12640
rect 21600 12628 21606 12640
rect 21821 12631 21879 12637
rect 21821 12628 21833 12631
rect 21600 12600 21833 12628
rect 21600 12588 21606 12600
rect 21821 12597 21833 12600
rect 21867 12597 21879 12631
rect 21821 12591 21879 12597
rect 24854 12588 24860 12640
rect 24912 12628 24918 12640
rect 25038 12628 25044 12640
rect 24912 12600 25044 12628
rect 24912 12588 24918 12600
rect 25038 12588 25044 12600
rect 25096 12588 25102 12640
rect 1104 12538 28888 12560
rect 1104 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 20982 12538
rect 21034 12486 21046 12538
rect 21098 12486 21110 12538
rect 21162 12486 21174 12538
rect 21226 12486 28888 12538
rect 1104 12464 28888 12486
rect 3053 12427 3111 12433
rect 3053 12393 3065 12427
rect 3099 12424 3111 12427
rect 3602 12424 3608 12436
rect 3099 12396 3608 12424
rect 3099 12393 3111 12396
rect 3053 12387 3111 12393
rect 3602 12384 3608 12396
rect 3660 12384 3666 12436
rect 4062 12384 4068 12436
rect 4120 12424 4126 12436
rect 4338 12424 4344 12436
rect 4120 12396 4344 12424
rect 4120 12384 4126 12396
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 13722 12424 13728 12436
rect 13683 12396 13728 12424
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 18598 12384 18604 12436
rect 18656 12424 18662 12436
rect 19153 12427 19211 12433
rect 19153 12424 19165 12427
rect 18656 12396 19165 12424
rect 18656 12384 18662 12396
rect 19153 12393 19165 12396
rect 19199 12393 19211 12427
rect 20438 12424 20444 12436
rect 20399 12396 20444 12424
rect 19153 12387 19211 12393
rect 20438 12384 20444 12396
rect 20496 12384 20502 12436
rect 20714 12384 20720 12436
rect 20772 12424 20778 12436
rect 20901 12427 20959 12433
rect 20901 12424 20913 12427
rect 20772 12396 20913 12424
rect 20772 12384 20778 12396
rect 20901 12393 20913 12396
rect 20947 12393 20959 12427
rect 24762 12424 24768 12436
rect 20901 12387 20959 12393
rect 24596 12396 24768 12424
rect 24596 12368 24624 12396
rect 24762 12384 24768 12396
rect 24820 12384 24826 12436
rect 24946 12384 24952 12436
rect 25004 12424 25010 12436
rect 25004 12396 25452 12424
rect 25004 12384 25010 12396
rect 25424 12368 25452 12396
rect 26510 12384 26516 12436
rect 26568 12424 26574 12436
rect 26694 12424 26700 12436
rect 26568 12396 26700 12424
rect 26568 12384 26574 12396
rect 26694 12384 26700 12396
rect 26752 12384 26758 12436
rect 26970 12424 26976 12436
rect 26931 12396 26976 12424
rect 26970 12384 26976 12396
rect 27028 12384 27034 12436
rect 2682 12316 2688 12368
rect 2740 12356 2746 12368
rect 2866 12356 2872 12368
rect 2740 12328 2872 12356
rect 2740 12316 2746 12328
rect 2866 12316 2872 12328
rect 2924 12316 2930 12368
rect 17954 12316 17960 12368
rect 18012 12365 18018 12368
rect 18012 12359 18076 12365
rect 18012 12325 18030 12359
rect 18064 12325 18076 12359
rect 18012 12319 18076 12325
rect 18012 12316 18018 12319
rect 24302 12316 24308 12368
rect 24360 12356 24366 12368
rect 24486 12356 24492 12368
rect 24360 12328 24492 12356
rect 24360 12316 24366 12328
rect 24486 12316 24492 12328
rect 24544 12316 24550 12368
rect 24578 12316 24584 12368
rect 24636 12316 24642 12368
rect 25406 12316 25412 12368
rect 25464 12316 25470 12368
rect 26418 12316 26424 12368
rect 26476 12356 26482 12368
rect 26988 12356 27016 12384
rect 26476 12328 27016 12356
rect 26476 12316 26482 12328
rect 2314 12288 2320 12300
rect 2275 12260 2320 12288
rect 2314 12248 2320 12260
rect 2372 12248 2378 12300
rect 2409 12291 2467 12297
rect 2409 12257 2421 12291
rect 2455 12288 2467 12291
rect 2958 12288 2964 12300
rect 2455 12260 2964 12288
rect 2455 12257 2467 12260
rect 2409 12251 2467 12257
rect 2958 12248 2964 12260
rect 3016 12248 3022 12300
rect 4505 12291 4563 12297
rect 4505 12288 4517 12291
rect 3620 12260 4517 12288
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12220 1915 12223
rect 2590 12220 2596 12232
rect 1903 12192 2596 12220
rect 1903 12189 1915 12192
rect 1857 12183 1915 12189
rect 2590 12180 2596 12192
rect 2648 12220 2654 12232
rect 3510 12220 3516 12232
rect 2648 12192 3516 12220
rect 2648 12180 2654 12192
rect 3510 12180 3516 12192
rect 3568 12220 3574 12232
rect 3620 12229 3648 12260
rect 4505 12257 4517 12260
rect 4551 12257 4563 12291
rect 10594 12288 10600 12300
rect 10555 12260 10600 12288
rect 4505 12251 4563 12257
rect 10594 12248 10600 12260
rect 10652 12248 10658 12300
rect 15654 12288 15660 12300
rect 15615 12260 15660 12288
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 17773 12291 17831 12297
rect 17773 12257 17785 12291
rect 17819 12288 17831 12291
rect 17862 12288 17868 12300
rect 17819 12260 17868 12288
rect 17819 12257 17831 12260
rect 17773 12251 17831 12257
rect 17862 12248 17868 12260
rect 17920 12248 17926 12300
rect 21269 12291 21327 12297
rect 21269 12257 21281 12291
rect 21315 12288 21327 12291
rect 21634 12288 21640 12300
rect 21315 12260 21640 12288
rect 21315 12257 21327 12260
rect 21269 12251 21327 12257
rect 21634 12248 21640 12260
rect 21692 12248 21698 12300
rect 25222 12288 25228 12300
rect 25183 12260 25228 12288
rect 25222 12248 25228 12260
rect 25280 12248 25286 12300
rect 25317 12291 25375 12297
rect 25317 12257 25329 12291
rect 25363 12288 25375 12291
rect 25590 12288 25596 12300
rect 25363 12260 25596 12288
rect 25363 12257 25375 12260
rect 25317 12251 25375 12257
rect 25590 12248 25596 12260
rect 25648 12248 25654 12300
rect 26510 12248 26516 12300
rect 26568 12288 26574 12300
rect 26881 12291 26939 12297
rect 26881 12288 26893 12291
rect 26568 12260 26893 12288
rect 26568 12248 26574 12260
rect 26881 12257 26893 12260
rect 26927 12257 26939 12291
rect 26881 12251 26939 12257
rect 3605 12223 3663 12229
rect 3605 12220 3617 12223
rect 3568 12192 3617 12220
rect 3568 12180 3574 12192
rect 3605 12189 3617 12192
rect 3651 12189 3663 12223
rect 4246 12220 4252 12232
rect 4207 12192 4252 12220
rect 3605 12183 3663 12189
rect 4246 12180 4252 12192
rect 4304 12180 4310 12232
rect 10410 12180 10416 12232
rect 10468 12220 10474 12232
rect 10689 12223 10747 12229
rect 10689 12220 10701 12223
rect 10468 12192 10701 12220
rect 10468 12180 10474 12192
rect 10689 12189 10701 12192
rect 10735 12189 10747 12223
rect 10689 12183 10747 12189
rect 10778 12180 10784 12232
rect 10836 12220 10842 12232
rect 15749 12223 15807 12229
rect 10836 12192 10881 12220
rect 10836 12180 10842 12192
rect 15749 12189 15761 12223
rect 15795 12220 15807 12223
rect 15838 12220 15844 12232
rect 15795 12192 15844 12220
rect 15795 12189 15807 12192
rect 15749 12183 15807 12189
rect 15838 12180 15844 12192
rect 15896 12180 15902 12232
rect 15930 12180 15936 12232
rect 15988 12220 15994 12232
rect 16666 12220 16672 12232
rect 15988 12192 16672 12220
rect 15988 12180 15994 12192
rect 16666 12180 16672 12192
rect 16724 12180 16730 12232
rect 21358 12220 21364 12232
rect 21319 12192 21364 12220
rect 21358 12180 21364 12192
rect 21416 12180 21422 12232
rect 21542 12220 21548 12232
rect 21503 12192 21548 12220
rect 21542 12180 21548 12192
rect 21600 12180 21606 12232
rect 22462 12220 22468 12232
rect 22423 12192 22468 12220
rect 22462 12180 22468 12192
rect 22520 12180 22526 12232
rect 23934 12180 23940 12232
rect 23992 12220 23998 12232
rect 24486 12220 24492 12232
rect 23992 12192 24492 12220
rect 23992 12180 23998 12192
rect 24486 12180 24492 12192
rect 24544 12180 24550 12232
rect 25501 12223 25559 12229
rect 25501 12189 25513 12223
rect 25547 12189 25559 12223
rect 27062 12220 27068 12232
rect 27023 12192 27068 12220
rect 25501 12183 25559 12189
rect 5626 12152 5632 12164
rect 5587 12124 5632 12152
rect 5626 12112 5632 12124
rect 5684 12112 5690 12164
rect 14734 12152 14740 12164
rect 14647 12124 14740 12152
rect 14734 12112 14740 12124
rect 14792 12152 14798 12164
rect 15289 12155 15347 12161
rect 15289 12152 15301 12155
rect 14792 12124 15301 12152
rect 14792 12112 14798 12124
rect 15289 12121 15301 12124
rect 15335 12121 15347 12155
rect 15289 12115 15347 12121
rect 23842 12112 23848 12164
rect 23900 12152 23906 12164
rect 24762 12152 24768 12164
rect 23900 12124 24768 12152
rect 23900 12112 23906 12124
rect 24762 12112 24768 12124
rect 24820 12152 24826 12164
rect 25516 12152 25544 12183
rect 27062 12180 27068 12192
rect 27120 12180 27126 12232
rect 25961 12155 26019 12161
rect 25961 12152 25973 12155
rect 24820 12124 25973 12152
rect 24820 12112 24826 12124
rect 25961 12121 25973 12124
rect 26007 12152 26019 12155
rect 26050 12152 26056 12164
rect 26007 12124 26056 12152
rect 26007 12121 26019 12124
rect 25961 12115 26019 12121
rect 26050 12112 26056 12124
rect 26108 12152 26114 12164
rect 27080 12152 27108 12180
rect 26108 12124 27108 12152
rect 26108 12112 26114 12124
rect 1946 12084 1952 12096
rect 1907 12056 1952 12084
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 6914 12084 6920 12096
rect 6875 12056 6920 12084
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 10229 12087 10287 12093
rect 10229 12053 10241 12087
rect 10275 12084 10287 12087
rect 10318 12084 10324 12096
rect 10275 12056 10324 12084
rect 10275 12053 10287 12056
rect 10229 12047 10287 12053
rect 10318 12044 10324 12056
rect 10376 12044 10382 12096
rect 12710 12044 12716 12096
rect 12768 12084 12774 12096
rect 14277 12087 14335 12093
rect 14277 12084 14289 12087
rect 12768 12056 14289 12084
rect 12768 12044 12774 12056
rect 14277 12053 14289 12056
rect 14323 12084 14335 12087
rect 14918 12084 14924 12096
rect 14323 12056 14924 12084
rect 14323 12053 14335 12056
rect 14277 12047 14335 12053
rect 14918 12044 14924 12056
rect 14976 12084 14982 12096
rect 15378 12084 15384 12096
rect 14976 12056 15384 12084
rect 14976 12044 14982 12056
rect 15378 12044 15384 12056
rect 15436 12044 15442 12096
rect 16298 12084 16304 12096
rect 16259 12056 16304 12084
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 24210 12084 24216 12096
rect 24171 12056 24216 12084
rect 24210 12044 24216 12056
rect 24268 12044 24274 12096
rect 24854 12084 24860 12096
rect 24815 12056 24860 12084
rect 24854 12044 24860 12056
rect 24912 12044 24918 12096
rect 26513 12087 26571 12093
rect 26513 12053 26525 12087
rect 26559 12084 26571 12087
rect 27154 12084 27160 12096
rect 26559 12056 27160 12084
rect 26559 12053 26571 12056
rect 26513 12047 26571 12053
rect 27154 12044 27160 12056
rect 27212 12044 27218 12096
rect 27522 12084 27528 12096
rect 27483 12056 27528 12084
rect 27522 12044 27528 12056
rect 27580 12044 27586 12096
rect 1104 11994 28888 12016
rect 1104 11942 5982 11994
rect 6034 11942 6046 11994
rect 6098 11942 6110 11994
rect 6162 11942 6174 11994
rect 6226 11942 15982 11994
rect 16034 11942 16046 11994
rect 16098 11942 16110 11994
rect 16162 11942 16174 11994
rect 16226 11942 25982 11994
rect 26034 11942 26046 11994
rect 26098 11942 26110 11994
rect 26162 11942 26174 11994
rect 26226 11942 28888 11994
rect 1104 11920 28888 11942
rect 1673 11883 1731 11889
rect 1673 11849 1685 11883
rect 1719 11880 1731 11883
rect 2314 11880 2320 11892
rect 1719 11852 2320 11880
rect 1719 11849 1731 11852
rect 1673 11843 1731 11849
rect 2314 11840 2320 11852
rect 2372 11840 2378 11892
rect 2590 11840 2596 11892
rect 2648 11880 2654 11892
rect 3145 11883 3203 11889
rect 3145 11880 3157 11883
rect 2648 11852 3157 11880
rect 2648 11840 2654 11852
rect 3145 11849 3157 11852
rect 3191 11849 3203 11883
rect 3970 11880 3976 11892
rect 3931 11852 3976 11880
rect 3145 11843 3203 11849
rect 3160 11812 3188 11843
rect 3970 11840 3976 11852
rect 4028 11840 4034 11892
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 4893 11883 4951 11889
rect 4893 11880 4905 11883
rect 4304 11852 4905 11880
rect 4304 11840 4310 11852
rect 4893 11849 4905 11852
rect 4939 11849 4951 11883
rect 4893 11843 4951 11849
rect 5442 11840 5448 11892
rect 5500 11880 5506 11892
rect 6549 11883 6607 11889
rect 6549 11880 6561 11883
rect 5500 11852 6561 11880
rect 5500 11840 5506 11852
rect 6549 11849 6561 11852
rect 6595 11849 6607 11883
rect 6549 11843 6607 11849
rect 4341 11815 4399 11821
rect 4341 11812 4353 11815
rect 3160 11784 4353 11812
rect 4341 11781 4353 11784
rect 4387 11781 4399 11815
rect 6564 11812 6592 11843
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 10781 11883 10839 11889
rect 10781 11880 10793 11883
rect 10652 11852 10793 11880
rect 10652 11840 10658 11852
rect 10781 11849 10793 11852
rect 10827 11849 10839 11883
rect 15102 11880 15108 11892
rect 15063 11852 15108 11880
rect 10781 11843 10839 11849
rect 8202 11812 8208 11824
rect 6564 11784 8208 11812
rect 4341 11775 4399 11781
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 3142 11744 3148 11756
rect 2455 11716 3148 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 3142 11704 3148 11716
rect 3200 11704 3206 11756
rect 4430 11744 4436 11756
rect 4391 11716 4436 11744
rect 4430 11704 4436 11716
rect 4488 11704 4494 11756
rect 6914 11704 6920 11756
rect 6972 11744 6978 11756
rect 7392 11753 7420 11784
rect 8202 11772 8208 11784
rect 8260 11772 8266 11824
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 6972 11716 7297 11744
rect 6972 11704 6978 11716
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11713 7435 11747
rect 8478 11744 8484 11756
rect 8439 11716 8484 11744
rect 7377 11707 7435 11713
rect 8478 11704 8484 11716
rect 8536 11704 8542 11756
rect 10796 11744 10824 11843
rect 15102 11840 15108 11852
rect 15160 11840 15166 11892
rect 16666 11880 16672 11892
rect 16627 11852 16672 11880
rect 16666 11840 16672 11852
rect 16724 11840 16730 11892
rect 21358 11840 21364 11892
rect 21416 11880 21422 11892
rect 21453 11883 21511 11889
rect 21453 11880 21465 11883
rect 21416 11852 21465 11880
rect 21416 11840 21422 11852
rect 21453 11849 21465 11852
rect 21499 11849 21511 11883
rect 21453 11843 21511 11849
rect 24121 11883 24179 11889
rect 24121 11849 24133 11883
rect 24167 11880 24179 11883
rect 25222 11880 25228 11892
rect 24167 11852 25228 11880
rect 24167 11849 24179 11852
rect 24121 11843 24179 11849
rect 25222 11840 25228 11852
rect 25280 11840 25286 11892
rect 26326 11840 26332 11892
rect 26384 11880 26390 11892
rect 26697 11883 26755 11889
rect 26697 11880 26709 11883
rect 26384 11852 26709 11880
rect 26384 11840 26390 11852
rect 26697 11849 26709 11852
rect 26743 11849 26755 11883
rect 26697 11843 26755 11849
rect 14918 11772 14924 11824
rect 14976 11812 14982 11824
rect 14976 11784 16344 11812
rect 14976 11772 14982 11784
rect 16316 11756 16344 11784
rect 17402 11772 17408 11824
rect 17460 11812 17466 11824
rect 17497 11815 17555 11821
rect 17497 11812 17509 11815
rect 17460 11784 17509 11812
rect 17460 11772 17466 11784
rect 17497 11781 17509 11784
rect 17543 11812 17555 11815
rect 17954 11812 17960 11824
rect 17543 11784 17960 11812
rect 17543 11781 17555 11784
rect 17497 11775 17555 11781
rect 17954 11772 17960 11784
rect 18012 11812 18018 11824
rect 20625 11815 20683 11821
rect 20625 11812 20637 11815
rect 18012 11784 20637 11812
rect 18012 11772 18018 11784
rect 20625 11781 20637 11784
rect 20671 11812 20683 11815
rect 21542 11812 21548 11824
rect 20671 11784 21548 11812
rect 20671 11781 20683 11784
rect 20625 11775 20683 11781
rect 21542 11772 21548 11784
rect 21600 11772 21606 11824
rect 25593 11815 25651 11821
rect 25593 11781 25605 11815
rect 25639 11781 25651 11815
rect 25593 11775 25651 11781
rect 26237 11815 26295 11821
rect 26237 11781 26249 11815
rect 26283 11812 26295 11815
rect 26418 11812 26424 11824
rect 26283 11784 26424 11812
rect 26283 11781 26295 11784
rect 26237 11775 26295 11781
rect 10965 11747 11023 11753
rect 10965 11744 10977 11747
rect 10796 11716 10977 11744
rect 10965 11713 10977 11716
rect 11011 11713 11023 11747
rect 13630 11744 13636 11756
rect 13591 11716 13636 11744
rect 10965 11707 11023 11713
rect 13630 11704 13636 11716
rect 13688 11744 13694 11756
rect 13688 11716 13860 11744
rect 13688 11704 13694 11716
rect 3329 11679 3387 11685
rect 3329 11645 3341 11679
rect 3375 11676 3387 11679
rect 3970 11676 3976 11688
rect 3375 11648 3976 11676
rect 3375 11645 3387 11648
rect 3329 11639 3387 11645
rect 3970 11636 3976 11648
rect 4028 11636 4034 11688
rect 13832 11685 13860 11716
rect 15010 11704 15016 11756
rect 15068 11744 15074 11756
rect 16114 11744 16120 11756
rect 15068 11716 16120 11744
rect 15068 11704 15074 11716
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 16298 11744 16304 11756
rect 16259 11716 16304 11744
rect 16298 11704 16304 11716
rect 16356 11704 16362 11756
rect 17865 11747 17923 11753
rect 17865 11713 17877 11747
rect 17911 11744 17923 11747
rect 19061 11747 19119 11753
rect 19061 11744 19073 11747
rect 17911 11716 19073 11744
rect 17911 11713 17923 11716
rect 17865 11707 17923 11713
rect 19061 11713 19073 11716
rect 19107 11744 19119 11747
rect 19150 11744 19156 11756
rect 19107 11716 19156 11744
rect 19107 11713 19119 11716
rect 19061 11707 19119 11713
rect 19150 11704 19156 11716
rect 19208 11744 19214 11756
rect 20806 11744 20812 11756
rect 19208 11716 20812 11744
rect 19208 11704 19214 11716
rect 20806 11704 20812 11716
rect 20864 11744 20870 11756
rect 20993 11747 21051 11753
rect 20993 11744 21005 11747
rect 20864 11716 21005 11744
rect 20864 11704 20870 11716
rect 20993 11713 21005 11716
rect 21039 11744 21051 11747
rect 22097 11747 22155 11753
rect 22097 11744 22109 11747
rect 21039 11716 22109 11744
rect 21039 11713 21051 11716
rect 20993 11707 21051 11713
rect 22097 11713 22109 11716
rect 22143 11744 22155 11747
rect 22278 11744 22284 11756
rect 22143 11716 22284 11744
rect 22143 11713 22155 11716
rect 22097 11707 22155 11713
rect 22278 11704 22284 11716
rect 22336 11704 22342 11756
rect 25608 11744 25636 11775
rect 26418 11772 26424 11784
rect 26476 11772 26482 11824
rect 26528 11784 27384 11812
rect 26528 11744 26556 11784
rect 26694 11744 26700 11756
rect 25608 11716 26700 11744
rect 26694 11704 26700 11716
rect 26752 11704 26758 11756
rect 27154 11744 27160 11756
rect 27115 11716 27160 11744
rect 27154 11704 27160 11716
rect 27212 11704 27218 11756
rect 27356 11753 27384 11784
rect 27341 11747 27399 11753
rect 27341 11713 27353 11747
rect 27387 11744 27399 11747
rect 27709 11747 27767 11753
rect 27709 11744 27721 11747
rect 27387 11716 27721 11744
rect 27387 11713 27399 11716
rect 27341 11707 27399 11713
rect 27709 11713 27721 11716
rect 27755 11713 27767 11747
rect 27709 11707 27767 11713
rect 13817 11679 13875 11685
rect 13817 11645 13829 11679
rect 13863 11645 13875 11679
rect 13817 11639 13875 11645
rect 14274 11636 14280 11688
rect 14332 11676 14338 11688
rect 16025 11679 16083 11685
rect 16025 11676 16037 11679
rect 14332 11648 16037 11676
rect 14332 11636 14338 11648
rect 16025 11645 16037 11648
rect 16071 11676 16083 11679
rect 17037 11679 17095 11685
rect 17037 11676 17049 11679
rect 16071 11648 17049 11676
rect 16071 11645 16083 11648
rect 16025 11639 16083 11645
rect 17037 11645 17049 11648
rect 17083 11645 17095 11679
rect 21266 11676 21272 11688
rect 21227 11648 21272 11676
rect 17037 11639 17095 11645
rect 21266 11636 21272 11648
rect 21324 11676 21330 11688
rect 21821 11679 21879 11685
rect 21821 11676 21833 11679
rect 21324 11648 21833 11676
rect 21324 11636 21330 11648
rect 21821 11645 21833 11648
rect 21867 11676 21879 11679
rect 23842 11676 23848 11688
rect 21867 11648 23848 11676
rect 21867 11645 21879 11648
rect 21821 11639 21879 11645
rect 23842 11636 23848 11648
rect 23900 11636 23906 11688
rect 24210 11676 24216 11688
rect 24171 11648 24216 11676
rect 24210 11636 24216 11648
rect 24268 11636 24274 11688
rect 24480 11679 24538 11685
rect 24480 11645 24492 11679
rect 24526 11676 24538 11679
rect 24762 11676 24768 11688
rect 24526 11648 24768 11676
rect 24526 11645 24538 11648
rect 24480 11639 24538 11645
rect 24762 11636 24768 11648
rect 24820 11636 24826 11688
rect 24854 11636 24860 11688
rect 24912 11676 24918 11688
rect 27065 11679 27123 11685
rect 27065 11676 27077 11679
rect 24912 11648 27077 11676
rect 24912 11636 24918 11648
rect 27065 11645 27077 11648
rect 27111 11676 27123 11679
rect 27522 11676 27528 11688
rect 27111 11648 27528 11676
rect 27111 11645 27123 11648
rect 27065 11639 27123 11645
rect 27522 11636 27528 11648
rect 27580 11636 27586 11688
rect 6273 11611 6331 11617
rect 6273 11577 6285 11611
rect 6319 11608 6331 11611
rect 8726 11611 8784 11617
rect 8726 11608 8738 11611
rect 6319 11580 7236 11608
rect 6319 11577 6331 11580
rect 6273 11571 6331 11577
rect 7208 11552 7236 11580
rect 8312 11580 8738 11608
rect 8312 11552 8340 11580
rect 8726 11577 8738 11580
rect 8772 11577 8784 11611
rect 8726 11571 8784 11577
rect 18138 11568 18144 11620
rect 18196 11608 18202 11620
rect 18325 11611 18383 11617
rect 18325 11608 18337 11611
rect 18196 11580 18337 11608
rect 18196 11568 18202 11580
rect 18325 11577 18337 11580
rect 18371 11608 18383 11611
rect 18785 11611 18843 11617
rect 18785 11608 18797 11611
rect 18371 11580 18797 11608
rect 18371 11577 18383 11580
rect 18325 11571 18383 11577
rect 18785 11577 18797 11580
rect 18831 11608 18843 11611
rect 19058 11608 19064 11620
rect 18831 11580 19064 11608
rect 18831 11577 18843 11580
rect 18785 11571 18843 11577
rect 19058 11568 19064 11580
rect 19116 11568 19122 11620
rect 20257 11611 20315 11617
rect 20257 11577 20269 11611
rect 20303 11608 20315 11611
rect 21634 11608 21640 11620
rect 20303 11580 21640 11608
rect 20303 11577 20315 11580
rect 20257 11571 20315 11577
rect 21634 11568 21640 11580
rect 21692 11568 21698 11620
rect 25774 11568 25780 11620
rect 25832 11608 25838 11620
rect 27246 11608 27252 11620
rect 25832 11580 27252 11608
rect 25832 11568 25838 11580
rect 27246 11568 27252 11580
rect 27304 11568 27310 11620
rect 1762 11540 1768 11552
rect 1723 11512 1768 11540
rect 1762 11500 1768 11512
rect 1820 11500 1826 11552
rect 1946 11500 1952 11552
rect 2004 11540 2010 11552
rect 2130 11540 2136 11552
rect 2004 11512 2136 11540
rect 2004 11500 2010 11512
rect 2130 11500 2136 11512
rect 2188 11500 2194 11552
rect 2222 11500 2228 11552
rect 2280 11540 2286 11552
rect 2869 11543 2927 11549
rect 2280 11512 2325 11540
rect 2280 11500 2286 11512
rect 2869 11509 2881 11543
rect 2915 11540 2927 11543
rect 2958 11540 2964 11552
rect 2915 11512 2964 11540
rect 2915 11509 2927 11512
rect 2869 11503 2927 11509
rect 2958 11500 2964 11512
rect 3016 11500 3022 11552
rect 3510 11540 3516 11552
rect 3471 11512 3516 11540
rect 3510 11500 3516 11512
rect 3568 11500 3574 11552
rect 6822 11540 6828 11552
rect 6783 11512 6828 11540
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 7190 11540 7196 11552
rect 7151 11512 7196 11540
rect 7190 11500 7196 11512
rect 7248 11500 7254 11552
rect 8294 11540 8300 11552
rect 8255 11512 8300 11540
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 9582 11500 9588 11552
rect 9640 11540 9646 11552
rect 9861 11543 9919 11549
rect 9861 11540 9873 11543
rect 9640 11512 9873 11540
rect 9640 11500 9646 11512
rect 9861 11509 9873 11512
rect 9907 11509 9919 11543
rect 10410 11540 10416 11552
rect 10371 11512 10416 11540
rect 9861 11503 9919 11509
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 15194 11500 15200 11552
rect 15252 11540 15258 11552
rect 15657 11543 15715 11549
rect 15657 11540 15669 11543
rect 15252 11512 15669 11540
rect 15252 11500 15258 11512
rect 15657 11509 15669 11512
rect 15703 11509 15715 11543
rect 18414 11540 18420 11552
rect 18375 11512 18420 11540
rect 15657 11503 15715 11509
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 18874 11500 18880 11552
rect 18932 11540 18938 11552
rect 19429 11543 19487 11549
rect 19429 11540 19441 11543
rect 18932 11512 19441 11540
rect 18932 11500 18938 11512
rect 19429 11509 19441 11512
rect 19475 11509 19487 11543
rect 19429 11503 19487 11509
rect 21450 11500 21456 11552
rect 21508 11540 21514 11552
rect 21913 11543 21971 11549
rect 21913 11540 21925 11543
rect 21508 11512 21925 11540
rect 21508 11500 21514 11512
rect 21913 11509 21925 11512
rect 21959 11540 21971 11543
rect 22002 11540 22008 11552
rect 21959 11512 22008 11540
rect 21959 11509 21971 11512
rect 21913 11503 21971 11509
rect 22002 11500 22008 11512
rect 22060 11500 22066 11552
rect 26510 11540 26516 11552
rect 26471 11512 26516 11540
rect 26510 11500 26516 11512
rect 26568 11500 26574 11552
rect 1104 11450 28888 11472
rect 1104 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 20982 11450
rect 21034 11398 21046 11450
rect 21098 11398 21110 11450
rect 21162 11398 21174 11450
rect 21226 11398 28888 11450
rect 1104 11376 28888 11398
rect 1949 11339 2007 11345
rect 1949 11305 1961 11339
rect 1995 11336 2007 11339
rect 2222 11336 2228 11348
rect 1995 11308 2228 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 2222 11296 2228 11308
rect 2280 11336 2286 11348
rect 3329 11339 3387 11345
rect 3329 11336 3341 11339
rect 2280 11308 3341 11336
rect 2280 11296 2286 11308
rect 3329 11305 3341 11308
rect 3375 11305 3387 11339
rect 3329 11299 3387 11305
rect 6549 11339 6607 11345
rect 6549 11305 6561 11339
rect 6595 11336 6607 11339
rect 6914 11336 6920 11348
rect 6595 11308 6920 11336
rect 6595 11305 6607 11308
rect 6549 11299 6607 11305
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 8478 11336 8484 11348
rect 8439 11308 8484 11336
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 9674 11336 9680 11348
rect 9635 11308 9680 11336
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 16114 11296 16120 11348
rect 16172 11336 16178 11348
rect 16485 11339 16543 11345
rect 16485 11336 16497 11339
rect 16172 11308 16497 11336
rect 16172 11296 16178 11308
rect 16485 11305 16497 11308
rect 16531 11305 16543 11339
rect 16758 11336 16764 11348
rect 16719 11308 16764 11336
rect 16485 11299 16543 11305
rect 16758 11296 16764 11308
rect 16816 11296 16822 11348
rect 17862 11336 17868 11348
rect 17823 11308 17868 11336
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 21177 11339 21235 11345
rect 21177 11305 21189 11339
rect 21223 11336 21235 11339
rect 21358 11336 21364 11348
rect 21223 11308 21364 11336
rect 21223 11305 21235 11308
rect 21177 11299 21235 11305
rect 21358 11296 21364 11308
rect 21416 11296 21422 11348
rect 21634 11336 21640 11348
rect 21595 11308 21640 11336
rect 21634 11296 21640 11308
rect 21692 11296 21698 11348
rect 22005 11339 22063 11345
rect 22005 11305 22017 11339
rect 22051 11336 22063 11339
rect 22094 11336 22100 11348
rect 22051 11308 22100 11336
rect 22051 11305 22063 11308
rect 22005 11299 22063 11305
rect 22094 11296 22100 11308
rect 22152 11336 22158 11348
rect 22462 11336 22468 11348
rect 22152 11308 22468 11336
rect 22152 11296 22158 11308
rect 22462 11296 22468 11308
rect 22520 11296 22526 11348
rect 24305 11339 24363 11345
rect 24305 11305 24317 11339
rect 24351 11336 24363 11339
rect 24762 11336 24768 11348
rect 24351 11308 24768 11336
rect 24351 11305 24363 11308
rect 24305 11299 24363 11305
rect 24762 11296 24768 11308
rect 24820 11296 24826 11348
rect 25682 11336 25688 11348
rect 24872 11308 25688 11336
rect 1394 11228 1400 11280
rect 1452 11268 1458 11280
rect 1673 11271 1731 11277
rect 1673 11268 1685 11271
rect 1452 11240 1685 11268
rect 1452 11228 1458 11240
rect 1673 11237 1685 11240
rect 1719 11268 1731 11271
rect 2958 11268 2964 11280
rect 1719 11240 2964 11268
rect 1719 11237 1731 11240
rect 1673 11231 1731 11237
rect 2958 11228 2964 11240
rect 3016 11228 3022 11280
rect 3053 11271 3111 11277
rect 3053 11237 3065 11271
rect 3099 11268 3111 11271
rect 3142 11268 3148 11280
rect 3099 11240 3148 11268
rect 3099 11237 3111 11240
rect 3053 11231 3111 11237
rect 3142 11228 3148 11240
rect 3200 11228 3206 11280
rect 17129 11271 17187 11277
rect 17129 11237 17141 11271
rect 17175 11268 17187 11271
rect 17218 11268 17224 11280
rect 17175 11240 17224 11268
rect 17175 11237 17187 11240
rect 17129 11231 17187 11237
rect 17218 11228 17224 11240
rect 17276 11268 17282 11280
rect 18414 11268 18420 11280
rect 17276 11240 18420 11268
rect 17276 11228 17282 11240
rect 18414 11228 18420 11240
rect 18472 11228 18478 11280
rect 2222 11160 2228 11212
rect 2280 11200 2286 11212
rect 2317 11203 2375 11209
rect 2317 11200 2329 11203
rect 2280 11172 2329 11200
rect 2280 11160 2286 11172
rect 2317 11169 2329 11172
rect 2363 11200 2375 11203
rect 2682 11200 2688 11212
rect 2363 11172 2688 11200
rect 2363 11169 2375 11172
rect 2317 11163 2375 11169
rect 2682 11160 2688 11172
rect 2740 11160 2746 11212
rect 6914 11200 6920 11212
rect 6875 11172 6920 11200
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 10045 11203 10103 11209
rect 10045 11169 10057 11203
rect 10091 11200 10103 11203
rect 10318 11200 10324 11212
rect 10091 11172 10324 11200
rect 10091 11169 10103 11172
rect 10045 11163 10103 11169
rect 10318 11160 10324 11172
rect 10376 11200 10382 11212
rect 10962 11200 10968 11212
rect 10376 11172 10968 11200
rect 10376 11160 10382 11172
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 12710 11209 12716 11212
rect 12704 11163 12716 11209
rect 12768 11200 12774 11212
rect 12768 11172 12804 11200
rect 12710 11160 12716 11163
rect 12768 11160 12774 11172
rect 15654 11160 15660 11212
rect 15712 11200 15718 11212
rect 16117 11203 16175 11209
rect 16117 11200 16129 11203
rect 15712 11172 16129 11200
rect 15712 11160 15718 11172
rect 16117 11169 16129 11172
rect 16163 11169 16175 11203
rect 16117 11163 16175 11169
rect 17954 11160 17960 11212
rect 18012 11200 18018 11212
rect 18690 11200 18696 11212
rect 18012 11172 18696 11200
rect 18012 11160 18018 11172
rect 18690 11160 18696 11172
rect 18748 11160 18754 11212
rect 21726 11160 21732 11212
rect 21784 11200 21790 11212
rect 22097 11203 22155 11209
rect 22097 11200 22109 11203
rect 21784 11172 22109 11200
rect 21784 11160 21790 11172
rect 22097 11169 22109 11172
rect 22143 11200 22155 11203
rect 24872 11200 24900 11308
rect 25682 11296 25688 11308
rect 25740 11296 25746 11348
rect 26694 11336 26700 11348
rect 26655 11308 26700 11336
rect 26694 11296 26700 11308
rect 26752 11296 26758 11348
rect 27062 11336 27068 11348
rect 27023 11308 27068 11336
rect 27062 11296 27068 11308
rect 27120 11296 27126 11348
rect 27154 11296 27160 11348
rect 27212 11336 27218 11348
rect 27433 11339 27491 11345
rect 27433 11336 27445 11339
rect 27212 11308 27445 11336
rect 27212 11296 27218 11308
rect 27433 11305 27445 11308
rect 27479 11305 27491 11339
rect 27614 11336 27620 11348
rect 27575 11308 27620 11336
rect 27433 11299 27491 11305
rect 27614 11296 27620 11308
rect 27672 11296 27678 11348
rect 24949 11271 25007 11277
rect 24949 11237 24961 11271
rect 24995 11268 25007 11271
rect 25498 11268 25504 11280
rect 24995 11240 25504 11268
rect 24995 11237 25007 11240
rect 24949 11231 25007 11237
rect 25498 11228 25504 11240
rect 25556 11228 25562 11280
rect 25590 11228 25596 11280
rect 25648 11268 25654 11280
rect 27338 11268 27344 11280
rect 25648 11240 27344 11268
rect 25648 11228 25654 11240
rect 27338 11228 27344 11240
rect 27396 11228 27402 11280
rect 25314 11200 25320 11212
rect 22143 11172 24900 11200
rect 25275 11172 25320 11200
rect 22143 11169 22155 11172
rect 22097 11163 22155 11169
rect 25314 11160 25320 11172
rect 25372 11160 25378 11212
rect 26510 11200 26516 11212
rect 26471 11172 26516 11200
rect 26510 11160 26516 11172
rect 26568 11160 26574 11212
rect 2409 11135 2467 11141
rect 2409 11101 2421 11135
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 2424 11064 2452 11095
rect 2498 11092 2504 11144
rect 2556 11132 2562 11144
rect 7006 11132 7012 11144
rect 2556 11104 2601 11132
rect 6967 11104 7012 11132
rect 2556 11092 2562 11104
rect 7006 11092 7012 11104
rect 7064 11092 7070 11144
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11101 7159 11135
rect 10134 11132 10140 11144
rect 10095 11104 10140 11132
rect 7101 11095 7159 11101
rect 2774 11064 2780 11076
rect 2424 11036 2780 11064
rect 2774 11024 2780 11036
rect 2832 11024 2838 11076
rect 6730 11024 6736 11076
rect 6788 11064 6794 11076
rect 7116 11064 7144 11095
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 10229 11135 10287 11141
rect 10229 11101 10241 11135
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 6788 11036 7144 11064
rect 6788 11024 6794 11036
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 10244 11064 10272 11095
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 15286 11132 15292 11144
rect 12492 11104 12537 11132
rect 15247 11104 15292 11132
rect 12492 11092 12498 11104
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 17221 11135 17279 11141
rect 17221 11101 17233 11135
rect 17267 11101 17279 11135
rect 17402 11132 17408 11144
rect 17363 11104 17408 11132
rect 17221 11095 17279 11101
rect 15838 11064 15844 11076
rect 9732 11036 10272 11064
rect 15799 11036 15844 11064
rect 9732 11024 9738 11036
rect 15838 11024 15844 11036
rect 15896 11024 15902 11076
rect 16850 11024 16856 11076
rect 16908 11064 16914 11076
rect 17236 11064 17264 11095
rect 17402 11092 17408 11104
rect 17460 11092 17466 11144
rect 18782 11132 18788 11144
rect 18743 11104 18788 11132
rect 18782 11092 18788 11104
rect 18840 11092 18846 11144
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11132 18935 11135
rect 19150 11132 19156 11144
rect 18923 11104 19156 11132
rect 18923 11101 18935 11104
rect 18877 11095 18935 11101
rect 18325 11067 18383 11073
rect 18325 11064 18337 11067
rect 16908 11036 18337 11064
rect 16908 11024 16914 11036
rect 18325 11033 18337 11036
rect 18371 11033 18383 11067
rect 18325 11027 18383 11033
rect 18414 11024 18420 11076
rect 18472 11064 18478 11076
rect 18892 11064 18920 11095
rect 19150 11092 19156 11104
rect 19208 11092 19214 11144
rect 22278 11132 22284 11144
rect 22191 11104 22284 11132
rect 22278 11092 22284 11104
rect 22336 11132 22342 11144
rect 22462 11132 22468 11144
rect 22336 11104 22468 11132
rect 22336 11092 22342 11104
rect 22462 11092 22468 11104
rect 22520 11092 22526 11144
rect 19426 11064 19432 11076
rect 18472 11036 18920 11064
rect 19387 11036 19432 11064
rect 18472 11024 18478 11036
rect 19426 11024 19432 11036
rect 19484 11024 19490 11076
rect 21450 11064 21456 11076
rect 21411 11036 21456 11064
rect 21450 11024 21456 11036
rect 21508 11024 21514 11076
rect 25498 11064 25504 11076
rect 25459 11036 25504 11064
rect 25498 11024 25504 11036
rect 25556 11024 25562 11076
rect 7653 10999 7711 11005
rect 7653 10965 7665 10999
rect 7699 10996 7711 10999
rect 7834 10996 7840 11008
rect 7699 10968 7840 10996
rect 7699 10965 7711 10968
rect 7653 10959 7711 10965
rect 7834 10956 7840 10968
rect 7892 10956 7898 11008
rect 10686 10996 10692 11008
rect 10647 10968 10692 10996
rect 10686 10956 10692 10968
rect 10744 10956 10750 11008
rect 13538 10956 13544 11008
rect 13596 10996 13602 11008
rect 13817 10999 13875 11005
rect 13817 10996 13829 10999
rect 13596 10968 13829 10996
rect 13596 10956 13602 10968
rect 13817 10965 13829 10968
rect 13863 10996 13875 10999
rect 14182 10996 14188 11008
rect 13863 10968 14188 10996
rect 13863 10965 13875 10968
rect 13817 10959 13875 10965
rect 14182 10956 14188 10968
rect 14240 10956 14246 11008
rect 14458 10996 14464 11008
rect 14419 10968 14464 10996
rect 14458 10956 14464 10968
rect 14516 10956 14522 11008
rect 1104 10906 28888 10928
rect 1104 10854 5982 10906
rect 6034 10854 6046 10906
rect 6098 10854 6110 10906
rect 6162 10854 6174 10906
rect 6226 10854 15982 10906
rect 16034 10854 16046 10906
rect 16098 10854 16110 10906
rect 16162 10854 16174 10906
rect 16226 10854 25982 10906
rect 26034 10854 26046 10906
rect 26098 10854 26110 10906
rect 26162 10854 26174 10906
rect 26226 10854 28888 10906
rect 1104 10832 28888 10854
rect 2041 10795 2099 10801
rect 2041 10761 2053 10795
rect 2087 10792 2099 10795
rect 2222 10792 2228 10804
rect 2087 10764 2228 10792
rect 2087 10761 2099 10764
rect 2041 10755 2099 10761
rect 2222 10752 2228 10764
rect 2280 10752 2286 10804
rect 2314 10752 2320 10804
rect 2372 10792 2378 10804
rect 2409 10795 2467 10801
rect 2409 10792 2421 10795
rect 2372 10764 2421 10792
rect 2372 10752 2378 10764
rect 2409 10761 2421 10764
rect 2455 10792 2467 10795
rect 2774 10792 2780 10804
rect 2455 10764 2780 10792
rect 2455 10761 2467 10764
rect 2409 10755 2467 10761
rect 2774 10752 2780 10764
rect 2832 10752 2838 10804
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7101 10795 7159 10801
rect 7101 10792 7113 10795
rect 6972 10764 7113 10792
rect 6972 10752 6978 10764
rect 7101 10761 7113 10764
rect 7147 10761 7159 10795
rect 7101 10755 7159 10761
rect 8849 10795 8907 10801
rect 8849 10761 8861 10795
rect 8895 10792 8907 10795
rect 10045 10795 10103 10801
rect 10045 10792 10057 10795
rect 8895 10764 10057 10792
rect 8895 10761 8907 10764
rect 8849 10755 8907 10761
rect 10045 10761 10057 10764
rect 10091 10792 10103 10795
rect 10134 10792 10140 10804
rect 10091 10764 10140 10792
rect 10091 10761 10103 10764
rect 10045 10755 10103 10761
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 11054 10792 11060 10804
rect 11015 10764 11060 10792
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 12710 10792 12716 10804
rect 12671 10764 12716 10792
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 14182 10792 14188 10804
rect 14095 10764 14188 10792
rect 14182 10752 14188 10764
rect 14240 10792 14246 10804
rect 14918 10792 14924 10804
rect 14240 10764 14924 10792
rect 14240 10752 14246 10764
rect 14918 10752 14924 10764
rect 14976 10752 14982 10804
rect 15286 10792 15292 10804
rect 15247 10764 15292 10792
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 16945 10795 17003 10801
rect 16945 10761 16957 10795
rect 16991 10792 17003 10795
rect 17402 10792 17408 10804
rect 16991 10764 17408 10792
rect 16991 10761 17003 10764
rect 16945 10755 17003 10761
rect 17402 10752 17408 10764
rect 17460 10752 17466 10804
rect 17497 10795 17555 10801
rect 17497 10761 17509 10795
rect 17543 10792 17555 10795
rect 17862 10792 17868 10804
rect 17543 10764 17868 10792
rect 17543 10761 17555 10764
rect 17497 10755 17555 10761
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 18874 10792 18880 10804
rect 18835 10764 18880 10792
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 21726 10792 21732 10804
rect 21687 10764 21732 10792
rect 21726 10752 21732 10764
rect 21784 10752 21790 10804
rect 22094 10752 22100 10804
rect 22152 10792 22158 10804
rect 25314 10792 25320 10804
rect 22152 10764 22197 10792
rect 25275 10764 25320 10792
rect 22152 10752 22158 10764
rect 25314 10752 25320 10764
rect 25372 10752 25378 10804
rect 26510 10752 26516 10804
rect 26568 10792 26574 10804
rect 27341 10795 27399 10801
rect 27341 10792 27353 10795
rect 26568 10764 27353 10792
rect 26568 10752 26574 10764
rect 27341 10761 27353 10764
rect 27387 10761 27399 10795
rect 27341 10755 27399 10761
rect 2498 10684 2504 10736
rect 2556 10724 2562 10736
rect 2685 10727 2743 10733
rect 2685 10724 2697 10727
rect 2556 10696 2697 10724
rect 2556 10684 2562 10696
rect 2685 10693 2697 10696
rect 2731 10693 2743 10727
rect 2685 10687 2743 10693
rect 6730 10684 6736 10736
rect 6788 10724 6794 10736
rect 9125 10727 9183 10733
rect 9125 10724 9137 10727
rect 6788 10696 9137 10724
rect 6788 10684 6794 10696
rect 9125 10693 9137 10696
rect 9171 10724 9183 10727
rect 9582 10724 9588 10736
rect 9171 10696 9588 10724
rect 9171 10693 9183 10696
rect 9125 10687 9183 10693
rect 9582 10684 9588 10696
rect 9640 10684 9646 10736
rect 13814 10684 13820 10736
rect 13872 10724 13878 10736
rect 14277 10727 14335 10733
rect 14277 10724 14289 10727
rect 13872 10696 14289 10724
rect 13872 10684 13878 10696
rect 14277 10693 14289 10696
rect 14323 10693 14335 10727
rect 15841 10727 15899 10733
rect 15841 10724 15853 10727
rect 14277 10687 14335 10693
rect 14660 10696 15853 10724
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 7653 10659 7711 10665
rect 7653 10656 7665 10659
rect 7616 10628 7665 10656
rect 7616 10616 7622 10628
rect 7653 10625 7665 10628
rect 7699 10656 7711 10659
rect 8294 10656 8300 10668
rect 7699 10628 8300 10656
rect 7699 10625 7711 10628
rect 7653 10619 7711 10625
rect 8294 10616 8300 10628
rect 8352 10656 8358 10668
rect 9493 10659 9551 10665
rect 9493 10656 9505 10659
rect 8352 10628 9505 10656
rect 8352 10616 8358 10628
rect 9493 10625 9505 10628
rect 9539 10656 9551 10659
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 9539 10628 10609 10656
rect 9539 10625 9551 10628
rect 9493 10619 9551 10625
rect 10597 10625 10609 10628
rect 10643 10656 10655 10659
rect 10686 10656 10692 10668
rect 10643 10628 10692 10656
rect 10643 10625 10655 10628
rect 10597 10619 10655 10625
rect 10686 10616 10692 10628
rect 10744 10656 10750 10668
rect 11882 10656 11888 10668
rect 10744 10628 11888 10656
rect 10744 10616 10750 10628
rect 11882 10616 11888 10628
rect 11940 10616 11946 10668
rect 1394 10588 1400 10600
rect 1355 10560 1400 10588
rect 1394 10548 1400 10560
rect 1452 10548 1458 10600
rect 3050 10588 3056 10600
rect 3011 10560 3056 10588
rect 3050 10548 3056 10560
rect 3108 10548 3114 10600
rect 3142 10548 3148 10600
rect 3200 10588 3206 10600
rect 3309 10591 3367 10597
rect 3309 10588 3321 10591
rect 3200 10560 3321 10588
rect 3200 10548 3206 10560
rect 3309 10557 3321 10560
rect 3355 10557 3367 10591
rect 3309 10551 3367 10557
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10588 6699 10591
rect 7466 10588 7472 10600
rect 6687 10560 7472 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 7466 10548 7472 10560
rect 7524 10548 7530 10600
rect 14458 10548 14464 10600
rect 14516 10588 14522 10600
rect 14660 10597 14688 10696
rect 15841 10693 15853 10696
rect 15887 10693 15899 10727
rect 15841 10687 15899 10693
rect 14918 10656 14924 10668
rect 14879 10628 14924 10656
rect 14918 10616 14924 10628
rect 14976 10616 14982 10668
rect 15378 10616 15384 10668
rect 15436 10656 15442 10668
rect 16298 10656 16304 10668
rect 15436 10628 16304 10656
rect 15436 10616 15442 10628
rect 16298 10616 16304 10628
rect 16356 10656 16362 10668
rect 16393 10659 16451 10665
rect 16393 10656 16405 10659
rect 16356 10628 16405 10656
rect 16356 10616 16362 10628
rect 16393 10625 16405 10628
rect 16439 10625 16451 10659
rect 19426 10656 19432 10668
rect 19387 10628 19432 10656
rect 16393 10619 16451 10625
rect 19426 10616 19432 10628
rect 19484 10616 19490 10668
rect 14645 10591 14703 10597
rect 14645 10588 14657 10591
rect 14516 10560 14657 10588
rect 14516 10548 14522 10560
rect 14645 10557 14657 10560
rect 14691 10557 14703 10591
rect 14645 10551 14703 10557
rect 15286 10548 15292 10600
rect 15344 10588 15350 10600
rect 16209 10591 16267 10597
rect 16209 10588 16221 10591
rect 15344 10560 16221 10588
rect 15344 10548 15350 10560
rect 16209 10557 16221 10560
rect 16255 10557 16267 10591
rect 16209 10551 16267 10557
rect 18417 10591 18475 10597
rect 18417 10557 18429 10591
rect 18463 10588 18475 10591
rect 18463 10560 19288 10588
rect 18463 10557 18475 10560
rect 18417 10551 18475 10557
rect 5905 10523 5963 10529
rect 5905 10489 5917 10523
rect 5951 10520 5963 10523
rect 7006 10520 7012 10532
rect 5951 10492 7012 10520
rect 5951 10489 5963 10492
rect 5905 10483 5963 10489
rect 7006 10480 7012 10492
rect 7064 10480 7070 10532
rect 10042 10480 10048 10532
rect 10100 10520 10106 10532
rect 10505 10523 10563 10529
rect 10505 10520 10517 10523
rect 10100 10492 10517 10520
rect 10100 10480 10106 10492
rect 10505 10489 10517 10492
rect 10551 10520 10563 10523
rect 10594 10520 10600 10532
rect 10551 10492 10600 10520
rect 10551 10489 10563 10492
rect 10505 10483 10563 10489
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 13817 10523 13875 10529
rect 13817 10489 13829 10523
rect 13863 10520 13875 10523
rect 14734 10520 14740 10532
rect 13863 10492 14740 10520
rect 13863 10489 13875 10492
rect 13817 10483 13875 10489
rect 14734 10480 14740 10492
rect 14792 10480 14798 10532
rect 15749 10523 15807 10529
rect 15749 10489 15761 10523
rect 15795 10520 15807 10523
rect 16301 10523 16359 10529
rect 16301 10520 16313 10523
rect 15795 10492 16313 10520
rect 15795 10489 15807 10492
rect 15749 10483 15807 10489
rect 16301 10489 16313 10492
rect 16347 10520 16359 10523
rect 16390 10520 16396 10532
rect 16347 10492 16396 10520
rect 16347 10489 16359 10492
rect 16301 10483 16359 10489
rect 16390 10480 16396 10492
rect 16448 10480 16454 10532
rect 17865 10523 17923 10529
rect 17865 10489 17877 10523
rect 17911 10520 17923 10523
rect 18782 10520 18788 10532
rect 17911 10492 18788 10520
rect 17911 10489 17923 10492
rect 17865 10483 17923 10489
rect 18782 10480 18788 10492
rect 18840 10480 18846 10532
rect 19260 10529 19288 10560
rect 23842 10548 23848 10600
rect 23900 10588 23906 10600
rect 26421 10591 26479 10597
rect 26421 10588 26433 10591
rect 23900 10560 26433 10588
rect 23900 10548 23906 10560
rect 26421 10557 26433 10560
rect 26467 10588 26479 10591
rect 26973 10591 27031 10597
rect 26973 10588 26985 10591
rect 26467 10560 26985 10588
rect 26467 10557 26479 10560
rect 26421 10551 26479 10557
rect 26973 10557 26985 10560
rect 27019 10557 27031 10591
rect 27522 10588 27528 10600
rect 27483 10560 27528 10588
rect 26973 10551 27031 10557
rect 27522 10548 27528 10560
rect 27580 10588 27586 10600
rect 28077 10591 28135 10597
rect 28077 10588 28089 10591
rect 27580 10560 28089 10588
rect 27580 10548 27586 10560
rect 28077 10557 28089 10560
rect 28123 10557 28135 10591
rect 28077 10551 28135 10557
rect 19245 10523 19303 10529
rect 19245 10489 19257 10523
rect 19291 10520 19303 10523
rect 19518 10520 19524 10532
rect 19291 10492 19524 10520
rect 19291 10489 19303 10492
rect 19245 10483 19303 10489
rect 19518 10480 19524 10492
rect 19576 10480 19582 10532
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 4430 10452 4436 10464
rect 4391 10424 4436 10452
rect 4430 10412 4436 10424
rect 4488 10412 4494 10464
rect 6270 10452 6276 10464
rect 6231 10424 6276 10452
rect 6270 10412 6276 10424
rect 6328 10412 6334 10464
rect 7561 10455 7619 10461
rect 7561 10421 7573 10455
rect 7607 10452 7619 10455
rect 7834 10452 7840 10464
rect 7607 10424 7840 10452
rect 7607 10421 7619 10424
rect 7561 10415 7619 10421
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 9858 10452 9864 10464
rect 9819 10424 9864 10452
rect 9858 10412 9864 10424
rect 9916 10452 9922 10464
rect 10413 10455 10471 10461
rect 10413 10452 10425 10455
rect 9916 10424 10425 10452
rect 9916 10412 9922 10424
rect 10413 10421 10425 10424
rect 10459 10421 10471 10455
rect 10413 10415 10471 10421
rect 13081 10455 13139 10461
rect 13081 10421 13093 10455
rect 13127 10452 13139 10455
rect 13262 10452 13268 10464
rect 13127 10424 13268 10452
rect 13127 10421 13139 10424
rect 13081 10415 13139 10421
rect 13262 10412 13268 10424
rect 13320 10412 13326 10464
rect 18693 10455 18751 10461
rect 18693 10421 18705 10455
rect 18739 10452 18751 10455
rect 19150 10452 19156 10464
rect 18739 10424 19156 10452
rect 18739 10421 18751 10424
rect 18693 10415 18751 10421
rect 19150 10412 19156 10424
rect 19208 10452 19214 10464
rect 19337 10455 19395 10461
rect 19337 10452 19349 10455
rect 19208 10424 19349 10452
rect 19208 10412 19214 10424
rect 19337 10421 19349 10424
rect 19383 10421 19395 10455
rect 22462 10452 22468 10464
rect 22423 10424 22468 10452
rect 19337 10415 19395 10421
rect 22462 10412 22468 10424
rect 22520 10412 22526 10464
rect 23474 10412 23480 10464
rect 23532 10452 23538 10464
rect 23661 10455 23719 10461
rect 23661 10452 23673 10455
rect 23532 10424 23673 10452
rect 23532 10412 23538 10424
rect 23661 10421 23673 10424
rect 23707 10421 23719 10455
rect 26602 10452 26608 10464
rect 26563 10424 26608 10452
rect 23661 10415 23719 10421
rect 26602 10412 26608 10424
rect 26660 10412 26666 10464
rect 27706 10452 27712 10464
rect 27667 10424 27712 10452
rect 27706 10412 27712 10424
rect 27764 10412 27770 10464
rect 1104 10362 28888 10384
rect 1104 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 20982 10362
rect 21034 10310 21046 10362
rect 21098 10310 21110 10362
rect 21162 10310 21174 10362
rect 21226 10310 28888 10362
rect 1104 10288 28888 10310
rect 2038 10248 2044 10260
rect 1999 10220 2044 10248
rect 2038 10208 2044 10220
rect 2096 10208 2102 10260
rect 2130 10208 2136 10260
rect 2188 10248 2194 10260
rect 2593 10251 2651 10257
rect 2593 10248 2605 10251
rect 2188 10220 2605 10248
rect 2188 10208 2194 10220
rect 2593 10217 2605 10220
rect 2639 10217 2651 10251
rect 3142 10248 3148 10260
rect 3103 10220 3148 10248
rect 2593 10211 2651 10217
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 6641 10251 6699 10257
rect 6641 10217 6653 10251
rect 6687 10248 6699 10251
rect 6730 10248 6736 10260
rect 6687 10220 6736 10248
rect 6687 10217 6699 10220
rect 6641 10211 6699 10217
rect 6730 10208 6736 10220
rect 6788 10208 6794 10260
rect 6914 10248 6920 10260
rect 6875 10220 6920 10248
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7193 10251 7251 10257
rect 7193 10248 7205 10251
rect 7064 10220 7205 10248
rect 7064 10208 7070 10220
rect 7193 10217 7205 10220
rect 7239 10217 7251 10251
rect 11882 10248 11888 10260
rect 11843 10220 11888 10248
rect 7193 10211 7251 10217
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 14734 10208 14740 10260
rect 14792 10248 14798 10260
rect 15289 10251 15347 10257
rect 15289 10248 15301 10251
rect 14792 10220 15301 10248
rect 14792 10208 14798 10220
rect 15289 10217 15301 10220
rect 15335 10217 15347 10251
rect 16298 10248 16304 10260
rect 16259 10220 16304 10248
rect 15289 10211 15347 10217
rect 16298 10208 16304 10220
rect 16356 10208 16362 10260
rect 16850 10248 16856 10260
rect 16811 10220 16856 10248
rect 16850 10208 16856 10220
rect 16908 10208 16914 10260
rect 17218 10248 17224 10260
rect 17179 10220 17224 10248
rect 17218 10208 17224 10220
rect 17276 10208 17282 10260
rect 18414 10248 18420 10260
rect 18375 10220 18420 10248
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 18782 10248 18788 10260
rect 18743 10220 18788 10248
rect 18782 10208 18788 10220
rect 18840 10208 18846 10260
rect 19058 10208 19064 10260
rect 19116 10248 19122 10260
rect 19153 10251 19211 10257
rect 19153 10248 19165 10251
rect 19116 10220 19165 10248
rect 19116 10208 19122 10220
rect 19153 10217 19165 10220
rect 19199 10217 19211 10251
rect 19153 10211 19211 10217
rect 22462 10208 22468 10260
rect 22520 10248 22526 10260
rect 22741 10251 22799 10257
rect 22741 10248 22753 10251
rect 22520 10220 22753 10248
rect 22520 10208 22526 10220
rect 22741 10217 22753 10220
rect 22787 10217 22799 10251
rect 22741 10211 22799 10217
rect 23474 10208 23480 10260
rect 23532 10248 23538 10260
rect 24213 10251 24271 10257
rect 24213 10248 24225 10251
rect 23532 10220 24225 10248
rect 23532 10208 23538 10220
rect 24213 10217 24225 10220
rect 24259 10217 24271 10251
rect 24213 10211 24271 10217
rect 1762 10140 1768 10192
rect 1820 10180 1826 10192
rect 1949 10183 2007 10189
rect 1949 10180 1961 10183
rect 1820 10152 1961 10180
rect 1820 10140 1826 10152
rect 1949 10149 1961 10152
rect 1995 10149 2007 10183
rect 1949 10143 2007 10149
rect 3050 10140 3056 10192
rect 3108 10180 3114 10192
rect 3421 10183 3479 10189
rect 3421 10180 3433 10183
rect 3108 10152 3433 10180
rect 3108 10140 3114 10152
rect 3421 10149 3433 10152
rect 3467 10180 3479 10183
rect 3602 10180 3608 10192
rect 3467 10152 3608 10180
rect 3467 10149 3479 10152
rect 3421 10143 3479 10149
rect 3602 10140 3608 10152
rect 3660 10140 3666 10192
rect 5534 10140 5540 10192
rect 5592 10180 5598 10192
rect 7466 10180 7472 10192
rect 5592 10152 7472 10180
rect 5592 10140 5598 10152
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 7561 10183 7619 10189
rect 7561 10149 7573 10183
rect 7607 10180 7619 10183
rect 7742 10180 7748 10192
rect 7607 10152 7748 10180
rect 7607 10149 7619 10152
rect 7561 10143 7619 10149
rect 7742 10140 7748 10152
rect 7800 10140 7806 10192
rect 9401 10183 9459 10189
rect 9401 10149 9413 10183
rect 9447 10180 9459 10183
rect 10686 10180 10692 10192
rect 9447 10152 10692 10180
rect 9447 10149 9459 10152
rect 9401 10143 9459 10149
rect 10686 10140 10692 10152
rect 10744 10189 10750 10192
rect 10744 10183 10808 10189
rect 10744 10149 10762 10183
rect 10796 10149 10808 10183
rect 10744 10143 10808 10149
rect 10744 10140 10750 10143
rect 13630 10140 13636 10192
rect 13688 10180 13694 10192
rect 13909 10183 13967 10189
rect 13909 10180 13921 10183
rect 13688 10152 13921 10180
rect 13688 10140 13694 10152
rect 13909 10149 13921 10152
rect 13955 10180 13967 10183
rect 15102 10180 15108 10192
rect 13955 10152 15108 10180
rect 13955 10149 13967 10152
rect 13909 10143 13967 10149
rect 15102 10140 15108 10152
rect 15160 10140 15166 10192
rect 18230 10140 18236 10192
rect 18288 10180 18294 10192
rect 19076 10180 19104 10208
rect 18288 10152 19104 10180
rect 18288 10140 18294 10152
rect 24118 10140 24124 10192
rect 24176 10180 24182 10192
rect 24305 10183 24363 10189
rect 24305 10180 24317 10183
rect 24176 10152 24317 10180
rect 24176 10140 24182 10152
rect 24305 10149 24317 10152
rect 24351 10149 24363 10183
rect 24305 10143 24363 10149
rect 24854 10140 24860 10192
rect 24912 10180 24918 10192
rect 27430 10180 27436 10192
rect 24912 10152 27436 10180
rect 24912 10140 24918 10152
rect 27430 10140 27436 10152
rect 27488 10140 27494 10192
rect 8846 10072 8852 10124
rect 8904 10112 8910 10124
rect 8941 10115 8999 10121
rect 8941 10112 8953 10115
rect 8904 10084 8953 10112
rect 8904 10072 8910 10084
rect 8941 10081 8953 10084
rect 8987 10081 8999 10115
rect 13814 10112 13820 10124
rect 13775 10084 13820 10112
rect 8941 10075 8999 10081
rect 13814 10072 13820 10084
rect 13872 10072 13878 10124
rect 15654 10112 15660 10124
rect 15615 10084 15660 10112
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 16482 10112 16488 10124
rect 15764 10084 16488 10112
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10044 2283 10047
rect 2314 10044 2320 10056
rect 2271 10016 2320 10044
rect 2271 10013 2283 10016
rect 2225 10007 2283 10013
rect 2314 10004 2320 10016
rect 2372 10004 2378 10056
rect 7650 10044 7656 10056
rect 7611 10016 7656 10044
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 6270 9936 6276 9988
rect 6328 9976 6334 9988
rect 7558 9976 7564 9988
rect 6328 9948 7564 9976
rect 6328 9936 6334 9948
rect 7558 9936 7564 9948
rect 7616 9976 7622 9988
rect 7760 9976 7788 10007
rect 10410 10004 10416 10056
rect 10468 10044 10474 10056
rect 10505 10047 10563 10053
rect 10505 10044 10517 10047
rect 10468 10016 10517 10044
rect 10468 10004 10474 10016
rect 10505 10013 10517 10016
rect 10551 10013 10563 10047
rect 13998 10044 14004 10056
rect 13959 10016 14004 10044
rect 10505 10007 10563 10013
rect 13998 10004 14004 10016
rect 14056 10004 14062 10056
rect 15562 10004 15568 10056
rect 15620 10044 15626 10056
rect 15764 10053 15792 10084
rect 16482 10072 16488 10084
rect 16540 10072 16546 10124
rect 18598 10072 18604 10124
rect 18656 10112 18662 10124
rect 18782 10112 18788 10124
rect 18656 10084 18788 10112
rect 18656 10072 18662 10084
rect 18782 10072 18788 10084
rect 18840 10112 18846 10124
rect 19245 10115 19303 10121
rect 19245 10112 19257 10115
rect 18840 10084 19257 10112
rect 18840 10072 18846 10084
rect 19245 10081 19257 10084
rect 19291 10081 19303 10115
rect 20530 10112 20536 10124
rect 20491 10084 20536 10112
rect 19245 10075 19303 10081
rect 20530 10072 20536 10084
rect 20588 10072 20594 10124
rect 21450 10072 21456 10124
rect 21508 10112 21514 10124
rect 21617 10115 21675 10121
rect 21617 10112 21629 10115
rect 21508 10084 21629 10112
rect 21508 10072 21514 10084
rect 21617 10081 21629 10084
rect 21663 10081 21675 10115
rect 21617 10075 21675 10081
rect 26418 10072 26424 10124
rect 26476 10112 26482 10124
rect 26513 10115 26571 10121
rect 26513 10112 26525 10115
rect 26476 10084 26525 10112
rect 26476 10072 26482 10084
rect 26513 10081 26525 10084
rect 26559 10081 26571 10115
rect 26513 10075 26571 10081
rect 15749 10047 15807 10053
rect 15749 10044 15761 10047
rect 15620 10016 15761 10044
rect 15620 10004 15626 10016
rect 15749 10013 15761 10016
rect 15795 10013 15807 10047
rect 15749 10007 15807 10013
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10044 15991 10047
rect 16298 10044 16304 10056
rect 15979 10016 16304 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 16298 10004 16304 10016
rect 16356 10004 16362 10056
rect 19426 10044 19432 10056
rect 19387 10016 19432 10044
rect 19426 10004 19432 10016
rect 19484 10004 19490 10056
rect 20806 10004 20812 10056
rect 20864 10044 20870 10056
rect 21358 10044 21364 10056
rect 20864 10016 21364 10044
rect 20864 10004 20870 10016
rect 21358 10004 21364 10016
rect 21416 10004 21422 10056
rect 24210 10004 24216 10056
rect 24268 10044 24274 10056
rect 24397 10047 24455 10053
rect 24397 10044 24409 10047
rect 24268 10016 24409 10044
rect 24268 10004 24274 10016
rect 24397 10013 24409 10016
rect 24443 10013 24455 10047
rect 24397 10007 24455 10013
rect 7616 9948 7788 9976
rect 7616 9936 7622 9948
rect 23290 9936 23296 9988
rect 23348 9976 23354 9988
rect 23845 9979 23903 9985
rect 23845 9976 23857 9979
rect 23348 9948 23857 9976
rect 23348 9936 23354 9948
rect 23845 9945 23857 9948
rect 23891 9945 23903 9979
rect 23845 9939 23903 9945
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 1670 9908 1676 9920
rect 1627 9880 1676 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 1670 9868 1676 9880
rect 1728 9868 1734 9920
rect 5166 9868 5172 9920
rect 5224 9908 5230 9920
rect 8110 9908 8116 9920
rect 5224 9880 8116 9908
rect 5224 9868 5230 9880
rect 8110 9868 8116 9880
rect 8168 9868 8174 9920
rect 8297 9911 8355 9917
rect 8297 9877 8309 9911
rect 8343 9908 8355 9911
rect 8386 9908 8392 9920
rect 8343 9880 8392 9908
rect 8343 9877 8355 9880
rect 8297 9871 8355 9877
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 8478 9868 8484 9920
rect 8536 9908 8542 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 8536 9880 8769 9908
rect 8536 9868 8542 9880
rect 8757 9877 8769 9880
rect 8803 9908 8815 9911
rect 9582 9908 9588 9920
rect 8803 9880 9588 9908
rect 8803 9877 8815 9880
rect 8757 9871 8815 9877
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 10042 9908 10048 9920
rect 10003 9880 10048 9908
rect 10042 9868 10048 9880
rect 10100 9868 10106 9920
rect 13262 9908 13268 9920
rect 13223 9880 13268 9908
rect 13262 9868 13268 9880
rect 13320 9868 13326 9920
rect 13449 9911 13507 9917
rect 13449 9877 13461 9911
rect 13495 9908 13507 9911
rect 13722 9908 13728 9920
rect 13495 9880 13728 9908
rect 13495 9877 13507 9880
rect 13449 9871 13507 9877
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 20346 9908 20352 9920
rect 20307 9880 20352 9908
rect 20346 9868 20352 9880
rect 20404 9868 20410 9920
rect 23753 9911 23811 9917
rect 23753 9877 23765 9911
rect 23799 9908 23811 9911
rect 24026 9908 24032 9920
rect 23799 9880 24032 9908
rect 23799 9877 23811 9880
rect 23753 9871 23811 9877
rect 24026 9868 24032 9880
rect 24084 9908 24090 9920
rect 24394 9908 24400 9920
rect 24084 9880 24400 9908
rect 24084 9868 24090 9880
rect 24394 9868 24400 9880
rect 24452 9868 24458 9920
rect 26694 9908 26700 9920
rect 26655 9880 26700 9908
rect 26694 9868 26700 9880
rect 26752 9868 26758 9920
rect 1104 9818 28888 9840
rect 1104 9766 5982 9818
rect 6034 9766 6046 9818
rect 6098 9766 6110 9818
rect 6162 9766 6174 9818
rect 6226 9766 15982 9818
rect 16034 9766 16046 9818
rect 16098 9766 16110 9818
rect 16162 9766 16174 9818
rect 16226 9766 25982 9818
rect 26034 9766 26046 9818
rect 26098 9766 26110 9818
rect 26162 9766 26174 9818
rect 26226 9766 28888 9818
rect 1104 9744 28888 9766
rect 2314 9704 2320 9716
rect 2275 9676 2320 9704
rect 2314 9664 2320 9676
rect 2372 9664 2378 9716
rect 3602 9704 3608 9716
rect 3563 9676 3608 9704
rect 3602 9664 3608 9676
rect 3660 9664 3666 9716
rect 6270 9664 6276 9716
rect 6328 9704 6334 9716
rect 6549 9707 6607 9713
rect 6549 9704 6561 9707
rect 6328 9676 6561 9704
rect 6328 9664 6334 9676
rect 6549 9673 6561 9676
rect 6595 9673 6607 9707
rect 6549 9667 6607 9673
rect 7650 9664 7656 9716
rect 7708 9704 7714 9716
rect 7745 9707 7803 9713
rect 7745 9704 7757 9707
rect 7708 9676 7757 9704
rect 7708 9664 7714 9676
rect 7745 9673 7757 9676
rect 7791 9673 7803 9707
rect 7745 9667 7803 9673
rect 7834 9664 7840 9716
rect 7892 9704 7898 9716
rect 13814 9704 13820 9716
rect 7892 9676 8340 9704
rect 7892 9664 7898 9676
rect 2332 9568 2360 9664
rect 2866 9596 2872 9648
rect 2924 9636 2930 9648
rect 2958 9636 2964 9648
rect 2924 9608 2964 9636
rect 2924 9596 2930 9608
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 3142 9636 3148 9648
rect 3103 9608 3148 9636
rect 3142 9596 3148 9608
rect 3200 9596 3206 9648
rect 8312 9636 8340 9676
rect 13188 9676 13820 9704
rect 9309 9639 9367 9645
rect 9309 9636 9321 9639
rect 8312 9608 9321 9636
rect 9309 9605 9321 9608
rect 9355 9605 9367 9639
rect 9309 9599 9367 9605
rect 12713 9639 12771 9645
rect 12713 9605 12725 9639
rect 12759 9636 12771 9639
rect 13188 9636 13216 9676
rect 13814 9664 13820 9676
rect 13872 9664 13878 9716
rect 15381 9707 15439 9713
rect 15381 9673 15393 9707
rect 15427 9704 15439 9707
rect 15654 9704 15660 9716
rect 15427 9676 15660 9704
rect 15427 9673 15439 9676
rect 15381 9667 15439 9673
rect 15654 9664 15660 9676
rect 15712 9664 15718 9716
rect 16117 9707 16175 9713
rect 16117 9673 16129 9707
rect 16163 9704 16175 9707
rect 16298 9704 16304 9716
rect 16163 9676 16304 9704
rect 16163 9673 16175 9676
rect 16117 9667 16175 9673
rect 16298 9664 16304 9676
rect 16356 9664 16362 9716
rect 20441 9707 20499 9713
rect 20441 9673 20453 9707
rect 20487 9704 20499 9707
rect 20530 9704 20536 9716
rect 20487 9676 20536 9704
rect 20487 9673 20499 9676
rect 20441 9667 20499 9673
rect 20530 9664 20536 9676
rect 20588 9664 20594 9716
rect 24118 9664 24124 9716
rect 24176 9704 24182 9716
rect 24673 9707 24731 9713
rect 24673 9704 24685 9707
rect 24176 9676 24685 9704
rect 24176 9664 24182 9676
rect 24673 9673 24685 9676
rect 24719 9673 24731 9707
rect 24673 9667 24731 9673
rect 26510 9664 26516 9716
rect 26568 9704 26574 9716
rect 27525 9707 27583 9713
rect 27525 9704 27537 9707
rect 26568 9676 27537 9704
rect 26568 9664 26574 9676
rect 27525 9673 27537 9676
rect 27571 9673 27583 9707
rect 27525 9667 27583 9673
rect 12759 9608 13216 9636
rect 12759 9605 12771 9608
rect 12713 9599 12771 9605
rect 18690 9596 18696 9648
rect 18748 9636 18754 9648
rect 18785 9639 18843 9645
rect 18785 9636 18797 9639
rect 18748 9608 18797 9636
rect 18748 9596 18754 9608
rect 18785 9605 18797 9608
rect 18831 9605 18843 9639
rect 23661 9639 23719 9645
rect 23661 9636 23673 9639
rect 18785 9599 18843 9605
rect 22480 9608 23673 9636
rect 4065 9571 4123 9577
rect 4065 9568 4077 9571
rect 2332 9540 4077 9568
rect 4065 9537 4077 9540
rect 4111 9568 4123 9571
rect 4111 9540 4292 9568
rect 4111 9537 4123 9540
rect 4065 9531 4123 9537
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 2501 9503 2559 9509
rect 1443 9472 2084 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 2056 9441 2084 9472
rect 2501 9469 2513 9503
rect 2547 9500 2559 9503
rect 3142 9500 3148 9512
rect 2547 9472 3148 9500
rect 2547 9469 2559 9472
rect 2501 9463 2559 9469
rect 3142 9460 3148 9472
rect 3200 9460 3206 9512
rect 3602 9460 3608 9512
rect 3660 9500 3666 9512
rect 4157 9503 4215 9509
rect 4157 9500 4169 9503
rect 3660 9472 4169 9500
rect 3660 9460 3666 9472
rect 4157 9469 4169 9472
rect 4203 9469 4215 9503
rect 4264 9500 4292 9540
rect 7190 9528 7196 9580
rect 7248 9568 7254 9580
rect 7285 9571 7343 9577
rect 7285 9568 7297 9571
rect 7248 9540 7297 9568
rect 7248 9528 7254 9540
rect 7285 9537 7297 9540
rect 7331 9568 7343 9571
rect 8018 9568 8024 9580
rect 7331 9540 8024 9568
rect 7331 9537 7343 9540
rect 7285 9531 7343 9537
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 8294 9568 8300 9580
rect 8255 9540 8300 9568
rect 8294 9528 8300 9540
rect 8352 9528 8358 9580
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9568 10011 9571
rect 10686 9568 10692 9580
rect 9999 9540 10692 9568
rect 9999 9537 10011 9540
rect 9953 9531 10011 9537
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 19426 9568 19432 9580
rect 19339 9540 19432 9568
rect 19426 9528 19432 9540
rect 19484 9568 19490 9580
rect 19484 9540 19656 9568
rect 19484 9528 19490 9540
rect 4430 9509 4436 9512
rect 4424 9500 4436 9509
rect 4264 9472 4436 9500
rect 4157 9463 4215 9469
rect 4424 9463 4436 9472
rect 2041 9435 2099 9441
rect 2041 9401 2053 9435
rect 2087 9432 2099 9435
rect 2958 9432 2964 9444
rect 2087 9404 2964 9432
rect 2087 9401 2099 9404
rect 2041 9395 2099 9401
rect 2958 9392 2964 9404
rect 3016 9392 3022 9444
rect 4172 9432 4200 9463
rect 4430 9460 4436 9463
rect 4488 9460 4494 9512
rect 7374 9460 7380 9512
rect 7432 9500 7438 9512
rect 8205 9503 8263 9509
rect 8205 9500 8217 9503
rect 7432 9472 8217 9500
rect 7432 9460 7438 9472
rect 5350 9432 5356 9444
rect 4172 9404 5356 9432
rect 5350 9392 5356 9404
rect 5408 9392 5414 9444
rect 7576 9376 7604 9472
rect 8205 9469 8217 9472
rect 8251 9469 8263 9503
rect 8205 9463 8263 9469
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9500 9275 9503
rect 9858 9500 9864 9512
rect 9263 9472 9864 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 9858 9460 9864 9472
rect 9916 9460 9922 9512
rect 12434 9460 12440 9512
rect 12492 9500 12498 9512
rect 13173 9503 13231 9509
rect 13173 9500 13185 9503
rect 12492 9472 13185 9500
rect 12492 9460 12498 9472
rect 13173 9469 13185 9472
rect 13219 9500 13231 9503
rect 13262 9500 13268 9512
rect 13219 9472 13268 9500
rect 13219 9469 13231 9472
rect 13173 9463 13231 9469
rect 13262 9460 13268 9472
rect 13320 9460 13326 9512
rect 19153 9503 19211 9509
rect 19153 9469 19165 9503
rect 19199 9500 19211 9503
rect 19242 9500 19248 9512
rect 19199 9472 19248 9500
rect 19199 9469 19211 9472
rect 19153 9463 19211 9469
rect 19242 9460 19248 9472
rect 19300 9460 19306 9512
rect 19628 9444 19656 9540
rect 22186 9528 22192 9580
rect 22244 9568 22250 9580
rect 22480 9577 22508 9608
rect 23661 9605 23673 9608
rect 23707 9605 23719 9639
rect 23661 9599 23719 9605
rect 23934 9596 23940 9648
rect 23992 9636 23998 9648
rect 24302 9636 24308 9648
rect 23992 9608 24308 9636
rect 23992 9596 23998 9608
rect 24302 9596 24308 9608
rect 24360 9596 24366 9648
rect 24486 9636 24492 9648
rect 24447 9608 24492 9636
rect 24486 9596 24492 9608
rect 24544 9596 24550 9648
rect 24578 9596 24584 9648
rect 24636 9636 24642 9648
rect 24946 9636 24952 9648
rect 24636 9608 24952 9636
rect 24636 9596 24642 9608
rect 24946 9596 24952 9608
rect 25004 9596 25010 9648
rect 26970 9636 26976 9648
rect 26931 9608 26976 9636
rect 26970 9596 26976 9608
rect 27028 9596 27034 9648
rect 22465 9571 22523 9577
rect 22465 9568 22477 9571
rect 22244 9540 22477 9568
rect 22244 9528 22250 9540
rect 22465 9537 22477 9540
rect 22511 9537 22523 9571
rect 22465 9531 22523 9537
rect 22554 9528 22560 9580
rect 22612 9568 22618 9580
rect 23109 9571 23167 9577
rect 22612 9540 22657 9568
rect 22612 9528 22618 9540
rect 23109 9537 23121 9571
rect 23155 9568 23167 9571
rect 23382 9568 23388 9580
rect 23155 9540 23388 9568
rect 23155 9537 23167 9540
rect 23109 9531 23167 9537
rect 23382 9528 23388 9540
rect 23440 9528 23446 9580
rect 23477 9571 23535 9577
rect 23477 9537 23489 9571
rect 23523 9568 23535 9571
rect 23566 9568 23572 9580
rect 23523 9540 23572 9568
rect 23523 9537 23535 9540
rect 23477 9531 23535 9537
rect 23566 9528 23572 9540
rect 23624 9568 23630 9580
rect 24210 9568 24216 9580
rect 23624 9540 24072 9568
rect 24123 9540 24216 9568
rect 23624 9528 23630 9540
rect 20622 9460 20628 9512
rect 20680 9500 20686 9512
rect 22373 9503 22431 9509
rect 20680 9472 21956 9500
rect 20680 9460 20686 9472
rect 7742 9392 7748 9444
rect 7800 9432 7806 9444
rect 8757 9435 8815 9441
rect 8757 9432 8769 9435
rect 7800 9404 8769 9432
rect 7800 9392 7806 9404
rect 8757 9401 8769 9404
rect 8803 9401 8815 9435
rect 9950 9432 9956 9444
rect 8757 9395 8815 9401
rect 9692 9404 9956 9432
rect 9692 9376 9720 9404
rect 9950 9392 9956 9404
rect 10008 9392 10014 9444
rect 10410 9392 10416 9444
rect 10468 9432 10474 9444
rect 10873 9435 10931 9441
rect 10873 9432 10885 9435
rect 10468 9404 10885 9432
rect 10468 9392 10474 9404
rect 10873 9401 10885 9404
rect 10919 9401 10931 9435
rect 10873 9395 10931 9401
rect 13440 9435 13498 9441
rect 13440 9401 13452 9435
rect 13486 9432 13498 9435
rect 13538 9432 13544 9444
rect 13486 9404 13544 9432
rect 13486 9401 13498 9404
rect 13440 9395 13498 9401
rect 13538 9392 13544 9404
rect 13596 9392 13602 9444
rect 19610 9392 19616 9444
rect 19668 9432 19674 9444
rect 21928 9441 21956 9472
rect 22373 9469 22385 9503
rect 22419 9500 22431 9503
rect 22646 9500 22652 9512
rect 22419 9472 22652 9500
rect 22419 9469 22431 9472
rect 22373 9463 22431 9469
rect 22646 9460 22652 9472
rect 22704 9500 22710 9512
rect 23290 9500 23296 9512
rect 22704 9472 23296 9500
rect 22704 9460 22710 9472
rect 23290 9460 23296 9472
rect 23348 9460 23354 9512
rect 24044 9509 24072 9540
rect 24210 9528 24216 9540
rect 24268 9568 24274 9580
rect 24268 9540 25176 9568
rect 24268 9528 24274 9540
rect 24029 9503 24087 9509
rect 24029 9469 24041 9503
rect 24075 9469 24087 9503
rect 24029 9463 24087 9469
rect 19889 9435 19947 9441
rect 19889 9432 19901 9435
rect 19668 9404 19901 9432
rect 19668 9392 19674 9404
rect 19889 9401 19901 9404
rect 19935 9432 19947 9435
rect 21913 9435 21971 9441
rect 19935 9404 21496 9432
rect 19935 9401 19947 9404
rect 19889 9395 19947 9401
rect 21468 9376 21496 9404
rect 21913 9401 21925 9435
rect 21959 9432 21971 9435
rect 22554 9432 22560 9444
rect 21959 9404 22560 9432
rect 21959 9401 21971 9404
rect 21913 9395 21971 9401
rect 22554 9392 22560 9404
rect 22612 9392 22618 9444
rect 23842 9392 23848 9444
rect 23900 9432 23906 9444
rect 25148 9441 25176 9540
rect 25593 9503 25651 9509
rect 25593 9469 25605 9503
rect 25639 9500 25651 9503
rect 25682 9500 25688 9512
rect 25639 9472 25688 9500
rect 25639 9469 25651 9472
rect 25593 9463 25651 9469
rect 25682 9460 25688 9472
rect 25740 9460 25746 9512
rect 24489 9435 24547 9441
rect 24489 9432 24501 9435
rect 23900 9404 24501 9432
rect 23900 9392 23906 9404
rect 24489 9401 24501 9404
rect 24535 9401 24547 9435
rect 24489 9395 24547 9401
rect 25133 9435 25191 9441
rect 25133 9401 25145 9435
rect 25179 9432 25191 9435
rect 25501 9435 25559 9441
rect 25501 9432 25513 9435
rect 25179 9404 25513 9432
rect 25179 9401 25191 9404
rect 25133 9395 25191 9401
rect 25501 9401 25513 9404
rect 25547 9432 25559 9435
rect 25860 9435 25918 9441
rect 25860 9432 25872 9435
rect 25547 9404 25872 9432
rect 25547 9401 25559 9404
rect 25501 9395 25559 9401
rect 25860 9401 25872 9404
rect 25906 9432 25918 9435
rect 27522 9432 27528 9444
rect 25906 9404 27528 9432
rect 25906 9401 25918 9404
rect 25860 9395 25918 9401
rect 27522 9392 27528 9404
rect 27580 9392 27586 9444
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 2682 9364 2688 9376
rect 2643 9336 2688 9364
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 5534 9364 5540 9376
rect 5495 9336 5540 9364
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 7558 9364 7564 9376
rect 7519 9336 7564 9364
rect 7558 9324 7564 9336
rect 7616 9324 7622 9376
rect 8018 9324 8024 9376
rect 8076 9364 8082 9376
rect 8113 9367 8171 9373
rect 8113 9364 8125 9367
rect 8076 9336 8125 9364
rect 8076 9324 8082 9336
rect 8113 9333 8125 9336
rect 8159 9333 8171 9367
rect 9674 9364 9680 9376
rect 9635 9336 9680 9364
rect 8113 9327 8171 9333
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 9769 9367 9827 9373
rect 9769 9333 9781 9367
rect 9815 9364 9827 9367
rect 9858 9364 9864 9376
rect 9815 9336 9864 9364
rect 9815 9333 9827 9336
rect 9769 9327 9827 9333
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 10597 9367 10655 9373
rect 10597 9333 10609 9367
rect 10643 9364 10655 9367
rect 10686 9364 10692 9376
rect 10643 9336 10692 9364
rect 10643 9333 10655 9336
rect 10597 9327 10655 9333
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 13081 9367 13139 9373
rect 13081 9333 13093 9367
rect 13127 9364 13139 9367
rect 13998 9364 14004 9376
rect 13127 9336 14004 9364
rect 13127 9333 13139 9336
rect 13081 9327 13139 9333
rect 13998 9324 14004 9336
rect 14056 9364 14062 9376
rect 14458 9364 14464 9376
rect 14056 9336 14464 9364
rect 14056 9324 14062 9336
rect 14458 9324 14464 9336
rect 14516 9364 14522 9376
rect 14553 9367 14611 9373
rect 14553 9364 14565 9367
rect 14516 9336 14565 9364
rect 14516 9324 14522 9336
rect 14553 9333 14565 9336
rect 14599 9333 14611 9367
rect 14553 9327 14611 9333
rect 15562 9324 15568 9376
rect 15620 9364 15626 9376
rect 15657 9367 15715 9373
rect 15657 9364 15669 9367
rect 15620 9336 15669 9364
rect 15620 9324 15626 9336
rect 15657 9333 15669 9336
rect 15703 9333 15715 9367
rect 18230 9364 18236 9376
rect 18191 9336 18236 9364
rect 15657 9327 15715 9333
rect 18230 9324 18236 9336
rect 18288 9324 18294 9376
rect 18693 9367 18751 9373
rect 18693 9333 18705 9367
rect 18739 9364 18751 9367
rect 18782 9364 18788 9376
rect 18739 9336 18788 9364
rect 18739 9333 18751 9336
rect 18693 9327 18751 9333
rect 18782 9324 18788 9336
rect 18840 9324 18846 9376
rect 19150 9324 19156 9376
rect 19208 9364 19214 9376
rect 19245 9367 19303 9373
rect 19245 9364 19257 9367
rect 19208 9336 19257 9364
rect 19208 9324 19214 9336
rect 19245 9333 19257 9336
rect 19291 9333 19303 9367
rect 19245 9327 19303 9333
rect 20806 9324 20812 9376
rect 20864 9364 20870 9376
rect 21085 9367 21143 9373
rect 21085 9364 21097 9367
rect 20864 9336 21097 9364
rect 20864 9324 20870 9336
rect 21085 9333 21097 9336
rect 21131 9364 21143 9367
rect 21266 9364 21272 9376
rect 21131 9336 21272 9364
rect 21131 9333 21143 9336
rect 21085 9327 21143 9333
rect 21266 9324 21272 9336
rect 21324 9324 21330 9376
rect 21450 9364 21456 9376
rect 21411 9336 21456 9364
rect 21450 9324 21456 9336
rect 21508 9324 21514 9376
rect 22002 9364 22008 9376
rect 21963 9336 22008 9364
rect 22002 9324 22008 9336
rect 22060 9324 22066 9376
rect 24118 9364 24124 9376
rect 24079 9336 24124 9364
rect 24118 9324 24124 9336
rect 24176 9324 24182 9376
rect 1104 9274 28888 9296
rect 1104 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 20982 9274
rect 21034 9222 21046 9274
rect 21098 9222 21110 9274
rect 21162 9222 21174 9274
rect 21226 9222 28888 9274
rect 1104 9200 28888 9222
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 4522 9160 4528 9172
rect 4483 9132 4528 9160
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 7469 9163 7527 9169
rect 7469 9129 7481 9163
rect 7515 9160 7527 9163
rect 7650 9160 7656 9172
rect 7515 9132 7656 9160
rect 7515 9129 7527 9132
rect 7469 9123 7527 9129
rect 7650 9120 7656 9132
rect 7708 9120 7714 9172
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 7800 9132 7845 9160
rect 7800 9120 7806 9132
rect 8110 9120 8116 9172
rect 8168 9160 8174 9172
rect 8205 9163 8263 9169
rect 8205 9160 8217 9163
rect 8168 9132 8217 9160
rect 8168 9120 8174 9132
rect 8205 9129 8217 9132
rect 8251 9129 8263 9163
rect 8846 9160 8852 9172
rect 8807 9132 8852 9160
rect 8205 9123 8263 9129
rect 8846 9120 8852 9132
rect 8904 9120 8910 9172
rect 13630 9160 13636 9172
rect 13591 9132 13636 9160
rect 13630 9120 13636 9132
rect 13688 9120 13694 9172
rect 18877 9163 18935 9169
rect 18877 9129 18889 9163
rect 18923 9160 18935 9163
rect 19150 9160 19156 9172
rect 18923 9132 19156 9160
rect 18923 9129 18935 9132
rect 18877 9123 18935 9129
rect 19150 9120 19156 9132
rect 19208 9120 19214 9172
rect 19610 9160 19616 9172
rect 19571 9132 19616 9160
rect 19610 9120 19616 9132
rect 19668 9120 19674 9172
rect 22186 9160 22192 9172
rect 22147 9132 22192 9160
rect 22186 9120 22192 9132
rect 22244 9120 22250 9172
rect 22557 9163 22615 9169
rect 22557 9129 22569 9163
rect 22603 9160 22615 9163
rect 22646 9160 22652 9172
rect 22603 9132 22652 9160
rect 22603 9129 22615 9132
rect 22557 9123 22615 9129
rect 22646 9120 22652 9132
rect 22704 9120 22710 9172
rect 26694 9160 26700 9172
rect 26655 9132 26700 9160
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 1762 9052 1768 9104
rect 1820 9092 1826 9104
rect 2317 9095 2375 9101
rect 2317 9092 2329 9095
rect 1820 9064 2329 9092
rect 1820 9052 1826 9064
rect 2317 9061 2329 9064
rect 2363 9061 2375 9095
rect 8478 9092 8484 9104
rect 2317 9055 2375 9061
rect 7116 9064 8484 9092
rect 7116 9036 7144 9064
rect 8478 9052 8484 9064
rect 8536 9052 8542 9104
rect 13265 9095 13323 9101
rect 13265 9061 13277 9095
rect 13311 9092 13323 9095
rect 13538 9092 13544 9104
rect 13311 9064 13544 9092
rect 13311 9061 13323 9064
rect 13265 9055 13323 9061
rect 13538 9052 13544 9064
rect 13596 9052 13602 9104
rect 19334 9052 19340 9104
rect 19392 9092 19398 9104
rect 20438 9092 20444 9104
rect 19392 9064 20444 9092
rect 19392 9052 19398 9064
rect 20438 9052 20444 9064
rect 20496 9092 20502 9104
rect 25038 9092 25044 9104
rect 20496 9064 25044 9092
rect 20496 9052 20502 9064
rect 25038 9052 25044 9064
rect 25096 9052 25102 9104
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2038 9024 2044 9036
rect 1443 8996 2044 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 7098 9024 7104 9036
rect 7011 8996 7104 9024
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 8018 8984 8024 9036
rect 8076 9024 8082 9036
rect 8113 9027 8171 9033
rect 8113 9024 8125 9027
rect 8076 8996 8125 9024
rect 8076 8984 8082 8996
rect 8113 8993 8125 8996
rect 8159 9024 8171 9027
rect 8570 9024 8576 9036
rect 8159 8996 8576 9024
rect 8159 8993 8171 8996
rect 8113 8987 8171 8993
rect 8570 8984 8576 8996
rect 8628 8984 8634 9036
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 10502 9024 10508 9036
rect 9640 8996 10508 9024
rect 9640 8984 9646 8996
rect 10502 8984 10508 8996
rect 10560 9024 10566 9036
rect 10597 9027 10655 9033
rect 10597 9024 10609 9027
rect 10560 8996 10609 9024
rect 10560 8984 10566 8996
rect 10597 8993 10609 8996
rect 10643 8993 10655 9027
rect 10597 8987 10655 8993
rect 16850 8984 16856 9036
rect 16908 9024 16914 9036
rect 17017 9027 17075 9033
rect 17017 9024 17029 9027
rect 16908 8996 17029 9024
rect 16908 8984 16914 8996
rect 17017 8993 17029 8996
rect 17063 8993 17075 9027
rect 17017 8987 17075 8993
rect 20346 8984 20352 9036
rect 20404 9024 20410 9036
rect 21818 9024 21824 9036
rect 20404 8996 21824 9024
rect 20404 8984 20410 8996
rect 21818 8984 21824 8996
rect 21876 8984 21882 9036
rect 23290 8984 23296 9036
rect 23348 9024 23354 9036
rect 23569 9027 23627 9033
rect 23569 9024 23581 9027
rect 23348 8996 23581 9024
rect 23348 8984 23354 8996
rect 23569 8993 23581 8996
rect 23615 8993 23627 9027
rect 23569 8987 23627 8993
rect 26418 8984 26424 9036
rect 26476 9024 26482 9036
rect 26513 9027 26571 9033
rect 26513 9024 26525 9027
rect 26476 8996 26525 9024
rect 26476 8984 26482 8996
rect 26513 8993 26525 8996
rect 26559 8993 26571 9027
rect 26513 8987 26571 8993
rect 8386 8956 8392 8968
rect 8347 8928 8392 8956
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 16758 8956 16764 8968
rect 16719 8928 16764 8956
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 23658 8956 23664 8968
rect 23619 8928 23664 8956
rect 23658 8916 23664 8928
rect 23716 8916 23722 8968
rect 23845 8959 23903 8965
rect 23845 8925 23857 8959
rect 23891 8956 23903 8959
rect 24210 8956 24216 8968
rect 23891 8928 24216 8956
rect 23891 8925 23903 8928
rect 23845 8919 23903 8925
rect 24210 8916 24216 8928
rect 24268 8916 24274 8968
rect 2406 8848 2412 8900
rect 2464 8888 2470 8900
rect 2590 8888 2596 8900
rect 2464 8860 2596 8888
rect 2464 8848 2470 8860
rect 2590 8848 2596 8860
rect 2648 8888 2654 8900
rect 9309 8891 9367 8897
rect 9309 8888 9321 8891
rect 2648 8860 9321 8888
rect 2648 8848 2654 8860
rect 9309 8857 9321 8860
rect 9355 8888 9367 8891
rect 9674 8888 9680 8900
rect 9355 8860 9680 8888
rect 9355 8857 9367 8860
rect 9309 8851 9367 8857
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 1394 8780 1400 8832
rect 1452 8820 1458 8832
rect 1581 8823 1639 8829
rect 1581 8820 1593 8823
rect 1452 8792 1593 8820
rect 1452 8780 1458 8792
rect 1581 8789 1593 8792
rect 1627 8789 1639 8823
rect 1581 8783 1639 8789
rect 5350 8780 5356 8832
rect 5408 8820 5414 8832
rect 6917 8823 6975 8829
rect 6917 8820 6929 8823
rect 5408 8792 6929 8820
rect 5408 8780 5414 8792
rect 6917 8789 6929 8792
rect 6963 8789 6975 8823
rect 10410 8820 10416 8832
rect 10371 8792 10416 8820
rect 6917 8783 6975 8789
rect 10410 8780 10416 8792
rect 10468 8780 10474 8832
rect 14642 8820 14648 8832
rect 14603 8792 14648 8820
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 18138 8820 18144 8832
rect 18099 8792 18144 8820
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 19242 8820 19248 8832
rect 19203 8792 19248 8820
rect 19242 8780 19248 8792
rect 19300 8780 19306 8832
rect 20162 8780 20168 8832
rect 20220 8820 20226 8832
rect 21266 8820 21272 8832
rect 20220 8792 21272 8820
rect 20220 8780 20226 8792
rect 21266 8780 21272 8792
rect 21324 8820 21330 8832
rect 21637 8823 21695 8829
rect 21637 8820 21649 8823
rect 21324 8792 21649 8820
rect 21324 8780 21330 8792
rect 21637 8789 21649 8792
rect 21683 8789 21695 8823
rect 21637 8783 21695 8789
rect 21910 8780 21916 8832
rect 21968 8820 21974 8832
rect 22278 8820 22284 8832
rect 21968 8792 22284 8820
rect 21968 8780 21974 8792
rect 22278 8780 22284 8792
rect 22336 8780 22342 8832
rect 23198 8820 23204 8832
rect 23159 8792 23204 8820
rect 23198 8780 23204 8792
rect 23256 8780 23262 8832
rect 24210 8820 24216 8832
rect 24171 8792 24216 8820
rect 24210 8780 24216 8792
rect 24268 8780 24274 8832
rect 25682 8820 25688 8832
rect 25643 8792 25688 8820
rect 25682 8780 25688 8792
rect 25740 8780 25746 8832
rect 1104 8730 28888 8752
rect 1104 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 15982 8730
rect 16034 8678 16046 8730
rect 16098 8678 16110 8730
rect 16162 8678 16174 8730
rect 16226 8678 25982 8730
rect 26034 8678 26046 8730
rect 26098 8678 26110 8730
rect 26162 8678 26174 8730
rect 26226 8678 28888 8730
rect 1104 8656 28888 8678
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 4246 8616 4252 8628
rect 4207 8588 4252 8616
rect 4246 8576 4252 8588
rect 4304 8576 4310 8628
rect 7098 8616 7104 8628
rect 7059 8588 7104 8616
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 7837 8619 7895 8625
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 8110 8616 8116 8628
rect 7883 8588 8116 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 8386 8576 8392 8628
rect 8444 8616 8450 8628
rect 8573 8619 8631 8625
rect 8573 8616 8585 8619
rect 8444 8588 8585 8616
rect 8444 8576 8450 8588
rect 8573 8585 8585 8588
rect 8619 8616 8631 8619
rect 10686 8616 10692 8628
rect 8619 8588 10692 8616
rect 8619 8585 8631 8588
rect 8573 8579 8631 8585
rect 10686 8576 10692 8588
rect 10744 8616 10750 8628
rect 11149 8619 11207 8625
rect 11149 8616 11161 8619
rect 10744 8588 11161 8616
rect 10744 8576 10750 8588
rect 11149 8585 11161 8588
rect 11195 8585 11207 8619
rect 14458 8616 14464 8628
rect 14419 8588 14464 8616
rect 11149 8579 11207 8585
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 16025 8619 16083 8625
rect 16025 8585 16037 8619
rect 16071 8616 16083 8619
rect 16850 8616 16856 8628
rect 16071 8588 16856 8616
rect 16071 8585 16083 8588
rect 16025 8579 16083 8585
rect 16850 8576 16856 8588
rect 16908 8576 16914 8628
rect 19337 8619 19395 8625
rect 19337 8585 19349 8619
rect 19383 8616 19395 8619
rect 20346 8616 20352 8628
rect 19383 8588 20352 8616
rect 19383 8585 19395 8588
rect 19337 8579 19395 8585
rect 1578 8548 1584 8560
rect 1539 8520 1584 8548
rect 1578 8508 1584 8520
rect 1636 8508 1642 8560
rect 2406 8480 2412 8492
rect 1412 8452 2412 8480
rect 1412 8421 1440 8452
rect 2406 8440 2412 8452
rect 2464 8440 2470 8492
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8480 4031 8483
rect 5077 8483 5135 8489
rect 5077 8480 5089 8483
rect 4019 8452 5089 8480
rect 4019 8449 4031 8452
rect 3973 8443 4031 8449
rect 5077 8449 5089 8452
rect 5123 8480 5135 8483
rect 5534 8480 5540 8492
rect 5123 8452 5540 8480
rect 5123 8449 5135 8452
rect 5077 8443 5135 8449
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 14476 8480 14504 8576
rect 16758 8508 16764 8560
rect 16816 8548 16822 8560
rect 17129 8551 17187 8557
rect 17129 8548 17141 8551
rect 16816 8520 17141 8548
rect 16816 8508 16822 8520
rect 17129 8517 17141 8520
rect 17175 8548 17187 8551
rect 18785 8551 18843 8557
rect 18785 8548 18797 8551
rect 17175 8520 18797 8548
rect 17175 8517 17187 8520
rect 17129 8511 17187 8517
rect 18785 8517 18797 8520
rect 18831 8548 18843 8551
rect 19242 8548 19248 8560
rect 18831 8520 19248 8548
rect 18831 8517 18843 8520
rect 18785 8511 18843 8517
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 14476 8452 14780 8480
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8381 1455 8415
rect 1397 8375 1455 8381
rect 4246 8372 4252 8424
rect 4304 8412 4310 8424
rect 4893 8415 4951 8421
rect 4893 8412 4905 8415
rect 4304 8384 4905 8412
rect 4304 8372 4310 8384
rect 4893 8381 4905 8384
rect 4939 8381 4951 8415
rect 9769 8415 9827 8421
rect 9769 8412 9781 8415
rect 4893 8375 4951 8381
rect 9324 8384 9781 8412
rect 4522 8304 4528 8356
rect 4580 8344 4586 8356
rect 4801 8347 4859 8353
rect 4801 8344 4813 8347
rect 4580 8316 4813 8344
rect 4580 8304 4586 8316
rect 4801 8313 4813 8316
rect 4847 8313 4859 8347
rect 4801 8307 4859 8313
rect 9324 8288 9352 8384
rect 9769 8381 9781 8384
rect 9815 8412 9827 8415
rect 10410 8412 10416 8424
rect 9815 8384 10416 8412
rect 9815 8381 9827 8384
rect 9769 8375 9827 8381
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 14642 8412 14648 8424
rect 14603 8384 14648 8412
rect 14642 8372 14648 8384
rect 14700 8372 14706 8424
rect 14752 8412 14780 8452
rect 14901 8415 14959 8421
rect 14901 8412 14913 8415
rect 14752 8384 14913 8412
rect 14901 8381 14913 8384
rect 14947 8381 14959 8415
rect 14901 8375 14959 8381
rect 18969 8415 19027 8421
rect 18969 8381 18981 8415
rect 19015 8412 19027 8415
rect 19352 8412 19380 8579
rect 20346 8576 20352 8588
rect 20404 8576 20410 8628
rect 21450 8616 21456 8628
rect 21411 8588 21456 8616
rect 21450 8576 21456 8588
rect 21508 8576 21514 8628
rect 21818 8576 21824 8628
rect 21876 8616 21882 8628
rect 22005 8619 22063 8625
rect 22005 8616 22017 8619
rect 21876 8588 22017 8616
rect 21876 8576 21882 8588
rect 22005 8585 22017 8588
rect 22051 8585 22063 8619
rect 22005 8579 22063 8585
rect 21910 8508 21916 8560
rect 21968 8548 21974 8560
rect 23201 8551 23259 8557
rect 23201 8548 23213 8551
rect 21968 8520 23213 8548
rect 21968 8508 21974 8520
rect 23201 8517 23213 8520
rect 23247 8548 23259 8551
rect 23290 8548 23296 8560
rect 23247 8520 23296 8548
rect 23247 8517 23259 8520
rect 23201 8511 23259 8517
rect 23290 8508 23296 8520
rect 23348 8508 23354 8560
rect 23382 8508 23388 8560
rect 23440 8548 23446 8560
rect 23661 8551 23719 8557
rect 23661 8548 23673 8551
rect 23440 8520 23673 8548
rect 23440 8508 23446 8520
rect 23661 8517 23673 8520
rect 23707 8517 23719 8551
rect 23661 8511 23719 8517
rect 22925 8483 22983 8489
rect 22925 8449 22937 8483
rect 22971 8480 22983 8483
rect 24210 8480 24216 8492
rect 22971 8452 24216 8480
rect 22971 8449 22983 8452
rect 22925 8443 22983 8449
rect 24210 8440 24216 8452
rect 24268 8440 24274 8492
rect 19015 8384 19380 8412
rect 20073 8415 20131 8421
rect 19015 8381 19027 8384
rect 18969 8375 19027 8381
rect 20073 8381 20085 8415
rect 20119 8412 20131 8415
rect 20162 8412 20168 8424
rect 20119 8384 20168 8412
rect 20119 8381 20131 8384
rect 20073 8375 20131 8381
rect 20162 8372 20168 8384
rect 20220 8372 20226 8424
rect 9677 8347 9735 8353
rect 9677 8313 9689 8347
rect 9723 8344 9735 8347
rect 10014 8347 10072 8353
rect 10014 8344 10026 8347
rect 9723 8316 10026 8344
rect 9723 8313 9735 8316
rect 9677 8307 9735 8313
rect 10014 8313 10026 8316
rect 10060 8344 10072 8347
rect 10134 8344 10140 8356
rect 10060 8316 10140 8344
rect 10060 8313 10072 8316
rect 10014 8307 10072 8313
rect 10134 8304 10140 8316
rect 10192 8304 10198 8356
rect 19981 8347 20039 8353
rect 19981 8313 19993 8347
rect 20027 8344 20039 8347
rect 20318 8347 20376 8353
rect 20318 8344 20330 8347
rect 20027 8316 20330 8344
rect 20027 8313 20039 8316
rect 19981 8307 20039 8313
rect 20318 8313 20330 8316
rect 20364 8344 20376 8347
rect 20806 8344 20812 8356
rect 20364 8316 20812 8344
rect 20364 8313 20376 8316
rect 20318 8307 20376 8313
rect 20806 8304 20812 8316
rect 20864 8304 20870 8356
rect 24029 8347 24087 8353
rect 24029 8313 24041 8347
rect 24075 8344 24087 8347
rect 24486 8344 24492 8356
rect 24075 8316 24492 8344
rect 24075 8313 24087 8316
rect 24029 8307 24087 8313
rect 24486 8304 24492 8316
rect 24544 8344 24550 8356
rect 25041 8347 25099 8353
rect 25041 8344 25053 8347
rect 24544 8316 25053 8344
rect 24544 8304 24550 8316
rect 25041 8313 25053 8316
rect 25087 8313 25099 8347
rect 25041 8307 25099 8313
rect 26418 8304 26424 8356
rect 26476 8344 26482 8356
rect 26513 8347 26571 8353
rect 26513 8344 26525 8347
rect 26476 8316 26525 8344
rect 26476 8304 26482 8316
rect 26513 8313 26525 8316
rect 26559 8313 26571 8347
rect 26513 8307 26571 8313
rect 4430 8276 4436 8288
rect 4391 8248 4436 8276
rect 4430 8236 4436 8248
rect 4488 8236 4494 8288
rect 8018 8236 8024 8288
rect 8076 8276 8082 8288
rect 8113 8279 8171 8285
rect 8113 8276 8125 8279
rect 8076 8248 8125 8276
rect 8076 8236 8082 8248
rect 8113 8245 8125 8248
rect 8159 8245 8171 8279
rect 9306 8276 9312 8288
rect 9267 8248 9312 8276
rect 8113 8239 8171 8245
rect 9306 8236 9312 8248
rect 9364 8236 9370 8288
rect 24121 8279 24179 8285
rect 24121 8245 24133 8279
rect 24167 8276 24179 8279
rect 24394 8276 24400 8288
rect 24167 8248 24400 8276
rect 24167 8245 24179 8248
rect 24121 8239 24179 8245
rect 24394 8236 24400 8248
rect 24452 8276 24458 8288
rect 24673 8279 24731 8285
rect 24673 8276 24685 8279
rect 24452 8248 24685 8276
rect 24452 8236 24458 8248
rect 24673 8245 24685 8248
rect 24719 8245 24731 8279
rect 24673 8239 24731 8245
rect 1104 8186 28888 8208
rect 1104 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 20982 8186
rect 21034 8134 21046 8186
rect 21098 8134 21110 8186
rect 21162 8134 21174 8186
rect 21226 8134 28888 8186
rect 1104 8112 28888 8134
rect 1486 8032 1492 8084
rect 1544 8072 1550 8084
rect 1581 8075 1639 8081
rect 1581 8072 1593 8075
rect 1544 8044 1593 8072
rect 1544 8032 1550 8044
rect 1581 8041 1593 8044
rect 1627 8041 1639 8075
rect 1581 8035 1639 8041
rect 4430 8032 4436 8084
rect 4488 8072 4494 8084
rect 4525 8075 4583 8081
rect 4525 8072 4537 8075
rect 4488 8044 4537 8072
rect 4488 8032 4494 8044
rect 4525 8041 4537 8044
rect 4571 8041 4583 8075
rect 10502 8072 10508 8084
rect 10463 8044 10508 8072
rect 4525 8035 4583 8041
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 21542 8072 21548 8084
rect 21455 8044 21548 8072
rect 21542 8032 21548 8044
rect 21600 8072 21606 8084
rect 22002 8072 22008 8084
rect 21600 8044 22008 8072
rect 21600 8032 21606 8044
rect 22002 8032 22008 8044
rect 22060 8032 22066 8084
rect 23293 8075 23351 8081
rect 23293 8041 23305 8075
rect 23339 8072 23351 8075
rect 23658 8072 23664 8084
rect 23339 8044 23664 8072
rect 23339 8041 23351 8044
rect 23293 8035 23351 8041
rect 23658 8032 23664 8044
rect 23716 8072 23722 8084
rect 24029 8075 24087 8081
rect 24029 8072 24041 8075
rect 23716 8044 24041 8072
rect 23716 8032 23722 8044
rect 24029 8041 24041 8044
rect 24075 8041 24087 8075
rect 24029 8035 24087 8041
rect 24118 8032 24124 8084
rect 24176 8072 24182 8084
rect 24397 8075 24455 8081
rect 24397 8072 24409 8075
rect 24176 8044 24409 8072
rect 24176 8032 24182 8044
rect 24397 8041 24409 8044
rect 24443 8072 24455 8075
rect 24762 8072 24768 8084
rect 24443 8044 24768 8072
rect 24443 8041 24455 8044
rect 24397 8035 24455 8041
rect 24762 8032 24768 8044
rect 24820 8032 24826 8084
rect 26694 8072 26700 8084
rect 26655 8044 26700 8072
rect 26694 8032 26700 8044
rect 26752 8032 26758 8084
rect 5534 7964 5540 8016
rect 5592 8004 5598 8016
rect 5718 8004 5724 8016
rect 5592 7976 5724 8004
rect 5592 7964 5598 7976
rect 5718 7964 5724 7976
rect 5776 8004 5782 8016
rect 5966 8007 6024 8013
rect 5966 8004 5978 8007
rect 5776 7976 5978 8004
rect 5776 7964 5782 7976
rect 5966 7973 5978 7976
rect 6012 7973 6024 8007
rect 5966 7967 6024 7973
rect 23753 8007 23811 8013
rect 23753 7973 23765 8007
rect 23799 8004 23811 8007
rect 24210 8004 24216 8016
rect 23799 7976 24216 8004
rect 23799 7973 23811 7976
rect 23753 7967 23811 7973
rect 24210 7964 24216 7976
rect 24268 7964 24274 8016
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1946 7936 1952 7948
rect 1443 7908 1952 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1946 7896 1952 7908
rect 2004 7896 2010 7948
rect 4338 7896 4344 7948
rect 4396 7936 4402 7948
rect 4433 7939 4491 7945
rect 4433 7936 4445 7939
rect 4396 7908 4445 7936
rect 4396 7896 4402 7908
rect 4433 7905 4445 7908
rect 4479 7905 4491 7939
rect 4433 7899 4491 7905
rect 11514 7896 11520 7948
rect 11572 7936 11578 7948
rect 11681 7939 11739 7945
rect 11681 7936 11693 7939
rect 11572 7908 11693 7936
rect 11572 7896 11578 7908
rect 11681 7905 11693 7908
rect 11727 7905 11739 7939
rect 11681 7899 11739 7905
rect 15562 7896 15568 7948
rect 15620 7936 15626 7948
rect 16301 7939 16359 7945
rect 16301 7936 16313 7939
rect 15620 7908 16313 7936
rect 15620 7896 15626 7908
rect 16301 7905 16313 7908
rect 16347 7905 16359 7939
rect 21634 7936 21640 7948
rect 21595 7908 21640 7936
rect 16301 7899 16359 7905
rect 21634 7896 21640 7908
rect 21692 7896 21698 7948
rect 25866 7896 25872 7948
rect 25924 7936 25930 7948
rect 26513 7939 26571 7945
rect 26513 7936 26525 7939
rect 25924 7908 26525 7936
rect 25924 7896 25930 7908
rect 26513 7905 26525 7908
rect 26559 7905 26571 7939
rect 26513 7899 26571 7905
rect 4614 7868 4620 7880
rect 4575 7840 4620 7868
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 5350 7828 5356 7880
rect 5408 7868 5414 7880
rect 5721 7871 5779 7877
rect 5721 7868 5733 7871
rect 5408 7840 5733 7868
rect 5408 7828 5414 7840
rect 5721 7837 5733 7840
rect 5767 7837 5779 7871
rect 11422 7868 11428 7880
rect 11383 7840 11428 7868
rect 5721 7831 5779 7837
rect 11422 7828 11428 7840
rect 11480 7828 11486 7880
rect 16390 7868 16396 7880
rect 16351 7840 16396 7868
rect 16390 7828 16396 7840
rect 16448 7828 16454 7880
rect 16574 7868 16580 7880
rect 16535 7840 16580 7868
rect 16574 7828 16580 7840
rect 16632 7828 16638 7880
rect 21726 7868 21732 7880
rect 21687 7840 21732 7868
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 23934 7828 23940 7880
rect 23992 7868 23998 7880
rect 24489 7871 24547 7877
rect 24489 7868 24501 7871
rect 23992 7840 24501 7868
rect 23992 7828 23998 7840
rect 24489 7837 24501 7840
rect 24535 7837 24547 7871
rect 24489 7831 24547 7837
rect 24673 7871 24731 7877
rect 24673 7837 24685 7871
rect 24719 7868 24731 7871
rect 24719 7840 25084 7868
rect 24719 7837 24731 7840
rect 24673 7831 24731 7837
rect 25056 7744 25084 7840
rect 1762 7692 1768 7744
rect 1820 7732 1826 7744
rect 1949 7735 2007 7741
rect 1949 7732 1961 7735
rect 1820 7704 1961 7732
rect 1820 7692 1826 7704
rect 1949 7701 1961 7704
rect 1995 7701 2007 7735
rect 4062 7732 4068 7744
rect 4023 7704 4068 7732
rect 1949 7695 2007 7701
rect 4062 7692 4068 7704
rect 4120 7692 4126 7744
rect 6362 7692 6368 7744
rect 6420 7732 6426 7744
rect 7101 7735 7159 7741
rect 7101 7732 7113 7735
rect 6420 7704 7113 7732
rect 6420 7692 6426 7704
rect 7101 7701 7113 7704
rect 7147 7732 7159 7735
rect 7374 7732 7380 7744
rect 7147 7704 7380 7732
rect 7147 7701 7159 7704
rect 7101 7695 7159 7701
rect 7374 7692 7380 7704
rect 7432 7692 7438 7744
rect 12802 7732 12808 7744
rect 12763 7704 12808 7732
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 14553 7735 14611 7741
rect 14553 7701 14565 7735
rect 14599 7732 14611 7735
rect 14642 7732 14648 7744
rect 14599 7704 14648 7732
rect 14599 7701 14611 7704
rect 14553 7695 14611 7701
rect 14642 7692 14648 7704
rect 14700 7692 14706 7744
rect 15933 7735 15991 7741
rect 15933 7701 15945 7735
rect 15979 7732 15991 7735
rect 16298 7732 16304 7744
rect 15979 7704 16304 7732
rect 15979 7701 15991 7704
rect 15933 7695 15991 7701
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 20162 7732 20168 7744
rect 20123 7704 20168 7732
rect 20162 7692 20168 7704
rect 20220 7692 20226 7744
rect 20714 7692 20720 7744
rect 20772 7732 20778 7744
rect 21177 7735 21235 7741
rect 21177 7732 21189 7735
rect 20772 7704 21189 7732
rect 20772 7692 20778 7704
rect 21177 7701 21189 7704
rect 21223 7701 21235 7735
rect 25038 7732 25044 7744
rect 24999 7704 25044 7732
rect 21177 7695 21235 7701
rect 25038 7692 25044 7704
rect 25096 7692 25102 7744
rect 25682 7692 25688 7744
rect 25740 7732 25746 7744
rect 26145 7735 26203 7741
rect 26145 7732 26157 7735
rect 25740 7704 26157 7732
rect 25740 7692 25746 7704
rect 26145 7701 26157 7704
rect 26191 7701 26203 7735
rect 26145 7695 26203 7701
rect 26786 7692 26792 7744
rect 26844 7732 26850 7744
rect 27062 7732 27068 7744
rect 26844 7704 27068 7732
rect 26844 7692 26850 7704
rect 27062 7692 27068 7704
rect 27120 7692 27126 7744
rect 1104 7642 28888 7664
rect 1104 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 15982 7642
rect 16034 7590 16046 7642
rect 16098 7590 16110 7642
rect 16162 7590 16174 7642
rect 16226 7590 25982 7642
rect 26034 7590 26046 7642
rect 26098 7590 26110 7642
rect 26162 7590 26174 7642
rect 26226 7590 28888 7642
rect 1104 7568 28888 7590
rect 4157 7531 4215 7537
rect 4157 7497 4169 7531
rect 4203 7528 4215 7531
rect 4338 7528 4344 7540
rect 4203 7500 4344 7528
rect 4203 7497 4215 7500
rect 4157 7491 4215 7497
rect 4338 7488 4344 7500
rect 4396 7488 4402 7540
rect 4430 7488 4436 7540
rect 4488 7528 4494 7540
rect 4801 7531 4859 7537
rect 4801 7528 4813 7531
rect 4488 7500 4813 7528
rect 4488 7488 4494 7500
rect 4801 7497 4813 7500
rect 4847 7497 4859 7531
rect 5718 7528 5724 7540
rect 5679 7500 5724 7528
rect 4801 7491 4859 7497
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 10134 7528 10140 7540
rect 10095 7500 10140 7528
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 11514 7528 11520 7540
rect 11475 7500 11520 7528
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 12434 7528 12440 7540
rect 11808 7500 12440 7528
rect 5534 7420 5540 7472
rect 5592 7460 5598 7472
rect 6825 7463 6883 7469
rect 6825 7460 6837 7463
rect 5592 7432 6837 7460
rect 5592 7420 5598 7432
rect 6825 7429 6837 7432
rect 6871 7429 6883 7463
rect 6825 7423 6883 7429
rect 7374 7392 7380 7404
rect 7335 7364 7380 7392
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 1489 7327 1547 7333
rect 1489 7293 1501 7327
rect 1535 7324 1547 7327
rect 2682 7324 2688 7336
rect 1535 7296 2688 7324
rect 1535 7293 1547 7296
rect 1489 7287 1547 7293
rect 2682 7284 2688 7296
rect 2740 7324 2746 7336
rect 5350 7324 5356 7336
rect 2740 7296 5356 7324
rect 2740 7284 2746 7296
rect 5350 7284 5356 7296
rect 5408 7284 5414 7336
rect 6638 7324 6644 7336
rect 6551 7296 6644 7324
rect 6638 7284 6644 7296
rect 6696 7324 6702 7336
rect 7282 7324 7288 7336
rect 6696 7296 7288 7324
rect 6696 7284 6702 7296
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 8754 7324 8760 7336
rect 8715 7296 8760 7324
rect 8754 7284 8760 7296
rect 8812 7324 8818 7336
rect 9306 7324 9312 7336
rect 8812 7296 9312 7324
rect 8812 7284 8818 7296
rect 9306 7284 9312 7296
rect 9364 7324 9370 7336
rect 11422 7324 11428 7336
rect 9364 7296 11428 7324
rect 9364 7284 9370 7296
rect 11422 7284 11428 7296
rect 11480 7324 11486 7336
rect 11808 7333 11836 7500
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 20806 7488 20812 7540
rect 20864 7528 20870 7540
rect 21269 7531 21327 7537
rect 21269 7528 21281 7531
rect 20864 7500 21281 7528
rect 20864 7488 20870 7500
rect 21269 7497 21281 7500
rect 21315 7528 21327 7531
rect 21726 7528 21732 7540
rect 21315 7500 21732 7528
rect 21315 7497 21327 7500
rect 21269 7491 21327 7497
rect 21726 7488 21732 7500
rect 21784 7528 21790 7540
rect 21821 7531 21879 7537
rect 21821 7528 21833 7531
rect 21784 7500 21833 7528
rect 21784 7488 21790 7500
rect 21821 7497 21833 7500
rect 21867 7497 21879 7531
rect 24394 7528 24400 7540
rect 24355 7500 24400 7528
rect 21821 7491 21879 7497
rect 24394 7488 24400 7500
rect 24452 7488 24458 7540
rect 25501 7531 25559 7537
rect 25501 7497 25513 7531
rect 25547 7528 25559 7531
rect 25590 7528 25596 7540
rect 25547 7500 25596 7528
rect 25547 7497 25559 7500
rect 25501 7491 25559 7497
rect 25590 7488 25596 7500
rect 25648 7488 25654 7540
rect 27522 7528 27528 7540
rect 27483 7500 27528 7528
rect 27522 7488 27528 7500
rect 27580 7488 27586 7540
rect 13078 7420 13084 7472
rect 13136 7460 13142 7472
rect 14461 7463 14519 7469
rect 14461 7460 14473 7463
rect 13136 7432 14473 7460
rect 13136 7420 13142 7432
rect 14461 7429 14473 7432
rect 14507 7429 14519 7463
rect 14461 7423 14519 7429
rect 16117 7463 16175 7469
rect 16117 7429 16129 7463
rect 16163 7460 16175 7463
rect 16390 7460 16396 7472
rect 16163 7432 16396 7460
rect 16163 7429 16175 7432
rect 16117 7423 16175 7429
rect 16390 7420 16396 7432
rect 16448 7460 16454 7472
rect 17497 7463 17555 7469
rect 17497 7460 17509 7463
rect 16448 7432 17509 7460
rect 16448 7420 16454 7432
rect 17497 7429 17509 7432
rect 17543 7429 17555 7463
rect 24210 7460 24216 7472
rect 24171 7432 24216 7460
rect 17497 7423 17555 7429
rect 24210 7420 24216 7432
rect 24268 7420 24274 7472
rect 13262 7352 13268 7404
rect 13320 7392 13326 7404
rect 13541 7395 13599 7401
rect 13541 7392 13553 7395
rect 13320 7364 13553 7392
rect 13320 7352 13326 7364
rect 13541 7361 13553 7364
rect 13587 7392 13599 7395
rect 14642 7392 14648 7404
rect 13587 7364 14648 7392
rect 13587 7361 13599 7364
rect 13541 7355 13599 7361
rect 14642 7352 14648 7364
rect 14700 7392 14706 7404
rect 15013 7395 15071 7401
rect 15013 7392 15025 7395
rect 14700 7364 15025 7392
rect 14700 7352 14706 7364
rect 15013 7361 15025 7364
rect 15059 7361 15071 7395
rect 15013 7355 15071 7361
rect 16761 7395 16819 7401
rect 16761 7361 16773 7395
rect 16807 7392 16819 7395
rect 16850 7392 16856 7404
rect 16807 7364 16856 7392
rect 16807 7361 16819 7364
rect 16761 7355 16819 7361
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 19797 7395 19855 7401
rect 19797 7361 19809 7395
rect 19843 7392 19855 7395
rect 23477 7395 23535 7401
rect 19843 7364 20024 7392
rect 19843 7361 19855 7364
rect 19797 7355 19855 7361
rect 11793 7327 11851 7333
rect 11793 7324 11805 7327
rect 11480 7296 11805 7324
rect 11480 7284 11486 7296
rect 11793 7293 11805 7296
rect 11839 7293 11851 7327
rect 15746 7324 15752 7336
rect 11793 7287 11851 7293
rect 14200 7296 15752 7324
rect 1762 7265 1768 7268
rect 1756 7256 1768 7265
rect 1723 7228 1768 7256
rect 1756 7219 1768 7228
rect 1820 7256 1826 7268
rect 4433 7259 4491 7265
rect 4433 7256 4445 7259
rect 1820 7228 4445 7256
rect 1762 7216 1768 7219
rect 1820 7216 1826 7228
rect 4433 7225 4445 7228
rect 4479 7256 4491 7259
rect 4614 7256 4620 7268
rect 4479 7228 4620 7256
rect 4479 7225 4491 7228
rect 4433 7219 4491 7225
rect 4614 7216 4620 7228
rect 4672 7256 4678 7268
rect 6181 7259 6239 7265
rect 6181 7256 6193 7259
rect 4672 7228 6193 7256
rect 4672 7216 4678 7228
rect 6181 7225 6193 7228
rect 6227 7256 6239 7259
rect 6362 7256 6368 7268
rect 6227 7228 6368 7256
rect 6227 7225 6239 7228
rect 6181 7219 6239 7225
rect 6362 7216 6368 7228
rect 6420 7216 6426 7268
rect 8665 7259 8723 7265
rect 8665 7225 8677 7259
rect 8711 7256 8723 7259
rect 9002 7259 9060 7265
rect 9002 7256 9014 7259
rect 8711 7228 9014 7256
rect 8711 7225 8723 7228
rect 8665 7219 8723 7225
rect 9002 7225 9014 7228
rect 9048 7256 9060 7259
rect 9582 7256 9588 7268
rect 9048 7228 9588 7256
rect 9048 7225 9060 7228
rect 9002 7219 9060 7225
rect 9582 7216 9588 7228
rect 9640 7216 9646 7268
rect 12805 7259 12863 7265
rect 12805 7225 12817 7259
rect 12851 7256 12863 7259
rect 13265 7259 13323 7265
rect 13265 7256 13277 7259
rect 12851 7228 13277 7256
rect 12851 7225 12863 7228
rect 12805 7219 12863 7225
rect 13265 7225 13277 7228
rect 13311 7256 13323 7259
rect 13446 7256 13452 7268
rect 13311 7228 13452 7256
rect 13311 7225 13323 7228
rect 13265 7219 13323 7225
rect 13446 7216 13452 7228
rect 13504 7216 13510 7268
rect 2866 7188 2872 7200
rect 2827 7160 2872 7188
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 7190 7188 7196 7200
rect 7151 7160 7196 7188
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 12158 7188 12164 7200
rect 12119 7160 12164 7188
rect 12158 7148 12164 7160
rect 12216 7148 12222 7200
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13354 7188 13360 7200
rect 13315 7160 13360 7188
rect 13354 7148 13360 7160
rect 13412 7188 13418 7200
rect 14200 7188 14228 7296
rect 15746 7284 15752 7296
rect 15804 7284 15810 7336
rect 16574 7284 16580 7336
rect 16632 7324 16638 7336
rect 17221 7327 17279 7333
rect 17221 7324 17233 7327
rect 16632 7296 17233 7324
rect 16632 7284 16638 7296
rect 17221 7293 17233 7296
rect 17267 7324 17279 7327
rect 18138 7324 18144 7336
rect 17267 7296 18144 7324
rect 17267 7293 17279 7296
rect 17221 7287 17279 7293
rect 18138 7284 18144 7296
rect 18196 7284 18202 7336
rect 19334 7284 19340 7336
rect 19392 7324 19398 7336
rect 19886 7324 19892 7336
rect 19392 7296 19892 7324
rect 19392 7284 19398 7296
rect 19886 7284 19892 7296
rect 19944 7284 19950 7336
rect 19996 7324 20024 7364
rect 23477 7361 23489 7395
rect 23523 7392 23535 7395
rect 25038 7392 25044 7404
rect 23523 7364 25044 7392
rect 23523 7361 23535 7364
rect 23477 7355 23535 7361
rect 25038 7352 25044 7364
rect 25096 7352 25102 7404
rect 25682 7352 25688 7404
rect 25740 7392 25746 7404
rect 26145 7395 26203 7401
rect 26145 7392 26157 7395
rect 25740 7364 26157 7392
rect 25740 7352 25746 7364
rect 26145 7361 26157 7364
rect 26191 7361 26203 7395
rect 26145 7355 26203 7361
rect 20156 7327 20214 7333
rect 20156 7324 20168 7327
rect 19996 7296 20168 7324
rect 20156 7293 20168 7296
rect 20202 7324 20214 7327
rect 20622 7324 20628 7336
rect 20202 7296 20628 7324
rect 20202 7293 20214 7296
rect 20156 7287 20214 7293
rect 20622 7284 20628 7296
rect 20680 7284 20686 7336
rect 24210 7284 24216 7336
rect 24268 7324 24274 7336
rect 24857 7327 24915 7333
rect 24857 7324 24869 7327
rect 24268 7296 24869 7324
rect 24268 7284 24274 7296
rect 24857 7293 24869 7296
rect 24903 7293 24915 7327
rect 25958 7324 25964 7336
rect 25919 7296 25964 7324
rect 24857 7287 24915 7293
rect 25958 7284 25964 7296
rect 26016 7284 26022 7336
rect 14366 7256 14372 7268
rect 14279 7228 14372 7256
rect 14366 7216 14372 7228
rect 14424 7256 14430 7268
rect 14424 7228 14964 7256
rect 14424 7216 14430 7228
rect 14936 7200 14964 7228
rect 15378 7216 15384 7268
rect 15436 7256 15442 7268
rect 15933 7259 15991 7265
rect 15933 7256 15945 7259
rect 15436 7228 15945 7256
rect 15436 7216 15442 7228
rect 15933 7225 15945 7228
rect 15979 7256 15991 7259
rect 16666 7256 16672 7268
rect 15979 7228 16672 7256
rect 15979 7225 15991 7228
rect 15933 7219 15991 7225
rect 13412 7160 14228 7188
rect 13412 7148 13418 7160
rect 14550 7148 14556 7200
rect 14608 7188 14614 7200
rect 14829 7191 14887 7197
rect 14829 7188 14841 7191
rect 14608 7160 14841 7188
rect 14608 7148 14614 7160
rect 14829 7157 14841 7160
rect 14875 7157 14887 7191
rect 14829 7151 14887 7157
rect 14918 7148 14924 7200
rect 14976 7188 14982 7200
rect 15562 7188 15568 7200
rect 14976 7160 15021 7188
rect 15523 7160 15568 7188
rect 14976 7148 14982 7160
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 16114 7148 16120 7200
rect 16172 7188 16178 7200
rect 16592 7197 16620 7228
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 24765 7259 24823 7265
rect 24765 7225 24777 7259
rect 24811 7256 24823 7259
rect 25590 7256 25596 7268
rect 24811 7228 25596 7256
rect 24811 7225 24823 7228
rect 24765 7219 24823 7225
rect 25590 7216 25596 7228
rect 25648 7216 25654 7268
rect 26412 7259 26470 7265
rect 26412 7225 26424 7259
rect 26458 7256 26470 7259
rect 26786 7256 26792 7268
rect 26458 7228 26792 7256
rect 26458 7225 26470 7228
rect 26412 7219 26470 7225
rect 26786 7216 26792 7228
rect 26844 7216 26850 7268
rect 16485 7191 16543 7197
rect 16485 7188 16497 7191
rect 16172 7160 16497 7188
rect 16172 7148 16178 7160
rect 16485 7157 16497 7160
rect 16531 7157 16543 7191
rect 16485 7151 16543 7157
rect 16577 7191 16635 7197
rect 16577 7157 16589 7191
rect 16623 7157 16635 7191
rect 16577 7151 16635 7157
rect 18141 7191 18199 7197
rect 18141 7157 18153 7191
rect 18187 7188 18199 7191
rect 18966 7188 18972 7200
rect 18187 7160 18972 7188
rect 18187 7157 18199 7160
rect 18141 7151 18199 7157
rect 18966 7148 18972 7160
rect 19024 7148 19030 7200
rect 23934 7188 23940 7200
rect 23895 7160 23940 7188
rect 23934 7148 23940 7160
rect 23992 7148 23998 7200
rect 1104 7098 28888 7120
rect 1104 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 20982 7098
rect 21034 7046 21046 7098
rect 21098 7046 21110 7098
rect 21162 7046 21174 7098
rect 21226 7046 28888 7098
rect 1104 7024 28888 7046
rect 1946 6984 1952 6996
rect 1907 6956 1952 6984
rect 1946 6944 1952 6956
rect 2004 6944 2010 6996
rect 3329 6987 3387 6993
rect 3329 6953 3341 6987
rect 3375 6984 3387 6987
rect 3694 6984 3700 6996
rect 3375 6956 3700 6984
rect 3375 6953 3387 6956
rect 3329 6947 3387 6953
rect 3694 6944 3700 6956
rect 3752 6984 3758 6996
rect 4062 6984 4068 6996
rect 3752 6956 4068 6984
rect 3752 6944 3758 6956
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 6178 6984 6184 6996
rect 6139 6956 6184 6984
rect 6178 6944 6184 6956
rect 6236 6944 6242 6996
rect 12621 6987 12679 6993
rect 12621 6953 12633 6987
rect 12667 6984 12679 6987
rect 12894 6984 12900 6996
rect 12667 6956 12900 6984
rect 12667 6953 12679 6956
rect 12621 6947 12679 6953
rect 12894 6944 12900 6956
rect 12952 6944 12958 6996
rect 13262 6984 13268 6996
rect 13223 6956 13268 6984
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 13725 6987 13783 6993
rect 13725 6953 13737 6987
rect 13771 6984 13783 6987
rect 14550 6984 14556 6996
rect 13771 6956 14556 6984
rect 13771 6953 13783 6956
rect 13725 6947 13783 6953
rect 14550 6944 14556 6956
rect 14608 6944 14614 6996
rect 18966 6984 18972 6996
rect 18927 6956 18972 6984
rect 18966 6944 18972 6956
rect 19024 6984 19030 6996
rect 19334 6984 19340 6996
rect 19024 6956 19340 6984
rect 19024 6944 19030 6956
rect 19334 6944 19340 6956
rect 19392 6944 19398 6996
rect 19886 6984 19892 6996
rect 19847 6956 19892 6984
rect 19886 6944 19892 6956
rect 19944 6944 19950 6996
rect 21269 6987 21327 6993
rect 21269 6953 21281 6987
rect 21315 6984 21327 6987
rect 21634 6984 21640 6996
rect 21315 6956 21640 6984
rect 21315 6953 21327 6956
rect 21269 6947 21327 6953
rect 21634 6944 21640 6956
rect 21692 6944 21698 6996
rect 22833 6987 22891 6993
rect 22833 6953 22845 6987
rect 22879 6984 22891 6987
rect 23198 6984 23204 6996
rect 22879 6956 23204 6984
rect 22879 6953 22891 6956
rect 22833 6947 22891 6953
rect 23198 6944 23204 6956
rect 23256 6944 23262 6996
rect 24118 6984 24124 6996
rect 24079 6956 24124 6984
rect 24118 6944 24124 6956
rect 24176 6944 24182 6996
rect 24762 6984 24768 6996
rect 24723 6956 24768 6984
rect 24762 6944 24768 6956
rect 24820 6984 24826 6996
rect 24946 6984 24952 6996
rect 24820 6956 24952 6984
rect 24820 6944 24826 6956
rect 24946 6944 24952 6956
rect 25004 6944 25010 6996
rect 3878 6876 3884 6928
rect 3936 6916 3942 6928
rect 10045 6919 10103 6925
rect 3936 6888 4384 6916
rect 3936 6876 3942 6888
rect 4356 6860 4384 6888
rect 10045 6885 10057 6919
rect 10091 6916 10103 6919
rect 10091 6888 11100 6916
rect 10091 6885 10103 6888
rect 10045 6879 10103 6885
rect 11072 6860 11100 6888
rect 11514 6876 11520 6928
rect 11572 6916 11578 6928
rect 13280 6916 13308 6944
rect 21542 6916 21548 6928
rect 11572 6888 13308 6916
rect 21503 6888 21548 6916
rect 11572 6876 11578 6888
rect 21542 6876 21548 6888
rect 21600 6876 21606 6928
rect 23290 6876 23296 6928
rect 23348 6916 23354 6928
rect 23348 6888 26556 6916
rect 23348 6876 23354 6888
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 2130 6848 2136 6860
rect 1443 6820 2136 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 2130 6808 2136 6820
rect 2188 6808 2194 6860
rect 4338 6808 4344 6860
rect 4396 6848 4402 6860
rect 4433 6851 4491 6857
rect 4433 6848 4445 6851
rect 4396 6820 4445 6848
rect 4396 6808 4402 6820
rect 4433 6817 4445 6820
rect 4479 6817 4491 6851
rect 4433 6811 4491 6817
rect 4525 6851 4583 6857
rect 4525 6817 4537 6851
rect 4571 6848 4583 6851
rect 4706 6848 4712 6860
rect 4571 6820 4712 6848
rect 4571 6817 4583 6820
rect 4525 6811 4583 6817
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 6917 6851 6975 6857
rect 6917 6817 6929 6851
rect 6963 6848 6975 6851
rect 7190 6848 7196 6860
rect 6963 6820 7196 6848
rect 6963 6817 6975 6820
rect 6917 6811 6975 6817
rect 7190 6808 7196 6820
rect 7248 6848 7254 6860
rect 7377 6851 7435 6857
rect 7377 6848 7389 6851
rect 7248 6820 7389 6848
rect 7248 6808 7254 6820
rect 7377 6817 7389 6820
rect 7423 6817 7435 6851
rect 7377 6811 7435 6817
rect 11054 6808 11060 6860
rect 11112 6808 11118 6860
rect 12529 6851 12587 6857
rect 12529 6817 12541 6851
rect 12575 6848 12587 6851
rect 13078 6848 13084 6860
rect 12575 6820 13084 6848
rect 12575 6817 12587 6820
rect 12529 6811 12587 6817
rect 13078 6808 13084 6820
rect 13136 6808 13142 6860
rect 16577 6851 16635 6857
rect 16577 6817 16589 6851
rect 16623 6848 16635 6851
rect 16850 6848 16856 6860
rect 16623 6820 16856 6848
rect 16623 6817 16635 6820
rect 16577 6811 16635 6817
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 16945 6851 17003 6857
rect 16945 6817 16957 6851
rect 16991 6848 17003 6851
rect 17405 6851 17463 6857
rect 17405 6848 17417 6851
rect 16991 6820 17417 6848
rect 16991 6817 17003 6820
rect 16945 6811 17003 6817
rect 17405 6817 17417 6820
rect 17451 6848 17463 6851
rect 19058 6848 19064 6860
rect 17451 6820 18644 6848
rect 19019 6820 19064 6848
rect 17451 6817 17463 6820
rect 17405 6811 17463 6817
rect 4614 6780 4620 6792
rect 4575 6752 4620 6780
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 6270 6780 6276 6792
rect 6231 6752 6276 6780
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 6362 6740 6368 6792
rect 6420 6780 6426 6792
rect 10134 6780 10140 6792
rect 6420 6752 6465 6780
rect 10095 6752 10140 6780
rect 6420 6740 6426 6752
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 12802 6780 12808 6792
rect 10284 6752 10329 6780
rect 12763 6752 12808 6780
rect 10284 6740 10290 6752
rect 12802 6740 12808 6752
rect 12860 6740 12866 6792
rect 16114 6780 16120 6792
rect 16075 6752 16120 6780
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 17494 6780 17500 6792
rect 17455 6752 17500 6780
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 17586 6740 17592 6792
rect 17644 6780 17650 6792
rect 18138 6780 18144 6792
rect 17644 6752 17689 6780
rect 18099 6752 18144 6780
rect 17644 6740 17650 6752
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 1578 6712 1584 6724
rect 1539 6684 1584 6712
rect 1578 6672 1584 6684
rect 1636 6672 1642 6724
rect 18616 6721 18644 6820
rect 19058 6808 19064 6820
rect 19116 6808 19122 6860
rect 22922 6848 22928 6860
rect 22835 6820 22928 6848
rect 22922 6808 22928 6820
rect 22980 6848 22986 6860
rect 23382 6848 23388 6860
rect 22980 6820 23388 6848
rect 22980 6808 22986 6820
rect 23382 6808 23388 6820
rect 23440 6808 23446 6860
rect 23750 6808 23756 6860
rect 23808 6848 23814 6860
rect 24394 6848 24400 6860
rect 23808 6820 24400 6848
rect 23808 6808 23814 6820
rect 24394 6808 24400 6820
rect 24452 6848 24458 6860
rect 26528 6857 26556 6888
rect 24857 6851 24915 6857
rect 24857 6848 24869 6851
rect 24452 6820 24869 6848
rect 24452 6808 24458 6820
rect 24857 6817 24869 6820
rect 24903 6817 24915 6851
rect 24857 6811 24915 6817
rect 26513 6851 26571 6857
rect 26513 6817 26525 6851
rect 26559 6848 26571 6851
rect 26970 6848 26976 6860
rect 26559 6820 26976 6848
rect 26559 6817 26571 6820
rect 26513 6811 26571 6817
rect 26970 6808 26976 6820
rect 27028 6808 27034 6860
rect 19153 6783 19211 6789
rect 19153 6749 19165 6783
rect 19199 6749 19211 6783
rect 19153 6743 19211 6749
rect 18601 6715 18659 6721
rect 18601 6681 18613 6715
rect 18647 6681 18659 6715
rect 18601 6675 18659 6681
rect 18690 6672 18696 6724
rect 18748 6712 18754 6724
rect 19168 6712 19196 6743
rect 22554 6740 22560 6792
rect 22612 6780 22618 6792
rect 23017 6783 23075 6789
rect 23017 6780 23029 6783
rect 22612 6752 23029 6780
rect 22612 6740 22618 6752
rect 23017 6749 23029 6752
rect 23063 6749 23075 6783
rect 25038 6780 25044 6792
rect 24999 6752 25044 6780
rect 23017 6743 23075 6749
rect 25038 6740 25044 6752
rect 25096 6740 25102 6792
rect 18748 6684 19196 6712
rect 18748 6672 18754 6684
rect 21634 6672 21640 6724
rect 21692 6712 21698 6724
rect 22465 6715 22523 6721
rect 22465 6712 22477 6715
rect 21692 6684 22477 6712
rect 21692 6672 21698 6684
rect 22465 6681 22477 6684
rect 22511 6681 22523 6715
rect 22465 6675 22523 6681
rect 24397 6715 24455 6721
rect 24397 6681 24409 6715
rect 24443 6712 24455 6715
rect 24486 6712 24492 6724
rect 24443 6684 24492 6712
rect 24443 6681 24455 6684
rect 24397 6675 24455 6681
rect 24486 6672 24492 6684
rect 24544 6672 24550 6724
rect 26694 6712 26700 6724
rect 26655 6684 26700 6712
rect 26694 6672 26700 6684
rect 26752 6672 26758 6724
rect 2409 6647 2467 6653
rect 2409 6613 2421 6647
rect 2455 6644 2467 6647
rect 2682 6644 2688 6656
rect 2455 6616 2688 6644
rect 2455 6613 2467 6616
rect 2409 6607 2467 6613
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 3602 6604 3608 6656
rect 3660 6644 3666 6656
rect 4065 6647 4123 6653
rect 4065 6644 4077 6647
rect 3660 6616 4077 6644
rect 3660 6604 3666 6616
rect 4065 6613 4077 6616
rect 4111 6613 4123 6647
rect 4065 6607 4123 6613
rect 5169 6647 5227 6653
rect 5169 6613 5181 6647
rect 5215 6644 5227 6647
rect 5442 6644 5448 6656
rect 5215 6616 5448 6644
rect 5215 6613 5227 6616
rect 5169 6607 5227 6613
rect 5442 6604 5448 6616
rect 5500 6644 5506 6656
rect 5813 6647 5871 6653
rect 5813 6644 5825 6647
rect 5500 6616 5825 6644
rect 5500 6604 5506 6616
rect 5813 6613 5825 6616
rect 5859 6613 5871 6647
rect 7282 6644 7288 6656
rect 7243 6616 7288 6644
rect 5813 6607 5871 6613
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 8754 6644 8760 6656
rect 8715 6616 8760 6644
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 9674 6644 9680 6656
rect 9635 6616 9680 6644
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 11054 6604 11060 6656
rect 11112 6644 11118 6656
rect 12161 6647 12219 6653
rect 12161 6644 12173 6647
rect 11112 6616 12173 6644
rect 11112 6604 11118 6616
rect 12161 6613 12173 6616
rect 12207 6613 12219 6647
rect 12161 6607 12219 6613
rect 16390 6604 16396 6656
rect 16448 6644 16454 6656
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 16448 6616 17049 6644
rect 16448 6604 16454 6616
rect 17037 6613 17049 6616
rect 17083 6613 17095 6647
rect 17037 6607 17095 6613
rect 20625 6647 20683 6653
rect 20625 6613 20637 6647
rect 20671 6644 20683 6647
rect 21082 6644 21088 6656
rect 20671 6616 21088 6644
rect 20671 6613 20683 6616
rect 20625 6607 20683 6613
rect 21082 6604 21088 6616
rect 21140 6604 21146 6656
rect 26237 6647 26295 6653
rect 26237 6613 26249 6647
rect 26283 6644 26295 6647
rect 26786 6644 26792 6656
rect 26283 6616 26792 6644
rect 26283 6613 26295 6616
rect 26237 6607 26295 6613
rect 26786 6604 26792 6616
rect 26844 6604 26850 6656
rect 1104 6554 28888 6576
rect 1104 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 15982 6554
rect 16034 6502 16046 6554
rect 16098 6502 16110 6554
rect 16162 6502 16174 6554
rect 16226 6502 25982 6554
rect 26034 6502 26046 6554
rect 26098 6502 26110 6554
rect 26162 6502 26174 6554
rect 26226 6502 28888 6554
rect 1104 6480 28888 6502
rect 2038 6440 2044 6452
rect 1999 6412 2044 6440
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 2130 6400 2136 6452
rect 2188 6440 2194 6452
rect 2317 6443 2375 6449
rect 2317 6440 2329 6443
rect 2188 6412 2329 6440
rect 2188 6400 2194 6412
rect 2317 6409 2329 6412
rect 2363 6409 2375 6443
rect 2317 6403 2375 6409
rect 5810 6400 5816 6452
rect 5868 6440 5874 6452
rect 5997 6443 6055 6449
rect 5997 6440 6009 6443
rect 5868 6412 6009 6440
rect 5868 6400 5874 6412
rect 5997 6409 6009 6412
rect 6043 6409 6055 6443
rect 5997 6403 6055 6409
rect 9033 6443 9091 6449
rect 9033 6409 9045 6443
rect 9079 6440 9091 6443
rect 9953 6443 10011 6449
rect 9953 6440 9965 6443
rect 9079 6412 9965 6440
rect 9079 6409 9091 6412
rect 9033 6403 9091 6409
rect 9953 6409 9965 6412
rect 9999 6440 10011 6443
rect 10134 6440 10140 6452
rect 9999 6412 10140 6440
rect 9999 6409 10011 6412
rect 9953 6403 10011 6409
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 11054 6440 11060 6452
rect 11015 6412 11060 6440
rect 11054 6400 11060 6412
rect 11112 6400 11118 6452
rect 12713 6443 12771 6449
rect 12713 6409 12725 6443
rect 12759 6440 12771 6443
rect 12894 6440 12900 6452
rect 12759 6412 12900 6440
rect 12759 6409 12771 6412
rect 12713 6403 12771 6409
rect 12894 6400 12900 6412
rect 12952 6400 12958 6452
rect 13078 6440 13084 6452
rect 13039 6412 13084 6440
rect 13078 6400 13084 6412
rect 13136 6400 13142 6452
rect 17494 6440 17500 6452
rect 17455 6412 17500 6440
rect 17494 6400 17500 6412
rect 17552 6440 17558 6452
rect 18049 6443 18107 6449
rect 18049 6440 18061 6443
rect 17552 6412 18061 6440
rect 17552 6400 17558 6412
rect 18049 6409 18061 6412
rect 18095 6409 18107 6443
rect 19058 6440 19064 6452
rect 19019 6412 19064 6440
rect 18049 6403 18107 6409
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 19334 6400 19340 6452
rect 19392 6440 19398 6452
rect 19429 6443 19487 6449
rect 19429 6440 19441 6443
rect 19392 6412 19441 6440
rect 19392 6400 19398 6412
rect 19429 6409 19441 6412
rect 19475 6409 19487 6443
rect 20438 6440 20444 6452
rect 20399 6412 20444 6440
rect 19429 6403 19487 6409
rect 20438 6400 20444 6412
rect 20496 6400 20502 6452
rect 22554 6440 22560 6452
rect 22515 6412 22560 6440
rect 22554 6400 22560 6412
rect 22612 6400 22618 6452
rect 22922 6440 22928 6452
rect 22883 6412 22928 6440
rect 22922 6400 22928 6412
rect 22980 6400 22986 6452
rect 23198 6440 23204 6452
rect 23159 6412 23204 6440
rect 23198 6400 23204 6412
rect 23256 6400 23262 6452
rect 24394 6440 24400 6452
rect 24355 6412 24400 6440
rect 24394 6400 24400 6412
rect 24452 6440 24458 6452
rect 24670 6440 24676 6452
rect 24452 6412 24676 6440
rect 24452 6400 24458 6412
rect 24670 6400 24676 6412
rect 24728 6400 24734 6452
rect 25038 6400 25044 6452
rect 25096 6440 25102 6452
rect 25225 6443 25283 6449
rect 25225 6440 25237 6443
rect 25096 6412 25237 6440
rect 25096 6400 25102 6412
rect 25225 6409 25237 6412
rect 25271 6440 25283 6443
rect 26786 6440 26792 6452
rect 25271 6412 26792 6440
rect 25271 6409 25283 6412
rect 25225 6403 25283 6409
rect 26786 6400 26792 6412
rect 26844 6400 26850 6452
rect 26970 6440 26976 6452
rect 26931 6412 26976 6440
rect 26970 6400 26976 6412
rect 27028 6400 27034 6452
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 4985 6375 5043 6381
rect 4985 6372 4997 6375
rect 4120 6344 4997 6372
rect 4120 6332 4126 6344
rect 4985 6341 4997 6344
rect 5031 6341 5043 6375
rect 4985 6335 5043 6341
rect 9769 6375 9827 6381
rect 9769 6341 9781 6375
rect 9815 6372 9827 6375
rect 10226 6372 10232 6384
rect 9815 6344 10232 6372
rect 9815 6341 9827 6344
rect 9769 6335 9827 6341
rect 10226 6332 10232 6344
rect 10284 6332 10290 6384
rect 15749 6375 15807 6381
rect 15749 6341 15761 6375
rect 15795 6372 15807 6375
rect 17129 6375 17187 6381
rect 17129 6372 17141 6375
rect 15795 6344 17141 6372
rect 15795 6341 15807 6344
rect 15749 6335 15807 6341
rect 3694 6304 3700 6316
rect 3655 6276 3700 6304
rect 3694 6264 3700 6276
rect 3752 6264 3758 6316
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6273 3939 6307
rect 5442 6304 5448 6316
rect 5403 6276 5448 6304
rect 3881 6267 3939 6273
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2038 6236 2044 6248
rect 1443 6208 2044 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2038 6196 2044 6208
rect 2096 6196 2102 6248
rect 2777 6239 2835 6245
rect 2777 6205 2789 6239
rect 2823 6236 2835 6239
rect 3602 6236 3608 6248
rect 2823 6208 3608 6236
rect 2823 6205 2835 6208
rect 2777 6199 2835 6205
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 3896 6236 3924 6267
rect 5442 6264 5448 6276
rect 5500 6264 5506 6316
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6304 6699 6307
rect 7650 6304 7656 6316
rect 6687 6276 7512 6304
rect 7611 6276 7656 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 5074 6236 5080 6248
rect 3896 6208 5080 6236
rect 2866 6128 2872 6180
rect 2924 6168 2930 6180
rect 3145 6171 3203 6177
rect 3145 6168 3157 6171
rect 2924 6140 3157 6168
rect 2924 6128 2930 6140
rect 3145 6137 3157 6140
rect 3191 6168 3203 6171
rect 3896 6168 3924 6208
rect 5074 6196 5080 6208
rect 5132 6236 5138 6248
rect 5552 6236 5580 6267
rect 5132 6208 5580 6236
rect 5132 6196 5138 6208
rect 7282 6196 7288 6248
rect 7340 6236 7346 6248
rect 7484 6245 7512 6276
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 9582 6264 9588 6316
rect 9640 6304 9646 6316
rect 10505 6307 10563 6313
rect 10505 6304 10517 6307
rect 9640 6276 10517 6304
rect 9640 6264 9646 6276
rect 10505 6273 10517 6276
rect 10551 6304 10563 6307
rect 12161 6307 12219 6313
rect 12161 6304 12173 6307
rect 10551 6276 12173 6304
rect 10551 6273 10563 6276
rect 10505 6267 10563 6273
rect 12161 6273 12173 6276
rect 12207 6304 12219 6307
rect 12802 6304 12808 6316
rect 12207 6276 12808 6304
rect 12207 6273 12219 6276
rect 12161 6267 12219 6273
rect 12802 6264 12808 6276
rect 12860 6264 12866 6316
rect 15381 6307 15439 6313
rect 15381 6273 15393 6307
rect 15427 6304 15439 6307
rect 16298 6304 16304 6316
rect 15427 6276 16304 6304
rect 15427 6273 15439 6276
rect 15381 6267 15439 6273
rect 16298 6264 16304 6276
rect 16356 6264 16362 6316
rect 16500 6313 16528 6344
rect 17129 6341 17141 6344
rect 17175 6372 17187 6375
rect 17218 6372 17224 6384
rect 17175 6344 17224 6372
rect 17175 6341 17187 6344
rect 17129 6335 17187 6341
rect 17218 6332 17224 6344
rect 17276 6372 17282 6384
rect 17586 6372 17592 6384
rect 17276 6344 17592 6372
rect 17276 6332 17282 6344
rect 17586 6332 17592 6344
rect 17644 6332 17650 6384
rect 16485 6307 16543 6313
rect 16485 6273 16497 6307
rect 16531 6273 16543 6307
rect 16485 6267 16543 6273
rect 18138 6264 18144 6316
rect 18196 6304 18202 6316
rect 18598 6304 18604 6316
rect 18196 6276 18604 6304
rect 18196 6264 18202 6276
rect 18598 6264 18604 6276
rect 18656 6264 18662 6316
rect 21082 6304 21088 6316
rect 21043 6276 21088 6304
rect 21082 6264 21088 6276
rect 21140 6264 21146 6316
rect 26234 6304 26240 6316
rect 26195 6276 26240 6304
rect 26234 6264 26240 6276
rect 26292 6304 26298 6316
rect 26292 6276 26464 6304
rect 26292 6264 26298 6276
rect 7377 6239 7435 6245
rect 7377 6236 7389 6239
rect 7340 6208 7389 6236
rect 7340 6196 7346 6208
rect 7377 6205 7389 6208
rect 7423 6205 7435 6239
rect 7377 6199 7435 6205
rect 7469 6239 7527 6245
rect 7469 6205 7481 6239
rect 7515 6236 7527 6239
rect 7834 6236 7840 6248
rect 7515 6208 7840 6236
rect 7515 6205 7527 6208
rect 7469 6199 7527 6205
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 17865 6239 17923 6245
rect 17865 6205 17877 6239
rect 17911 6236 17923 6239
rect 18414 6236 18420 6248
rect 17911 6208 18420 6236
rect 17911 6205 17923 6208
rect 17865 6199 17923 6205
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 20438 6196 20444 6248
rect 20496 6236 20502 6248
rect 26436 6245 26464 6276
rect 20993 6239 21051 6245
rect 20993 6236 21005 6239
rect 20496 6208 21005 6236
rect 20496 6196 20502 6208
rect 20993 6205 21005 6208
rect 21039 6205 21051 6239
rect 20993 6199 21051 6205
rect 26421 6239 26479 6245
rect 26421 6205 26433 6239
rect 26467 6205 26479 6239
rect 26421 6199 26479 6205
rect 3191 6140 3924 6168
rect 5353 6171 5411 6177
rect 3191 6137 3203 6140
rect 3145 6131 3203 6137
rect 5353 6137 5365 6171
rect 5399 6168 5411 6171
rect 5442 6168 5448 6180
rect 5399 6140 5448 6168
rect 5399 6137 5411 6140
rect 5353 6131 5411 6137
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 9401 6171 9459 6177
rect 9401 6137 9413 6171
rect 9447 6168 9459 6171
rect 10413 6171 10471 6177
rect 10413 6168 10425 6171
rect 9447 6140 10425 6168
rect 9447 6137 9459 6140
rect 9401 6131 9459 6137
rect 10413 6137 10425 6140
rect 10459 6168 10471 6171
rect 10778 6168 10784 6180
rect 10459 6140 10784 6168
rect 10459 6137 10471 6140
rect 10413 6131 10471 6137
rect 10778 6128 10784 6140
rect 10836 6128 10842 6180
rect 15013 6171 15071 6177
rect 15013 6137 15025 6171
rect 15059 6168 15071 6171
rect 15746 6168 15752 6180
rect 15059 6140 15752 6168
rect 15059 6137 15071 6140
rect 15013 6131 15071 6137
rect 15746 6128 15752 6140
rect 15804 6168 15810 6180
rect 16209 6171 16267 6177
rect 16209 6168 16221 6171
rect 15804 6140 16221 6168
rect 15804 6128 15810 6140
rect 16209 6137 16221 6140
rect 16255 6137 16267 6171
rect 16209 6131 16267 6137
rect 1394 6060 1400 6112
rect 1452 6100 1458 6112
rect 1581 6103 1639 6109
rect 1581 6100 1593 6103
rect 1452 6072 1593 6100
rect 1452 6060 1458 6072
rect 1581 6069 1593 6072
rect 1627 6069 1639 6103
rect 3234 6100 3240 6112
rect 3195 6072 3240 6100
rect 1581 6063 1639 6069
rect 3234 6060 3240 6072
rect 3292 6060 3298 6112
rect 4338 6100 4344 6112
rect 4299 6072 4344 6100
rect 4338 6060 4344 6072
rect 4396 6060 4402 6112
rect 4706 6100 4712 6112
rect 4667 6072 4712 6100
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 7009 6103 7067 6109
rect 7009 6069 7021 6103
rect 7055 6100 7067 6103
rect 7374 6100 7380 6112
rect 7055 6072 7380 6100
rect 7055 6069 7067 6072
rect 7009 6063 7067 6069
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 7650 6060 7656 6112
rect 7708 6100 7714 6112
rect 8021 6103 8079 6109
rect 8021 6100 8033 6103
rect 7708 6072 8033 6100
rect 7708 6060 7714 6072
rect 8021 6069 8033 6072
rect 8067 6069 8079 6103
rect 10318 6100 10324 6112
rect 10279 6072 10324 6100
rect 8021 6063 8079 6069
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 15838 6100 15844 6112
rect 15799 6072 15844 6100
rect 15838 6060 15844 6072
rect 15896 6060 15902 6112
rect 17954 6060 17960 6112
rect 18012 6100 18018 6112
rect 18506 6100 18512 6112
rect 18012 6072 18512 6100
rect 18012 6060 18018 6072
rect 18506 6060 18512 6072
rect 18564 6060 18570 6112
rect 20530 6100 20536 6112
rect 20491 6072 20536 6100
rect 20530 6060 20536 6072
rect 20588 6060 20594 6112
rect 20806 6060 20812 6112
rect 20864 6100 20870 6112
rect 20901 6103 20959 6109
rect 20901 6100 20913 6103
rect 20864 6072 20913 6100
rect 20864 6060 20870 6072
rect 20901 6069 20913 6072
rect 20947 6069 20959 6103
rect 24762 6100 24768 6112
rect 24723 6072 24768 6100
rect 20901 6063 20959 6069
rect 24762 6060 24768 6072
rect 24820 6060 24826 6112
rect 26602 6100 26608 6112
rect 26563 6072 26608 6100
rect 26602 6060 26608 6072
rect 26660 6060 26666 6112
rect 1104 6010 28888 6032
rect 1104 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 20982 6010
rect 21034 5958 21046 6010
rect 21098 5958 21110 6010
rect 21162 5958 21174 6010
rect 21226 5958 28888 6010
rect 1104 5936 28888 5958
rect 4341 5899 4399 5905
rect 4341 5865 4353 5899
rect 4387 5896 4399 5899
rect 4614 5896 4620 5908
rect 4387 5868 4620 5896
rect 4387 5865 4399 5868
rect 4341 5859 4399 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5074 5896 5080 5908
rect 5035 5868 5080 5896
rect 5074 5856 5080 5868
rect 5132 5856 5138 5908
rect 5442 5896 5448 5908
rect 5403 5868 5448 5896
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 5905 5899 5963 5905
rect 5905 5865 5917 5899
rect 5951 5896 5963 5899
rect 6270 5896 6276 5908
rect 5951 5868 6276 5896
rect 5951 5865 5963 5868
rect 5905 5859 5963 5865
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 9582 5856 9588 5908
rect 9640 5896 9646 5908
rect 9953 5899 10011 5905
rect 9953 5896 9965 5899
rect 9640 5868 9965 5896
rect 9640 5856 9646 5868
rect 9953 5865 9965 5868
rect 9999 5865 10011 5899
rect 10318 5896 10324 5908
rect 10279 5868 10324 5896
rect 9953 5859 10011 5865
rect 10318 5856 10324 5868
rect 10376 5896 10382 5908
rect 10597 5899 10655 5905
rect 10597 5896 10609 5899
rect 10376 5868 10609 5896
rect 10376 5856 10382 5868
rect 10597 5865 10609 5868
rect 10643 5865 10655 5899
rect 10597 5859 10655 5865
rect 10686 5856 10692 5908
rect 10744 5896 10750 5908
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 10744 5868 11069 5896
rect 10744 5856 10750 5868
rect 11057 5865 11069 5868
rect 11103 5896 11115 5899
rect 12161 5899 12219 5905
rect 12161 5896 12173 5899
rect 11103 5868 12173 5896
rect 11103 5865 11115 5868
rect 11057 5859 11115 5865
rect 12161 5865 12173 5868
rect 12207 5865 12219 5899
rect 12161 5859 12219 5865
rect 12342 5856 12348 5908
rect 12400 5896 12406 5908
rect 12621 5899 12679 5905
rect 12621 5896 12633 5899
rect 12400 5868 12633 5896
rect 12400 5856 12406 5868
rect 12621 5865 12633 5868
rect 12667 5896 12679 5899
rect 12710 5896 12716 5908
rect 12667 5868 12716 5896
rect 12667 5865 12679 5868
rect 12621 5859 12679 5865
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 17218 5896 17224 5908
rect 17179 5868 17224 5896
rect 17218 5856 17224 5868
rect 17276 5856 17282 5908
rect 17954 5856 17960 5908
rect 18012 5896 18018 5908
rect 18049 5899 18107 5905
rect 18049 5896 18061 5899
rect 18012 5868 18061 5896
rect 18012 5856 18018 5868
rect 18049 5865 18061 5868
rect 18095 5865 18107 5899
rect 18598 5896 18604 5908
rect 18559 5868 18604 5896
rect 18049 5859 18107 5865
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 19242 5856 19248 5908
rect 19300 5896 19306 5908
rect 19613 5899 19671 5905
rect 19613 5896 19625 5899
rect 19300 5868 19625 5896
rect 19300 5856 19306 5868
rect 19613 5865 19625 5868
rect 19659 5896 19671 5899
rect 20530 5896 20536 5908
rect 19659 5868 20536 5896
rect 19659 5865 19671 5868
rect 19613 5859 19671 5865
rect 20530 5856 20536 5868
rect 20588 5856 20594 5908
rect 20625 5899 20683 5905
rect 20625 5865 20637 5899
rect 20671 5896 20683 5899
rect 20806 5896 20812 5908
rect 20671 5868 20812 5896
rect 20671 5865 20683 5868
rect 20625 5859 20683 5865
rect 20806 5856 20812 5868
rect 20864 5896 20870 5908
rect 20901 5899 20959 5905
rect 20901 5896 20913 5899
rect 20864 5868 20913 5896
rect 20864 5856 20870 5868
rect 20901 5865 20913 5868
rect 20947 5865 20959 5899
rect 20901 5859 20959 5865
rect 1756 5831 1814 5837
rect 1756 5797 1768 5831
rect 1802 5828 1814 5831
rect 2774 5828 2780 5840
rect 1802 5800 2780 5828
rect 1802 5797 1814 5800
rect 1756 5791 1814 5797
rect 2774 5788 2780 5800
rect 2832 5788 2838 5840
rect 4632 5828 4660 5856
rect 6181 5831 6239 5837
rect 6181 5828 6193 5831
rect 4632 5800 6193 5828
rect 6181 5797 6193 5800
rect 6227 5797 6239 5831
rect 6181 5791 6239 5797
rect 7377 5831 7435 5837
rect 7377 5797 7389 5831
rect 7423 5828 7435 5831
rect 7742 5828 7748 5840
rect 7423 5800 7748 5828
rect 7423 5797 7435 5800
rect 7377 5791 7435 5797
rect 7742 5788 7748 5800
rect 7800 5788 7806 5840
rect 12526 5828 12532 5840
rect 12487 5800 12532 5828
rect 12526 5788 12532 5800
rect 12584 5788 12590 5840
rect 16108 5831 16166 5837
rect 16108 5797 16120 5831
rect 16154 5828 16166 5831
rect 16298 5828 16304 5840
rect 16154 5800 16304 5828
rect 16154 5797 16166 5800
rect 16108 5791 16166 5797
rect 16298 5788 16304 5800
rect 16356 5828 16362 5840
rect 16482 5828 16488 5840
rect 16356 5800 16488 5828
rect 16356 5788 16362 5800
rect 16482 5788 16488 5800
rect 16540 5788 16546 5840
rect 1489 5763 1547 5769
rect 1489 5729 1501 5763
rect 1535 5760 1547 5763
rect 2682 5760 2688 5772
rect 1535 5732 2688 5760
rect 1535 5729 1547 5732
rect 1489 5723 1547 5729
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 7466 5720 7472 5772
rect 7524 5760 7530 5772
rect 10962 5760 10968 5772
rect 7524 5732 7569 5760
rect 10923 5732 10968 5760
rect 7524 5720 7530 5732
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 13262 5760 13268 5772
rect 12492 5732 13268 5760
rect 12492 5720 12498 5732
rect 13262 5720 13268 5732
rect 13320 5760 13326 5772
rect 13633 5763 13691 5769
rect 13633 5760 13645 5763
rect 13320 5732 13645 5760
rect 13320 5720 13326 5732
rect 13633 5729 13645 5732
rect 13679 5729 13691 5763
rect 13633 5723 13691 5729
rect 15654 5720 15660 5772
rect 15712 5760 15718 5772
rect 15841 5763 15899 5769
rect 15841 5760 15853 5763
rect 15712 5732 15853 5760
rect 15712 5720 15718 5732
rect 15841 5729 15853 5732
rect 15887 5729 15899 5763
rect 15841 5723 15899 5729
rect 22462 5720 22468 5772
rect 22520 5760 22526 5772
rect 22629 5763 22687 5769
rect 22629 5760 22641 5763
rect 22520 5732 22641 5760
rect 22520 5720 22526 5732
rect 22629 5729 22641 5732
rect 22675 5729 22687 5763
rect 26510 5760 26516 5772
rect 26471 5732 26516 5760
rect 22629 5723 22687 5729
rect 26510 5720 26516 5732
rect 26568 5720 26574 5772
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 7484 5692 7512 5720
rect 7650 5692 7656 5704
rect 6972 5664 7512 5692
rect 7611 5664 7656 5692
rect 6972 5652 6978 5664
rect 7650 5652 7656 5664
rect 7708 5652 7714 5704
rect 11241 5695 11299 5701
rect 11241 5661 11253 5695
rect 11287 5692 11299 5695
rect 11514 5692 11520 5704
rect 11287 5664 11520 5692
rect 11287 5661 11299 5664
rect 11241 5655 11299 5661
rect 11514 5652 11520 5664
rect 11572 5652 11578 5704
rect 12805 5695 12863 5701
rect 12805 5661 12817 5695
rect 12851 5692 12863 5695
rect 19702 5692 19708 5704
rect 12851 5664 13400 5692
rect 19663 5664 19708 5692
rect 12851 5661 12863 5664
rect 12805 5655 12863 5661
rect 2866 5556 2872 5568
rect 2827 5528 2872 5556
rect 2866 5516 2872 5528
rect 2924 5516 2930 5568
rect 7006 5556 7012 5568
rect 6967 5528 7012 5556
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 13372 5565 13400 5664
rect 19702 5652 19708 5664
rect 19760 5652 19766 5704
rect 19797 5695 19855 5701
rect 19797 5661 19809 5695
rect 19843 5661 19855 5695
rect 19797 5655 19855 5661
rect 19426 5584 19432 5636
rect 19484 5624 19490 5636
rect 19812 5624 19840 5655
rect 22370 5652 22376 5704
rect 22428 5692 22434 5704
rect 22428 5664 22473 5692
rect 22428 5652 22434 5664
rect 23842 5652 23848 5704
rect 23900 5692 23906 5704
rect 27430 5692 27436 5704
rect 23900 5664 27436 5692
rect 23900 5652 23906 5664
rect 27430 5652 27436 5664
rect 27488 5652 27494 5704
rect 19484 5596 19840 5624
rect 19484 5584 19490 5596
rect 13357 5559 13415 5565
rect 13357 5525 13369 5559
rect 13403 5556 13415 5559
rect 13630 5556 13636 5568
rect 13403 5528 13636 5556
rect 13403 5525 13415 5528
rect 13357 5519 13415 5525
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 19245 5559 19303 5565
rect 19245 5525 19257 5559
rect 19291 5556 19303 5559
rect 19334 5556 19340 5568
rect 19291 5528 19340 5556
rect 19291 5525 19303 5528
rect 19245 5519 19303 5525
rect 19334 5516 19340 5528
rect 19392 5516 19398 5568
rect 23753 5559 23811 5565
rect 23753 5525 23765 5559
rect 23799 5556 23811 5559
rect 23842 5556 23848 5568
rect 23799 5528 23848 5556
rect 23799 5525 23811 5528
rect 23753 5519 23811 5525
rect 23842 5516 23848 5528
rect 23900 5516 23906 5568
rect 25498 5556 25504 5568
rect 25459 5528 25504 5556
rect 25498 5516 25504 5528
rect 25556 5516 25562 5568
rect 26694 5556 26700 5568
rect 26655 5528 26700 5556
rect 26694 5516 26700 5528
rect 26752 5516 26758 5568
rect 1104 5466 28888 5488
rect 1104 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 15982 5466
rect 16034 5414 16046 5466
rect 16098 5414 16110 5466
rect 16162 5414 16174 5466
rect 16226 5414 25982 5466
rect 26034 5414 26046 5466
rect 26098 5414 26110 5466
rect 26162 5414 26174 5466
rect 26226 5414 28888 5466
rect 1104 5392 28888 5414
rect 1578 5352 1584 5364
rect 1539 5324 1584 5352
rect 1578 5312 1584 5324
rect 1636 5312 1642 5364
rect 2777 5355 2835 5361
rect 2777 5321 2789 5355
rect 2823 5352 2835 5355
rect 2866 5352 2872 5364
rect 2823 5324 2872 5352
rect 2823 5321 2835 5324
rect 2777 5315 2835 5321
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 3973 5355 4031 5361
rect 3973 5321 3985 5355
rect 4019 5352 4031 5355
rect 4062 5352 4068 5364
rect 4019 5324 4068 5352
rect 4019 5321 4031 5324
rect 3973 5315 4031 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 6638 5352 6644 5364
rect 6551 5324 6644 5352
rect 6638 5312 6644 5324
rect 6696 5352 6702 5364
rect 6914 5352 6920 5364
rect 6696 5324 6920 5352
rect 6696 5312 6702 5324
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 7653 5355 7711 5361
rect 7653 5321 7665 5355
rect 7699 5352 7711 5355
rect 7742 5352 7748 5364
rect 7699 5324 7748 5352
rect 7699 5321 7711 5324
rect 7653 5315 7711 5321
rect 7742 5312 7748 5324
rect 7800 5312 7806 5364
rect 10778 5352 10784 5364
rect 10739 5324 10784 5352
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 12342 5352 12348 5364
rect 12299 5324 12348 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 12526 5312 12532 5364
rect 12584 5352 12590 5364
rect 12621 5355 12679 5361
rect 12621 5352 12633 5355
rect 12584 5324 12633 5352
rect 12584 5312 12590 5324
rect 12621 5321 12633 5324
rect 12667 5321 12679 5355
rect 14642 5352 14648 5364
rect 14603 5324 14648 5352
rect 12621 5315 12679 5321
rect 14642 5312 14648 5324
rect 14700 5312 14706 5364
rect 15746 5312 15752 5364
rect 15804 5352 15810 5364
rect 16025 5355 16083 5361
rect 16025 5352 16037 5355
rect 15804 5324 16037 5352
rect 15804 5312 15810 5324
rect 16025 5321 16037 5324
rect 16071 5321 16083 5355
rect 16025 5315 16083 5321
rect 16298 5312 16304 5364
rect 16356 5352 16362 5364
rect 17037 5355 17095 5361
rect 17037 5352 17049 5355
rect 16356 5324 17049 5352
rect 16356 5312 16362 5324
rect 2884 5284 2912 5312
rect 10689 5287 10747 5293
rect 2884 5256 3464 5284
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5216 2467 5219
rect 2774 5216 2780 5228
rect 2455 5188 2780 5216
rect 2455 5185 2467 5188
rect 2409 5179 2467 5185
rect 2774 5176 2780 5188
rect 2832 5176 2838 5228
rect 3234 5176 3240 5228
rect 3292 5216 3298 5228
rect 3436 5225 3464 5256
rect 10689 5253 10701 5287
rect 10735 5284 10747 5287
rect 10962 5284 10968 5296
rect 10735 5256 10968 5284
rect 10735 5253 10747 5256
rect 10689 5247 10747 5253
rect 10962 5244 10968 5256
rect 11020 5244 11026 5296
rect 15565 5287 15623 5293
rect 15565 5253 15577 5287
rect 15611 5284 15623 5287
rect 16316 5284 16344 5312
rect 15611 5256 16344 5284
rect 15611 5253 15623 5256
rect 15565 5247 15623 5253
rect 3329 5219 3387 5225
rect 3329 5216 3341 5219
rect 3292 5188 3341 5216
rect 3292 5176 3298 5188
rect 3329 5185 3341 5188
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 3421 5219 3479 5225
rect 3421 5185 3433 5219
rect 3467 5185 3479 5219
rect 3421 5179 3479 5185
rect 7101 5219 7159 5225
rect 7101 5185 7113 5219
rect 7147 5216 7159 5219
rect 7282 5216 7288 5228
rect 7147 5188 7288 5216
rect 7147 5185 7159 5188
rect 7101 5179 7159 5185
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 10321 5219 10379 5225
rect 10321 5185 10333 5219
rect 10367 5216 10379 5219
rect 11425 5219 11483 5225
rect 11425 5216 11437 5219
rect 10367 5188 11437 5216
rect 10367 5185 10379 5188
rect 10321 5179 10379 5185
rect 11425 5185 11437 5188
rect 11471 5216 11483 5219
rect 11514 5216 11520 5228
rect 11471 5188 11520 5216
rect 11471 5185 11483 5188
rect 11425 5179 11483 5185
rect 11514 5176 11520 5188
rect 11572 5176 11578 5228
rect 13262 5216 13268 5228
rect 13223 5188 13268 5216
rect 13262 5176 13268 5188
rect 13320 5176 13326 5228
rect 16684 5225 16712 5324
rect 17037 5321 17049 5324
rect 17083 5321 17095 5355
rect 17037 5315 17095 5321
rect 18969 5355 19027 5361
rect 18969 5321 18981 5355
rect 19015 5352 19027 5355
rect 19242 5352 19248 5364
rect 19015 5324 19248 5352
rect 19015 5321 19027 5324
rect 18969 5315 19027 5321
rect 19242 5312 19248 5324
rect 19300 5312 19306 5364
rect 19702 5352 19708 5364
rect 19663 5324 19708 5352
rect 19702 5312 19708 5324
rect 19760 5352 19766 5364
rect 20533 5355 20591 5361
rect 20533 5352 20545 5355
rect 19760 5324 20545 5352
rect 19760 5312 19766 5324
rect 20533 5321 20545 5324
rect 20579 5321 20591 5355
rect 20533 5315 20591 5321
rect 26510 5312 26516 5364
rect 26568 5352 26574 5364
rect 27341 5355 27399 5361
rect 27341 5352 27353 5355
rect 26568 5324 27353 5352
rect 26568 5312 26574 5324
rect 27341 5321 27353 5324
rect 27387 5321 27399 5355
rect 27341 5315 27399 5321
rect 20073 5287 20131 5293
rect 20073 5253 20085 5287
rect 20119 5284 20131 5287
rect 22462 5284 22468 5296
rect 20119 5256 21220 5284
rect 22423 5256 22468 5284
rect 20119 5253 20131 5256
rect 20073 5247 20131 5253
rect 16669 5219 16727 5225
rect 16669 5185 16681 5219
rect 16715 5185 16727 5219
rect 20346 5216 20352 5228
rect 20307 5188 20352 5216
rect 16669 5179 16727 5185
rect 20346 5176 20352 5188
rect 20404 5216 20410 5228
rect 21192 5225 21220 5256
rect 22462 5244 22468 5256
rect 22520 5244 22526 5296
rect 26786 5284 26792 5296
rect 26747 5256 26792 5284
rect 26786 5244 26792 5256
rect 26844 5244 26850 5296
rect 21177 5219 21235 5225
rect 20404 5188 20944 5216
rect 20404 5176 20410 5188
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 8110 5148 8116 5160
rect 1443 5120 2084 5148
rect 8071 5120 8116 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 2056 5021 2084 5120
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 15194 5108 15200 5160
rect 15252 5148 15258 5160
rect 15933 5151 15991 5157
rect 15933 5148 15945 5151
rect 15252 5120 15945 5148
rect 15252 5108 15258 5120
rect 15933 5117 15945 5120
rect 15979 5148 15991 5151
rect 16393 5151 16451 5157
rect 16393 5148 16405 5151
rect 15979 5120 16405 5148
rect 15979 5117 15991 5120
rect 15933 5111 15991 5117
rect 16393 5117 16405 5120
rect 16439 5148 16451 5151
rect 16482 5148 16488 5160
rect 16439 5120 16488 5148
rect 16439 5117 16451 5120
rect 16393 5111 16451 5117
rect 16482 5108 16488 5120
rect 16540 5108 16546 5160
rect 20916 5157 20944 5188
rect 21177 5185 21189 5219
rect 21223 5216 21235 5219
rect 21266 5216 21272 5228
rect 21223 5188 21272 5216
rect 21223 5185 21235 5188
rect 21177 5179 21235 5185
rect 21266 5176 21272 5188
rect 21324 5216 21330 5228
rect 22480 5216 22508 5244
rect 21324 5188 22508 5216
rect 21324 5176 21330 5188
rect 20901 5151 20959 5157
rect 20901 5117 20913 5151
rect 20947 5117 20959 5151
rect 25409 5151 25467 5157
rect 25409 5148 25421 5151
rect 20901 5111 20959 5117
rect 23584 5120 25421 5148
rect 3237 5083 3295 5089
rect 3237 5049 3249 5083
rect 3283 5080 3295 5083
rect 4062 5080 4068 5092
rect 3283 5052 4068 5080
rect 3283 5049 3295 5052
rect 3237 5043 3295 5049
rect 4062 5040 4068 5052
rect 4120 5040 4126 5092
rect 7650 5080 7656 5092
rect 6196 5052 7656 5080
rect 2041 5015 2099 5021
rect 2041 4981 2053 5015
rect 2087 5012 2099 5015
rect 2130 5012 2136 5024
rect 2087 4984 2136 5012
rect 2087 4981 2099 4984
rect 2041 4975 2099 4981
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 2869 5015 2927 5021
rect 2869 4981 2881 5015
rect 2915 5012 2927 5015
rect 3142 5012 3148 5024
rect 2915 4984 3148 5012
rect 2915 4981 2927 4984
rect 2869 4975 2927 4981
rect 3142 4972 3148 4984
rect 3200 4972 3206 5024
rect 5810 4972 5816 5024
rect 5868 5012 5874 5024
rect 6196 5021 6224 5052
rect 7650 5040 7656 5052
rect 7708 5080 7714 5092
rect 7929 5083 7987 5089
rect 7929 5080 7941 5083
rect 7708 5052 7941 5080
rect 7708 5040 7714 5052
rect 7929 5049 7941 5052
rect 7975 5080 7987 5083
rect 8358 5083 8416 5089
rect 8358 5080 8370 5083
rect 7975 5052 8370 5080
rect 7975 5049 7987 5052
rect 7929 5043 7987 5049
rect 8358 5049 8370 5052
rect 8404 5049 8416 5083
rect 8358 5043 8416 5049
rect 11149 5083 11207 5089
rect 11149 5049 11161 5083
rect 11195 5080 11207 5083
rect 11195 5052 11928 5080
rect 11195 5049 11207 5052
rect 11149 5043 11207 5049
rect 11900 5024 11928 5052
rect 12066 5040 12072 5092
rect 12124 5080 12130 5092
rect 13081 5083 13139 5089
rect 13081 5080 13093 5083
rect 12124 5052 13093 5080
rect 12124 5040 12130 5052
rect 13081 5049 13093 5052
rect 13127 5080 13139 5083
rect 13532 5083 13590 5089
rect 13532 5080 13544 5083
rect 13127 5052 13544 5080
rect 13127 5049 13139 5052
rect 13081 5043 13139 5049
rect 13532 5049 13544 5052
rect 13578 5080 13590 5083
rect 13630 5080 13636 5092
rect 13578 5052 13636 5080
rect 13578 5049 13590 5052
rect 13532 5043 13590 5049
rect 13630 5040 13636 5052
rect 13688 5040 13694 5092
rect 15654 5040 15660 5092
rect 15712 5080 15718 5092
rect 16206 5080 16212 5092
rect 15712 5052 16212 5080
rect 15712 5040 15718 5052
rect 16206 5040 16212 5052
rect 16264 5080 16270 5092
rect 17405 5083 17463 5089
rect 17405 5080 17417 5083
rect 16264 5052 17417 5080
rect 16264 5040 16270 5052
rect 17405 5049 17417 5052
rect 17451 5049 17463 5083
rect 17405 5043 17463 5049
rect 20530 5040 20536 5092
rect 20588 5080 20594 5092
rect 20993 5083 21051 5089
rect 20993 5080 21005 5083
rect 20588 5052 21005 5080
rect 20588 5040 20594 5052
rect 20993 5049 21005 5052
rect 21039 5049 21051 5083
rect 20993 5043 21051 5049
rect 23584 5024 23612 5120
rect 25409 5117 25421 5120
rect 25455 5148 25467 5151
rect 25498 5148 25504 5160
rect 25455 5120 25504 5148
rect 25455 5117 25467 5120
rect 25409 5111 25467 5117
rect 25498 5108 25504 5120
rect 25556 5108 25562 5160
rect 25654 5083 25712 5089
rect 25654 5080 25666 5083
rect 25240 5052 25666 5080
rect 6181 5015 6239 5021
rect 6181 5012 6193 5015
rect 5868 4984 6193 5012
rect 5868 4972 5874 4984
rect 6181 4981 6193 4984
rect 6227 4981 6239 5015
rect 9490 5012 9496 5024
rect 9451 4984 9496 5012
rect 6181 4975 6239 4981
rect 9490 4972 9496 4984
rect 9548 4972 9554 5024
rect 11241 5015 11299 5021
rect 11241 4981 11253 5015
rect 11287 5012 11299 5015
rect 11330 5012 11336 5024
rect 11287 4984 11336 5012
rect 11287 4981 11299 4984
rect 11241 4975 11299 4981
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 11882 5012 11888 5024
rect 11843 4984 11888 5012
rect 11882 4972 11888 4984
rect 11940 4972 11946 5024
rect 16114 4972 16120 5024
rect 16172 5012 16178 5024
rect 16485 5015 16543 5021
rect 16485 5012 16497 5015
rect 16172 4984 16497 5012
rect 16172 4972 16178 4984
rect 16485 4981 16497 4984
rect 16531 5012 16543 5015
rect 16666 5012 16672 5024
rect 16531 4984 16672 5012
rect 16531 4981 16543 4984
rect 16485 4975 16543 4981
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 19337 5015 19395 5021
rect 19337 4981 19349 5015
rect 19383 5012 19395 5015
rect 19426 5012 19432 5024
rect 19383 4984 19432 5012
rect 19383 4981 19395 4984
rect 19337 4975 19395 4981
rect 19426 4972 19432 4984
rect 19484 4972 19490 5024
rect 20162 4972 20168 5024
rect 20220 5012 20226 5024
rect 22370 5012 22376 5024
rect 20220 4984 22376 5012
rect 20220 4972 20226 4984
rect 22370 4972 22376 4984
rect 22428 5012 22434 5024
rect 22741 5015 22799 5021
rect 22741 5012 22753 5015
rect 22428 4984 22753 5012
rect 22428 4972 22434 4984
rect 22741 4981 22753 4984
rect 22787 5012 22799 5015
rect 23566 5012 23572 5024
rect 22787 4984 23572 5012
rect 22787 4981 22799 4984
rect 22741 4975 22799 4981
rect 23566 4972 23572 4984
rect 23624 4972 23630 5024
rect 24946 4972 24952 5024
rect 25004 5012 25010 5024
rect 25240 5021 25268 5052
rect 25654 5049 25666 5052
rect 25700 5049 25712 5083
rect 25654 5043 25712 5049
rect 25225 5015 25283 5021
rect 25225 5012 25237 5015
rect 25004 4984 25237 5012
rect 25004 4972 25010 4984
rect 25225 4981 25237 4984
rect 25271 4981 25283 5015
rect 25225 4975 25283 4981
rect 1104 4922 28888 4944
rect 1104 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 20982 4922
rect 21034 4870 21046 4922
rect 21098 4870 21110 4922
rect 21162 4870 21174 4922
rect 21226 4870 28888 4922
rect 1104 4848 28888 4870
rect 1578 4808 1584 4820
rect 1539 4780 1584 4808
rect 1578 4768 1584 4780
rect 1636 4768 1642 4820
rect 3145 4811 3203 4817
rect 3145 4777 3157 4811
rect 3191 4808 3203 4811
rect 3234 4808 3240 4820
rect 3191 4780 3240 4808
rect 3191 4777 3203 4780
rect 3145 4771 3203 4777
rect 3234 4768 3240 4780
rect 3292 4768 3298 4820
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 7466 4808 7472 4820
rect 7064 4780 7472 4808
rect 7064 4768 7070 4780
rect 7466 4768 7472 4780
rect 7524 4808 7530 4820
rect 7561 4811 7619 4817
rect 7561 4808 7573 4811
rect 7524 4780 7573 4808
rect 7524 4768 7530 4780
rect 7561 4777 7573 4780
rect 7607 4777 7619 4811
rect 8110 4808 8116 4820
rect 8071 4780 8116 4808
rect 7561 4771 7619 4777
rect 8110 4768 8116 4780
rect 8168 4768 8174 4820
rect 10505 4811 10563 4817
rect 10505 4777 10517 4811
rect 10551 4808 10563 4811
rect 10686 4808 10692 4820
rect 10551 4780 10692 4808
rect 10551 4777 10563 4780
rect 10505 4771 10563 4777
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 11241 4811 11299 4817
rect 11241 4777 11253 4811
rect 11287 4808 11299 4811
rect 11330 4808 11336 4820
rect 11287 4780 11336 4808
rect 11287 4777 11299 4780
rect 11241 4771 11299 4777
rect 11330 4768 11336 4780
rect 11388 4808 11394 4820
rect 11425 4811 11483 4817
rect 11425 4808 11437 4811
rect 11388 4780 11437 4808
rect 11388 4768 11394 4780
rect 11425 4777 11437 4780
rect 11471 4777 11483 4811
rect 11790 4808 11796 4820
rect 11751 4780 11796 4808
rect 11425 4771 11483 4777
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 11882 4768 11888 4820
rect 11940 4808 11946 4820
rect 12989 4811 13047 4817
rect 12989 4808 13001 4811
rect 11940 4780 13001 4808
rect 11940 4768 11946 4780
rect 12989 4777 13001 4780
rect 13035 4777 13047 4811
rect 12989 4771 13047 4777
rect 13357 4811 13415 4817
rect 13357 4777 13369 4811
rect 13403 4808 13415 4811
rect 13446 4808 13452 4820
rect 13403 4780 13452 4808
rect 13403 4777 13415 4780
rect 13357 4771 13415 4777
rect 13446 4768 13452 4780
rect 13504 4808 13510 4820
rect 16114 4808 16120 4820
rect 13504 4780 16120 4808
rect 13504 4768 13510 4780
rect 16114 4768 16120 4780
rect 16172 4768 16178 4820
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 19613 4811 19671 4817
rect 19613 4808 19625 4811
rect 19392 4780 19625 4808
rect 19392 4768 19398 4780
rect 19613 4777 19625 4780
rect 19659 4777 19671 4811
rect 20530 4808 20536 4820
rect 20491 4780 20536 4808
rect 19613 4771 19671 4777
rect 20530 4768 20536 4780
rect 20588 4768 20594 4820
rect 10873 4743 10931 4749
rect 10873 4709 10885 4743
rect 10919 4740 10931 4743
rect 11514 4740 11520 4752
rect 10919 4712 11520 4740
rect 10919 4709 10931 4712
rect 10873 4703 10931 4709
rect 11514 4700 11520 4712
rect 11572 4700 11578 4752
rect 15378 4740 15384 4752
rect 11900 4712 15384 4740
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 2038 4672 2044 4684
rect 1443 4644 2044 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 2038 4632 2044 4644
rect 2096 4632 2102 4684
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4672 2559 4675
rect 2590 4672 2596 4684
rect 2547 4644 2596 4672
rect 2547 4641 2559 4644
rect 2501 4635 2559 4641
rect 2590 4632 2596 4644
rect 2648 4632 2654 4684
rect 4890 4681 4896 4684
rect 4884 4635 4896 4681
rect 4948 4672 4954 4684
rect 4948 4644 4984 4672
rect 4890 4632 4896 4635
rect 4948 4632 4954 4644
rect 7374 4632 7380 4684
rect 7432 4672 7438 4684
rect 7469 4675 7527 4681
rect 7469 4672 7481 4675
rect 7432 4644 7481 4672
rect 7432 4632 7438 4644
rect 7469 4641 7481 4644
rect 7515 4641 7527 4675
rect 7469 4635 7527 4641
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4604 2467 4607
rect 2682 4604 2688 4616
rect 2455 4576 2688 4604
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 4614 4604 4620 4616
rect 4575 4576 4620 4604
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 7190 4564 7196 4616
rect 7248 4604 7254 4616
rect 7745 4607 7803 4613
rect 7745 4604 7757 4607
rect 7248 4576 7757 4604
rect 7248 4564 7254 4576
rect 7745 4573 7757 4576
rect 7791 4604 7803 4607
rect 9490 4604 9496 4616
rect 7791 4576 9496 4604
rect 7791 4573 7803 4576
rect 7745 4567 7803 4573
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 11514 4564 11520 4616
rect 11572 4604 11578 4616
rect 11900 4613 11928 4712
rect 15378 4700 15384 4712
rect 15436 4700 15442 4752
rect 16476 4743 16534 4749
rect 16476 4709 16488 4743
rect 16522 4740 16534 4743
rect 17218 4740 17224 4752
rect 16522 4712 17224 4740
rect 16522 4709 16534 4712
rect 16476 4703 16534 4709
rect 17218 4700 17224 4712
rect 17276 4700 17282 4752
rect 13449 4675 13507 4681
rect 13449 4641 13461 4675
rect 13495 4672 13507 4675
rect 13538 4672 13544 4684
rect 13495 4644 13544 4672
rect 13495 4641 13507 4644
rect 13449 4635 13507 4641
rect 13538 4632 13544 4644
rect 13596 4632 13602 4684
rect 16206 4672 16212 4684
rect 16167 4644 16212 4672
rect 16206 4632 16212 4644
rect 16264 4632 16270 4684
rect 23566 4672 23572 4684
rect 23527 4644 23572 4672
rect 23566 4632 23572 4644
rect 23624 4632 23630 4684
rect 23842 4681 23848 4684
rect 23836 4672 23848 4681
rect 23803 4644 23848 4672
rect 23836 4635 23848 4644
rect 23842 4632 23848 4635
rect 23900 4632 23906 4684
rect 26510 4672 26516 4684
rect 26423 4644 26516 4672
rect 26510 4632 26516 4644
rect 26568 4672 26574 4684
rect 27154 4672 27160 4684
rect 26568 4644 27160 4672
rect 26568 4632 26574 4644
rect 27154 4632 27160 4644
rect 27212 4632 27218 4684
rect 11885 4607 11943 4613
rect 11885 4604 11897 4607
rect 11572 4576 11897 4604
rect 11572 4564 11578 4576
rect 11885 4573 11897 4576
rect 11931 4573 11943 4607
rect 12066 4604 12072 4616
rect 12027 4576 12072 4604
rect 11885 4567 11943 4573
rect 12066 4564 12072 4576
rect 12124 4564 12130 4616
rect 13630 4604 13636 4616
rect 13591 4576 13636 4604
rect 13630 4564 13636 4576
rect 13688 4564 13694 4616
rect 19702 4604 19708 4616
rect 19663 4576 19708 4604
rect 19702 4564 19708 4576
rect 19760 4564 19766 4616
rect 19886 4604 19892 4616
rect 19847 4576 19892 4604
rect 19886 4564 19892 4576
rect 19944 4564 19950 4616
rect 24946 4536 24952 4548
rect 24907 4508 24952 4536
rect 24946 4496 24952 4508
rect 25004 4496 25010 4548
rect 2685 4471 2743 4477
rect 2685 4437 2697 4471
rect 2731 4468 2743 4471
rect 2774 4468 2780 4480
rect 2731 4440 2780 4468
rect 2731 4437 2743 4440
rect 2685 4431 2743 4437
rect 2774 4428 2780 4440
rect 2832 4428 2838 4480
rect 5810 4428 5816 4480
rect 5868 4468 5874 4480
rect 5997 4471 6055 4477
rect 5997 4468 6009 4471
rect 5868 4440 6009 4468
rect 5868 4428 5874 4440
rect 5997 4437 6009 4440
rect 6043 4437 6055 4471
rect 7098 4468 7104 4480
rect 7059 4440 7104 4468
rect 5997 4431 6055 4437
rect 7098 4428 7104 4440
rect 7156 4428 7162 4480
rect 17586 4468 17592 4480
rect 17547 4440 17592 4468
rect 17586 4428 17592 4440
rect 17644 4428 17650 4480
rect 19242 4468 19248 4480
rect 19203 4440 19248 4468
rect 19242 4428 19248 4440
rect 19300 4428 19306 4480
rect 21358 4428 21364 4480
rect 21416 4468 21422 4480
rect 21634 4468 21640 4480
rect 21416 4440 21640 4468
rect 21416 4428 21422 4440
rect 21634 4428 21640 4440
rect 21692 4428 21698 4480
rect 26694 4468 26700 4480
rect 26655 4440 26700 4468
rect 26694 4428 26700 4440
rect 26752 4428 26758 4480
rect 1104 4378 28888 4400
rect 1104 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 15982 4378
rect 16034 4326 16046 4378
rect 16098 4326 16110 4378
rect 16162 4326 16174 4378
rect 16226 4326 25982 4378
rect 26034 4326 26046 4378
rect 26098 4326 26110 4378
rect 26162 4326 26174 4378
rect 26226 4326 28888 4378
rect 1104 4304 28888 4326
rect 2590 4264 2596 4276
rect 2551 4236 2596 4264
rect 2590 4224 2596 4236
rect 2648 4224 2654 4276
rect 4157 4267 4215 4273
rect 4157 4233 4169 4267
rect 4203 4264 4215 4267
rect 4338 4264 4344 4276
rect 4203 4236 4344 4264
rect 4203 4233 4215 4236
rect 4157 4227 4215 4233
rect 4338 4224 4344 4236
rect 4396 4264 4402 4276
rect 4801 4267 4859 4273
rect 4801 4264 4813 4267
rect 4396 4236 4813 4264
rect 4396 4224 4402 4236
rect 4801 4233 4813 4236
rect 4847 4264 4859 4267
rect 4890 4264 4896 4276
rect 4847 4236 4896 4264
rect 4847 4233 4859 4236
rect 4801 4227 4859 4233
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 7190 4264 7196 4276
rect 7151 4236 7196 4264
rect 7190 4224 7196 4236
rect 7248 4224 7254 4276
rect 7466 4264 7472 4276
rect 7427 4236 7472 4264
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 11514 4264 11520 4276
rect 11475 4236 11520 4264
rect 11514 4224 11520 4236
rect 11572 4224 11578 4276
rect 12066 4224 12072 4276
rect 12124 4264 12130 4276
rect 12161 4267 12219 4273
rect 12161 4264 12173 4267
rect 12124 4236 12173 4264
rect 12124 4224 12130 4236
rect 12161 4233 12173 4236
rect 12207 4233 12219 4267
rect 13446 4264 13452 4276
rect 13407 4236 13452 4264
rect 12161 4227 12219 4233
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 13630 4224 13636 4276
rect 13688 4264 13694 4276
rect 13725 4267 13783 4273
rect 13725 4264 13737 4267
rect 13688 4236 13737 4264
rect 13688 4224 13694 4236
rect 13725 4233 13737 4236
rect 13771 4233 13783 4267
rect 13725 4227 13783 4233
rect 17037 4267 17095 4273
rect 17037 4233 17049 4267
rect 17083 4264 17095 4267
rect 17218 4264 17224 4276
rect 17083 4236 17224 4264
rect 17083 4233 17095 4236
rect 17037 4227 17095 4233
rect 17218 4224 17224 4236
rect 17276 4224 17282 4276
rect 19337 4267 19395 4273
rect 19337 4233 19349 4267
rect 19383 4264 19395 4267
rect 19886 4264 19892 4276
rect 19383 4236 19892 4264
rect 19383 4233 19395 4236
rect 19337 4227 19395 4233
rect 19886 4224 19892 4236
rect 19944 4224 19950 4276
rect 21085 4267 21143 4273
rect 21085 4233 21097 4267
rect 21131 4264 21143 4267
rect 21266 4264 21272 4276
rect 21131 4236 21272 4264
rect 21131 4233 21143 4236
rect 21085 4227 21143 4233
rect 21266 4224 21272 4236
rect 21324 4224 21330 4276
rect 23566 4224 23572 4276
rect 23624 4264 23630 4276
rect 24213 4267 24271 4273
rect 24213 4264 24225 4267
rect 23624 4236 24225 4264
rect 23624 4224 23630 4236
rect 24213 4233 24225 4236
rect 24259 4233 24271 4267
rect 27154 4264 27160 4276
rect 27115 4236 27160 4264
rect 24213 4227 24271 4233
rect 27154 4224 27160 4236
rect 27212 4224 27218 4276
rect 4614 4156 4620 4208
rect 4672 4196 4678 4208
rect 5169 4199 5227 4205
rect 5169 4196 5181 4199
rect 4672 4168 5181 4196
rect 4672 4156 4678 4168
rect 5169 4165 5181 4168
rect 5215 4196 5227 4199
rect 5215 4168 7144 4196
rect 5215 4165 5227 4168
rect 5169 4159 5227 4165
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5276 4100 5917 4128
rect 5276 4072 5304 4100
rect 5905 4097 5917 4100
rect 5951 4128 5963 4131
rect 7006 4128 7012 4140
rect 5951 4100 7012 4128
rect 5951 4097 5963 4100
rect 5905 4091 5963 4097
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 7116 4128 7144 4168
rect 7374 4156 7380 4208
rect 7432 4196 7438 4208
rect 7837 4199 7895 4205
rect 7837 4196 7849 4199
rect 7432 4168 7849 4196
rect 7432 4156 7438 4168
rect 7837 4165 7849 4168
rect 7883 4165 7895 4199
rect 11790 4196 11796 4208
rect 11751 4168 11796 4196
rect 7837 4159 7895 4165
rect 11790 4156 11796 4168
rect 11848 4156 11854 4208
rect 13081 4199 13139 4205
rect 13081 4165 13093 4199
rect 13127 4196 13139 4199
rect 13538 4196 13544 4208
rect 13127 4168 13544 4196
rect 13127 4165 13139 4168
rect 13081 4159 13139 4165
rect 13538 4156 13544 4168
rect 13596 4156 13602 4208
rect 15841 4199 15899 4205
rect 15841 4165 15853 4199
rect 15887 4196 15899 4199
rect 19981 4199 20039 4205
rect 15887 4168 16519 4196
rect 15887 4165 15899 4168
rect 15841 4159 15899 4165
rect 16491 4140 16519 4168
rect 19981 4165 19993 4199
rect 20027 4165 20039 4199
rect 21284 4196 21312 4224
rect 21450 4196 21456 4208
rect 21284 4168 21456 4196
rect 19981 4159 20039 4165
rect 8110 4128 8116 4140
rect 7116 4100 8116 4128
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 16393 4131 16451 4137
rect 16393 4128 16405 4131
rect 15988 4100 16405 4128
rect 15988 4088 15994 4100
rect 16393 4097 16405 4100
rect 16439 4097 16451 4131
rect 16393 4091 16451 4097
rect 16482 4088 16488 4140
rect 16540 4128 16546 4140
rect 18969 4131 19027 4137
rect 16540 4100 16633 4128
rect 16540 4088 16546 4100
rect 18969 4097 18981 4131
rect 19015 4128 19027 4131
rect 19702 4128 19708 4140
rect 19015 4100 19708 4128
rect 19015 4097 19027 4100
rect 18969 4091 19027 4097
rect 19702 4088 19708 4100
rect 19760 4128 19766 4140
rect 19996 4128 20024 4159
rect 21450 4156 21456 4168
rect 21508 4196 21514 4208
rect 21508 4168 22140 4196
rect 21508 4156 21514 4168
rect 20622 4128 20628 4140
rect 19760 4100 20024 4128
rect 20583 4100 20628 4128
rect 19760 4088 19766 4100
rect 20622 4088 20628 4100
rect 20680 4088 20686 4140
rect 21358 4128 21364 4140
rect 21319 4100 21364 4128
rect 21358 4088 21364 4100
rect 21416 4088 21422 4140
rect 21634 4088 21640 4140
rect 21692 4128 21698 4140
rect 22112 4137 22140 4168
rect 22005 4131 22063 4137
rect 22005 4128 22017 4131
rect 21692 4100 22017 4128
rect 21692 4088 21698 4100
rect 22005 4097 22017 4100
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 22097 4131 22155 4137
rect 22097 4097 22109 4131
rect 22143 4097 22155 4131
rect 26789 4131 26847 4137
rect 26789 4128 26801 4131
rect 22097 4091 22155 4097
rect 26344 4100 26801 4128
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4029 1455 4063
rect 1397 4023 1455 4029
rect 1412 3992 1440 4023
rect 2682 4020 2688 4072
rect 2740 4060 2746 4072
rect 2777 4063 2835 4069
rect 2777 4060 2789 4063
rect 2740 4032 2789 4060
rect 2740 4020 2746 4032
rect 2777 4029 2789 4032
rect 2823 4029 2835 4063
rect 2777 4023 2835 4029
rect 2866 4020 2872 4072
rect 2924 4060 2930 4072
rect 3033 4063 3091 4069
rect 3033 4060 3045 4063
rect 2924 4032 3045 4060
rect 2924 4020 2930 4032
rect 3033 4029 3045 4032
rect 3079 4029 3091 4063
rect 3033 4023 3091 4029
rect 5258 4020 5264 4072
rect 5316 4060 5322 4072
rect 5316 4032 5409 4060
rect 5316 4020 5322 4032
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 19889 4063 19947 4069
rect 19889 4060 19901 4063
rect 19484 4032 19901 4060
rect 19484 4020 19490 4032
rect 19889 4029 19901 4032
rect 19935 4060 19947 4063
rect 20640 4060 20668 4088
rect 19935 4032 20668 4060
rect 21376 4060 21404 4088
rect 26344 4072 26372 4100
rect 26789 4097 26801 4100
rect 26835 4097 26847 4131
rect 26789 4091 26847 4097
rect 21913 4063 21971 4069
rect 21913 4060 21925 4063
rect 21376 4032 21925 4060
rect 19935 4029 19947 4032
rect 19889 4023 19947 4029
rect 21913 4029 21925 4032
rect 21959 4029 21971 4063
rect 23842 4060 23848 4072
rect 23803 4032 23848 4060
rect 21913 4023 21971 4029
rect 2038 3992 2044 4004
rect 1412 3964 2044 3992
rect 2038 3952 2044 3964
rect 2096 3952 2102 4004
rect 3970 3952 3976 4004
rect 4028 3992 4034 4004
rect 15473 3995 15531 4001
rect 4028 3964 5488 3992
rect 4028 3952 4034 3964
rect 1486 3884 1492 3936
rect 1544 3924 1550 3936
rect 5460 3933 5488 3964
rect 15473 3961 15485 3995
rect 15519 3992 15531 3995
rect 16298 3992 16304 4004
rect 15519 3964 16304 3992
rect 15519 3961 15531 3964
rect 15473 3955 15531 3961
rect 16298 3952 16304 3964
rect 16356 3952 16362 4004
rect 20346 3992 20352 4004
rect 20259 3964 20352 3992
rect 20346 3952 20352 3964
rect 20404 3992 20410 4004
rect 21928 3992 21956 4023
rect 23842 4020 23848 4032
rect 23900 4020 23906 4072
rect 26237 4063 26295 4069
rect 26237 4029 26249 4063
rect 26283 4060 26295 4063
rect 26326 4060 26332 4072
rect 26283 4032 26332 4060
rect 26283 4029 26295 4032
rect 26237 4023 26295 4029
rect 26326 4020 26332 4032
rect 26384 4020 26390 4072
rect 26602 4020 26608 4072
rect 26660 4060 26666 4072
rect 27341 4063 27399 4069
rect 27341 4060 27353 4063
rect 26660 4032 27353 4060
rect 26660 4020 26666 4032
rect 27341 4029 27353 4032
rect 27387 4060 27399 4063
rect 27893 4063 27951 4069
rect 27893 4060 27905 4063
rect 27387 4032 27905 4060
rect 27387 4029 27399 4032
rect 27341 4023 27399 4029
rect 27893 4029 27905 4032
rect 27939 4029 27951 4063
rect 27893 4023 27951 4029
rect 22002 3992 22008 4004
rect 20404 3964 21588 3992
rect 21928 3964 22008 3992
rect 20404 3952 20410 3964
rect 1581 3927 1639 3933
rect 1581 3924 1593 3927
rect 1544 3896 1593 3924
rect 1544 3884 1550 3896
rect 1581 3893 1593 3896
rect 1627 3893 1639 3927
rect 1581 3887 1639 3893
rect 5445 3927 5503 3933
rect 5445 3893 5457 3927
rect 5491 3893 5503 3927
rect 5445 3887 5503 3893
rect 15838 3884 15844 3936
rect 15896 3924 15902 3936
rect 15933 3927 15991 3933
rect 15933 3924 15945 3927
rect 15896 3896 15945 3924
rect 15896 3884 15902 3896
rect 15933 3893 15945 3896
rect 15979 3893 15991 3927
rect 15933 3887 15991 3893
rect 20438 3884 20444 3936
rect 20496 3924 20502 3936
rect 21560 3933 21588 3964
rect 22002 3952 22008 3964
rect 22060 3952 22066 4004
rect 21545 3927 21603 3933
rect 20496 3896 20541 3924
rect 20496 3884 20502 3896
rect 21545 3893 21557 3927
rect 21591 3893 21603 3927
rect 21545 3887 21603 3893
rect 26421 3927 26479 3933
rect 26421 3893 26433 3927
rect 26467 3924 26479 3927
rect 26694 3924 26700 3936
rect 26467 3896 26700 3924
rect 26467 3893 26479 3896
rect 26421 3887 26479 3893
rect 26694 3884 26700 3896
rect 26752 3884 26758 3936
rect 27522 3924 27528 3936
rect 27483 3896 27528 3924
rect 27522 3884 27528 3896
rect 27580 3884 27586 3936
rect 1104 3834 28888 3856
rect 1104 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 20982 3834
rect 21034 3782 21046 3834
rect 21098 3782 21110 3834
rect 21162 3782 21174 3834
rect 21226 3782 28888 3834
rect 1104 3760 28888 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 2866 3680 2872 3732
rect 2924 3720 2930 3732
rect 3053 3723 3111 3729
rect 3053 3720 3065 3723
rect 2924 3692 3065 3720
rect 2924 3680 2930 3692
rect 3053 3689 3065 3692
rect 3099 3689 3111 3723
rect 4338 3720 4344 3732
rect 4299 3692 4344 3720
rect 3053 3683 3111 3689
rect 4338 3680 4344 3692
rect 4396 3680 4402 3732
rect 5166 3680 5172 3732
rect 5224 3720 5230 3732
rect 5445 3723 5503 3729
rect 5445 3720 5457 3723
rect 5224 3692 5457 3720
rect 5224 3680 5230 3692
rect 5445 3689 5457 3692
rect 5491 3689 5503 3723
rect 5445 3683 5503 3689
rect 5626 3680 5632 3732
rect 5684 3720 5690 3732
rect 6181 3723 6239 3729
rect 6181 3720 6193 3723
rect 5684 3692 6193 3720
rect 5684 3680 5690 3692
rect 6181 3689 6193 3692
rect 6227 3720 6239 3723
rect 6822 3720 6828 3732
rect 6227 3692 6828 3720
rect 6227 3689 6239 3692
rect 6181 3683 6239 3689
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7377 3723 7435 3729
rect 7377 3689 7389 3723
rect 7423 3720 7435 3723
rect 7558 3720 7564 3732
rect 7423 3692 7564 3720
rect 7423 3689 7435 3692
rect 7377 3683 7435 3689
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 12066 3680 12072 3732
rect 12124 3720 12130 3732
rect 12161 3723 12219 3729
rect 12161 3720 12173 3723
rect 12124 3692 12173 3720
rect 12124 3680 12130 3692
rect 12161 3689 12173 3692
rect 12207 3689 12219 3723
rect 15930 3720 15936 3732
rect 15891 3692 15936 3720
rect 12161 3683 12219 3689
rect 15930 3680 15936 3692
rect 15988 3680 15994 3732
rect 19334 3720 19340 3732
rect 19295 3692 19340 3720
rect 19334 3680 19340 3692
rect 19392 3680 19398 3732
rect 20073 3723 20131 3729
rect 20073 3689 20085 3723
rect 20119 3720 20131 3723
rect 20438 3720 20444 3732
rect 20119 3692 20444 3720
rect 20119 3689 20131 3692
rect 20073 3683 20131 3689
rect 20438 3680 20444 3692
rect 20496 3720 20502 3732
rect 20901 3723 20959 3729
rect 20901 3720 20913 3723
rect 20496 3692 20913 3720
rect 20496 3680 20502 3692
rect 20901 3689 20913 3692
rect 20947 3689 20959 3723
rect 21269 3723 21327 3729
rect 21269 3720 21281 3723
rect 20901 3683 20959 3689
rect 21008 3692 21281 3720
rect 2682 3612 2688 3664
rect 2740 3652 2746 3664
rect 3513 3655 3571 3661
rect 3513 3652 3525 3655
rect 2740 3624 3525 3652
rect 2740 3612 2746 3624
rect 3513 3621 3525 3624
rect 3559 3652 3571 3655
rect 4614 3652 4620 3664
rect 3559 3624 4620 3652
rect 3559 3621 3571 3624
rect 3513 3615 3571 3621
rect 4614 3612 4620 3624
rect 4672 3612 4678 3664
rect 4982 3612 4988 3664
rect 5040 3652 5046 3664
rect 6457 3655 6515 3661
rect 6457 3652 6469 3655
rect 5040 3624 6469 3652
rect 5040 3612 5046 3624
rect 6457 3621 6469 3624
rect 6503 3621 6515 3655
rect 6457 3615 6515 3621
rect 15654 3612 15660 3664
rect 15712 3652 15718 3664
rect 16301 3655 16359 3661
rect 16301 3652 16313 3655
rect 15712 3624 16313 3652
rect 15712 3612 15718 3624
rect 16301 3621 16313 3624
rect 16347 3621 16359 3655
rect 16301 3615 16359 3621
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 2501 3587 2559 3593
rect 2501 3553 2513 3587
rect 2547 3584 2559 3587
rect 2590 3584 2596 3596
rect 2547 3556 2596 3584
rect 2547 3553 2559 3556
rect 2501 3547 2559 3553
rect 1412 3516 1440 3547
rect 2590 3544 2596 3556
rect 2648 3544 2654 3596
rect 6270 3584 6276 3596
rect 4816 3556 6276 3584
rect 2041 3519 2099 3525
rect 2041 3516 2053 3519
rect 1412 3488 2053 3516
rect 2041 3485 2053 3488
rect 2087 3516 2099 3519
rect 4816 3516 4844 3556
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 8018 3584 8024 3596
rect 7484 3556 8024 3584
rect 5537 3519 5595 3525
rect 5537 3516 5549 3519
rect 2087 3488 4844 3516
rect 4908 3488 5549 3516
rect 2087 3485 2099 3488
rect 2041 3479 2099 3485
rect 4908 3392 4936 3488
rect 5537 3485 5549 3488
rect 5583 3485 5595 3519
rect 5537 3479 5595 3485
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3516 5779 3519
rect 5810 3516 5816 3528
rect 5767 3488 5816 3516
rect 5767 3485 5779 3488
rect 5721 3479 5779 3485
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 6546 3476 6552 3528
rect 6604 3516 6610 3528
rect 7484 3525 7512 3556
rect 8018 3544 8024 3556
rect 8076 3544 8082 3596
rect 11054 3593 11060 3596
rect 11048 3584 11060 3593
rect 11015 3556 11060 3584
rect 11048 3547 11060 3556
rect 11054 3544 11060 3547
rect 11112 3544 11118 3596
rect 16316 3584 16344 3615
rect 16482 3612 16488 3664
rect 16540 3652 16546 3664
rect 17466 3655 17524 3661
rect 17466 3652 17478 3655
rect 16540 3624 17478 3652
rect 16540 3612 16546 3624
rect 17466 3621 17478 3624
rect 17512 3652 17524 3655
rect 17586 3652 17592 3664
rect 17512 3624 17592 3652
rect 17512 3621 17524 3624
rect 17466 3615 17524 3621
rect 17586 3612 17592 3624
rect 17644 3612 17650 3664
rect 20346 3652 20352 3664
rect 20307 3624 20352 3652
rect 20346 3612 20352 3624
rect 20404 3612 20410 3664
rect 20806 3612 20812 3664
rect 20864 3652 20870 3664
rect 21008 3652 21036 3692
rect 21269 3689 21281 3692
rect 21315 3720 21327 3723
rect 21818 3720 21824 3732
rect 21315 3692 21824 3720
rect 21315 3689 21327 3692
rect 21269 3683 21327 3689
rect 21818 3680 21824 3692
rect 21876 3680 21882 3732
rect 20864 3624 21036 3652
rect 21836 3652 21864 3680
rect 21836 3624 26556 3652
rect 20864 3612 20870 3624
rect 17221 3587 17279 3593
rect 17221 3584 17233 3587
rect 16316 3556 17233 3584
rect 17221 3553 17233 3556
rect 17267 3584 17279 3587
rect 17770 3584 17776 3596
rect 17267 3556 17776 3584
rect 17267 3553 17279 3556
rect 17221 3547 17279 3553
rect 17770 3544 17776 3556
rect 17828 3544 17834 3596
rect 25314 3584 25320 3596
rect 25275 3556 25320 3584
rect 25314 3544 25320 3556
rect 25372 3544 25378 3596
rect 26528 3593 26556 3624
rect 26513 3587 26571 3593
rect 26513 3553 26525 3587
rect 26559 3584 26571 3587
rect 27338 3584 27344 3596
rect 26559 3556 27344 3584
rect 26559 3553 26571 3556
rect 26513 3547 26571 3553
rect 27338 3544 27344 3556
rect 27396 3544 27402 3596
rect 7469 3519 7527 3525
rect 7469 3516 7481 3519
rect 6604 3488 7481 3516
rect 6604 3476 6610 3488
rect 7469 3485 7481 3488
rect 7515 3485 7527 3519
rect 7469 3479 7527 3485
rect 7561 3519 7619 3525
rect 7561 3485 7573 3519
rect 7607 3485 7619 3519
rect 7561 3479 7619 3485
rect 5828 3448 5856 3476
rect 7576 3448 7604 3479
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 10778 3516 10784 3528
rect 8812 3488 10784 3516
rect 8812 3476 8818 3488
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 21358 3516 21364 3528
rect 20772 3488 21364 3516
rect 20772 3476 20778 3488
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 21450 3476 21456 3528
rect 21508 3516 21514 3528
rect 21508 3488 21553 3516
rect 21508 3476 21514 3488
rect 25498 3448 25504 3460
rect 5828 3420 7604 3448
rect 25459 3420 25504 3448
rect 25498 3408 25504 3420
rect 25556 3408 25562 3460
rect 2682 3380 2688 3392
rect 2643 3352 2688 3380
rect 2682 3340 2688 3352
rect 2740 3340 2746 3392
rect 4890 3380 4896 3392
rect 4851 3352 4896 3380
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 5077 3383 5135 3389
rect 5077 3349 5089 3383
rect 5123 3380 5135 3383
rect 5442 3380 5448 3392
rect 5123 3352 5448 3380
rect 5123 3349 5135 3352
rect 5077 3343 5135 3349
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 6914 3380 6920 3392
rect 6875 3352 6920 3380
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 7009 3383 7067 3389
rect 7009 3349 7021 3383
rect 7055 3380 7067 3383
rect 7282 3380 7288 3392
rect 7055 3352 7288 3380
rect 7055 3349 7067 3352
rect 7009 3343 7067 3349
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 18598 3380 18604 3392
rect 18559 3352 18604 3380
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 26694 3380 26700 3392
rect 26655 3352 26700 3380
rect 26694 3340 26700 3352
rect 26752 3340 26758 3392
rect 1104 3290 28888 3312
rect 1104 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 15982 3290
rect 16034 3238 16046 3290
rect 16098 3238 16110 3290
rect 16162 3238 16174 3290
rect 16226 3238 25982 3290
rect 26034 3238 26046 3290
rect 26098 3238 26110 3290
rect 26162 3238 26174 3290
rect 26226 3238 28888 3290
rect 1104 3216 28888 3238
rect 2590 3176 2596 3188
rect 2551 3148 2596 3176
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 3881 3179 3939 3185
rect 3881 3145 3893 3179
rect 3927 3176 3939 3179
rect 4890 3176 4896 3188
rect 3927 3148 4896 3176
rect 3927 3145 3939 3148
rect 3881 3139 3939 3145
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 5166 3176 5172 3188
rect 5127 3148 5172 3176
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 7392 3148 10609 3176
rect 2608 3108 2636 3136
rect 6546 3108 6552 3120
rect 2608 3080 6552 3108
rect 6546 3068 6552 3080
rect 6604 3068 6610 3120
rect 1670 3000 1676 3052
rect 1728 3000 1734 3052
rect 4338 3000 4344 3052
rect 4396 3040 4402 3052
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 4396 3012 4445 3040
rect 4396 3000 4402 3012
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 5258 3040 5264 3052
rect 4433 3003 4491 3009
rect 4908 3012 5264 3040
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 1688 2972 1716 3000
rect 1854 2972 1860 2984
rect 1443 2944 1860 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 1854 2932 1860 2944
rect 1912 2932 1918 2984
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 2498 2972 2504 2984
rect 2271 2944 2504 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 2498 2932 2504 2944
rect 2556 2972 2562 2984
rect 2685 2975 2743 2981
rect 2685 2972 2697 2975
rect 2556 2944 2697 2972
rect 2556 2932 2562 2944
rect 2685 2941 2697 2944
rect 2731 2941 2743 2975
rect 2685 2935 2743 2941
rect 3421 2975 3479 2981
rect 3421 2941 3433 2975
rect 3467 2972 3479 2975
rect 4249 2975 4307 2981
rect 4249 2972 4261 2975
rect 3467 2944 4261 2972
rect 3467 2941 3479 2944
rect 3421 2935 3479 2941
rect 4249 2941 4261 2944
rect 4295 2972 4307 2975
rect 4908 2972 4936 3012
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 7392 3049 7420 3148
rect 10597 3145 10609 3148
rect 10643 3176 10655 3179
rect 11054 3176 11060 3188
rect 10643 3148 11060 3176
rect 10643 3145 10655 3148
rect 10597 3139 10655 3145
rect 11054 3136 11060 3148
rect 11112 3176 11118 3188
rect 11149 3179 11207 3185
rect 11149 3176 11161 3179
rect 11112 3148 11161 3176
rect 11112 3136 11118 3148
rect 11149 3145 11161 3148
rect 11195 3145 11207 3179
rect 13170 3176 13176 3188
rect 13131 3148 13176 3176
rect 11149 3139 11207 3145
rect 13170 3136 13176 3148
rect 13228 3136 13234 3188
rect 15197 3179 15255 3185
rect 15197 3145 15209 3179
rect 15243 3176 15255 3179
rect 15838 3176 15844 3188
rect 15243 3148 15844 3176
rect 15243 3145 15255 3148
rect 15197 3139 15255 3145
rect 7558 3068 7564 3120
rect 7616 3108 7622 3120
rect 7837 3111 7895 3117
rect 7837 3108 7849 3111
rect 7616 3080 7849 3108
rect 7616 3068 7622 3080
rect 7837 3077 7849 3080
rect 7883 3077 7895 3111
rect 7837 3071 7895 3077
rect 10778 3068 10784 3120
rect 10836 3108 10842 3120
rect 11517 3111 11575 3117
rect 11517 3108 11529 3111
rect 10836 3080 11529 3108
rect 10836 3068 10842 3080
rect 11517 3077 11529 3080
rect 11563 3077 11575 3111
rect 11517 3071 11575 3077
rect 7377 3043 7435 3049
rect 7377 3040 7389 3043
rect 6972 3012 7389 3040
rect 6972 3000 6978 3012
rect 7377 3009 7389 3012
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3040 9183 3043
rect 9171 3012 9352 3040
rect 9171 3009 9183 3012
rect 9125 3003 9183 3009
rect 4295 2944 4936 2972
rect 4295 2941 4307 2944
rect 4249 2935 4307 2941
rect 4982 2932 4988 2984
rect 5040 2972 5046 2984
rect 5445 2975 5503 2981
rect 5445 2972 5457 2975
rect 5040 2944 5457 2972
rect 5040 2932 5046 2944
rect 5445 2941 5457 2944
rect 5491 2941 5503 2975
rect 5718 2972 5724 2984
rect 5679 2944 5724 2972
rect 5445 2935 5503 2941
rect 5718 2932 5724 2944
rect 5776 2932 5782 2984
rect 7098 2932 7104 2984
rect 7156 2972 7162 2984
rect 7193 2975 7251 2981
rect 7193 2972 7205 2975
rect 7156 2944 7205 2972
rect 7156 2932 7162 2944
rect 7193 2941 7205 2944
rect 7239 2972 7251 2975
rect 8573 2975 8631 2981
rect 8573 2972 8585 2975
rect 7239 2944 8585 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 8573 2941 8585 2944
rect 8619 2941 8631 2975
rect 8573 2935 8631 2941
rect 8754 2932 8760 2984
rect 8812 2972 8818 2984
rect 9217 2975 9275 2981
rect 9217 2972 9229 2975
rect 8812 2944 9229 2972
rect 8812 2932 8818 2944
rect 9217 2941 9229 2944
rect 9263 2941 9275 2975
rect 9324 2972 9352 3012
rect 9490 2981 9496 2984
rect 9484 2972 9496 2981
rect 9324 2944 9496 2972
rect 9217 2935 9275 2941
rect 9484 2935 9496 2944
rect 9490 2932 9496 2935
rect 9548 2932 9554 2984
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 13170 2972 13176 2984
rect 12483 2944 13176 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 13170 2932 13176 2944
rect 13228 2932 13234 2984
rect 14369 2975 14427 2981
rect 14369 2941 14381 2975
rect 14415 2972 14427 2975
rect 15212 2972 15240 3139
rect 15838 3136 15844 3148
rect 15896 3136 15902 3188
rect 16577 3179 16635 3185
rect 16577 3145 16589 3179
rect 16623 3176 16635 3179
rect 16666 3176 16672 3188
rect 16623 3148 16672 3176
rect 16623 3145 16635 3148
rect 16577 3139 16635 3145
rect 16666 3136 16672 3148
rect 16724 3136 16730 3188
rect 17497 3179 17555 3185
rect 17497 3145 17509 3179
rect 17543 3176 17555 3179
rect 17586 3176 17592 3188
rect 17543 3148 17592 3176
rect 17543 3145 17555 3148
rect 17497 3139 17555 3145
rect 17586 3136 17592 3148
rect 17644 3136 17650 3188
rect 17770 3176 17776 3188
rect 17731 3148 17776 3176
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 21358 3136 21364 3188
rect 21416 3176 21422 3188
rect 22097 3179 22155 3185
rect 22097 3176 22109 3179
rect 21416 3148 22109 3176
rect 21416 3136 21422 3148
rect 22097 3145 22109 3148
rect 22143 3145 22155 3179
rect 22097 3139 22155 3145
rect 24305 3179 24363 3185
rect 24305 3145 24317 3179
rect 24351 3176 24363 3179
rect 24673 3179 24731 3185
rect 24673 3176 24685 3179
rect 24351 3148 24685 3176
rect 24351 3145 24363 3148
rect 24305 3139 24363 3145
rect 24673 3145 24685 3148
rect 24719 3176 24731 3179
rect 25406 3176 25412 3188
rect 24719 3148 25412 3176
rect 24719 3145 24731 3148
rect 24673 3139 24731 3145
rect 21450 3068 21456 3120
rect 21508 3108 21514 3120
rect 21545 3111 21603 3117
rect 21545 3108 21557 3111
rect 21508 3080 21557 3108
rect 21508 3068 21514 3080
rect 21545 3077 21557 3080
rect 21591 3077 21603 3111
rect 21545 3071 21603 3077
rect 18598 3000 18604 3052
rect 18656 3040 18662 3052
rect 19981 3043 20039 3049
rect 19981 3040 19993 3043
rect 18656 3012 19993 3040
rect 18656 3000 18662 3012
rect 19981 3009 19993 3012
rect 20027 3040 20039 3043
rect 20070 3040 20076 3052
rect 20027 3012 20076 3040
rect 20027 3009 20039 3012
rect 19981 3003 20039 3009
rect 20070 3000 20076 3012
rect 20128 3040 20134 3052
rect 20128 3012 20300 3040
rect 20128 3000 20134 3012
rect 16666 2972 16672 2984
rect 14415 2944 15240 2972
rect 16627 2944 16672 2972
rect 14415 2941 14427 2944
rect 14369 2935 14427 2941
rect 16666 2932 16672 2944
rect 16724 2932 16730 2984
rect 16945 2975 17003 2981
rect 16945 2941 16957 2975
rect 16991 2972 17003 2975
rect 17770 2972 17776 2984
rect 16991 2944 17776 2972
rect 16991 2941 17003 2944
rect 16945 2935 17003 2941
rect 17770 2932 17776 2944
rect 17828 2932 17834 2984
rect 18874 2972 18880 2984
rect 18787 2944 18880 2972
rect 18874 2932 18880 2944
rect 18932 2972 18938 2984
rect 19613 2975 19671 2981
rect 19613 2972 19625 2975
rect 18932 2944 19625 2972
rect 18932 2932 18938 2944
rect 19613 2941 19625 2944
rect 19659 2941 19671 2975
rect 20162 2972 20168 2984
rect 20123 2944 20168 2972
rect 19613 2935 19671 2941
rect 20162 2932 20168 2944
rect 20220 2932 20226 2984
rect 20272 2972 20300 3012
rect 24780 2981 24808 3148
rect 25406 3136 25412 3148
rect 25464 3136 25470 3188
rect 27338 3176 27344 3188
rect 27299 3148 27344 3176
rect 27338 3136 27344 3148
rect 27396 3136 27402 3188
rect 24949 3111 25007 3117
rect 24949 3077 24961 3111
rect 24995 3108 25007 3111
rect 26326 3108 26332 3120
rect 24995 3080 26332 3108
rect 24995 3077 25007 3080
rect 24949 3071 25007 3077
rect 26326 3068 26332 3080
rect 26384 3068 26390 3120
rect 25314 3040 25320 3052
rect 25275 3012 25320 3040
rect 25314 3000 25320 3012
rect 25372 3000 25378 3052
rect 20421 2975 20479 2981
rect 20421 2972 20433 2975
rect 20272 2944 20433 2972
rect 20421 2941 20433 2944
rect 20467 2941 20479 2975
rect 20421 2935 20479 2941
rect 23661 2975 23719 2981
rect 23661 2941 23673 2975
rect 23707 2972 23719 2975
rect 24765 2975 24823 2981
rect 24765 2972 24777 2975
rect 23707 2944 24777 2972
rect 23707 2941 23719 2944
rect 23661 2935 23719 2941
rect 24765 2941 24777 2944
rect 24811 2941 24823 2975
rect 26418 2972 26424 2984
rect 26379 2944 26424 2972
rect 24765 2935 24823 2941
rect 26418 2932 26424 2944
rect 26476 2972 26482 2984
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26476 2944 26985 2972
rect 26476 2932 26482 2944
rect 26973 2941 26985 2944
rect 27019 2941 27031 2975
rect 26973 2935 27031 2941
rect 27430 2932 27436 2984
rect 27488 2972 27494 2984
rect 27525 2975 27583 2981
rect 27525 2972 27537 2975
rect 27488 2944 27537 2972
rect 27488 2932 27494 2944
rect 27525 2941 27537 2944
rect 27571 2972 27583 2975
rect 28077 2975 28135 2981
rect 28077 2972 28089 2975
rect 27571 2944 28089 2972
rect 27571 2941 27583 2944
rect 27525 2935 27583 2941
rect 28077 2941 28089 2944
rect 28123 2941 28135 2975
rect 28077 2935 28135 2941
rect 1673 2907 1731 2913
rect 1673 2873 1685 2907
rect 1719 2904 1731 2907
rect 2038 2904 2044 2916
rect 1719 2876 2044 2904
rect 1719 2873 1731 2876
rect 1673 2867 1731 2873
rect 2038 2864 2044 2876
rect 2096 2864 2102 2916
rect 3789 2907 3847 2913
rect 3789 2873 3801 2907
rect 3835 2904 3847 2907
rect 4341 2907 4399 2913
rect 4341 2904 4353 2907
rect 3835 2876 4353 2904
rect 3835 2873 3847 2876
rect 3789 2867 3847 2873
rect 4341 2873 4353 2876
rect 4387 2904 4399 2907
rect 5534 2904 5540 2916
rect 4387 2876 5540 2904
rect 4387 2873 4399 2876
rect 4341 2867 4399 2873
rect 5534 2864 5540 2876
rect 5592 2864 5598 2916
rect 6914 2864 6920 2916
rect 6972 2904 6978 2916
rect 7285 2907 7343 2913
rect 7285 2904 7297 2907
rect 6972 2876 7297 2904
rect 6972 2864 6978 2876
rect 7285 2873 7297 2876
rect 7331 2904 7343 2907
rect 8205 2907 8263 2913
rect 8205 2904 8217 2907
rect 7331 2876 8217 2904
rect 7331 2873 7343 2876
rect 7285 2867 7343 2873
rect 8205 2873 8217 2876
rect 8251 2873 8263 2907
rect 8205 2867 8263 2873
rect 12066 2864 12072 2916
rect 12124 2904 12130 2916
rect 12713 2907 12771 2913
rect 12713 2904 12725 2907
rect 12124 2876 12725 2904
rect 12124 2864 12130 2876
rect 12713 2873 12725 2876
rect 12759 2873 12771 2907
rect 12713 2867 12771 2873
rect 14645 2907 14703 2913
rect 14645 2873 14657 2907
rect 14691 2904 14703 2907
rect 14918 2904 14924 2916
rect 14691 2876 14924 2904
rect 14691 2873 14703 2876
rect 14645 2867 14703 2873
rect 14918 2864 14924 2876
rect 14976 2864 14982 2916
rect 19150 2904 19156 2916
rect 19111 2876 19156 2904
rect 19150 2864 19156 2876
rect 19208 2864 19214 2916
rect 2866 2836 2872 2848
rect 2827 2808 2872 2836
rect 2866 2796 2872 2808
rect 2924 2796 2930 2848
rect 5166 2796 5172 2848
rect 5224 2836 5230 2848
rect 5810 2836 5816 2848
rect 5224 2808 5816 2836
rect 5224 2796 5230 2808
rect 5810 2796 5816 2808
rect 5868 2836 5874 2848
rect 6181 2839 6239 2845
rect 6181 2836 6193 2839
rect 5868 2808 6193 2836
rect 5868 2796 5874 2808
rect 6181 2805 6193 2808
rect 6227 2805 6239 2839
rect 6822 2836 6828 2848
rect 6783 2808 6828 2836
rect 6181 2799 6239 2805
rect 6822 2796 6828 2808
rect 6880 2796 6886 2848
rect 23842 2836 23848 2848
rect 23803 2808 23848 2836
rect 23842 2796 23848 2808
rect 23900 2796 23906 2848
rect 26602 2836 26608 2848
rect 26563 2808 26608 2836
rect 26602 2796 26608 2808
rect 26660 2796 26666 2848
rect 27706 2836 27712 2848
rect 27667 2808 27712 2836
rect 27706 2796 27712 2808
rect 27764 2796 27770 2848
rect 1104 2746 28888 2768
rect 1104 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 20982 2746
rect 21034 2694 21046 2746
rect 21098 2694 21110 2746
rect 21162 2694 21174 2746
rect 21226 2694 28888 2746
rect 1104 2672 28888 2694
rect 1854 2592 1860 2644
rect 1912 2632 1918 2644
rect 2317 2635 2375 2641
rect 2317 2632 2329 2635
rect 1912 2604 2329 2632
rect 1912 2592 1918 2604
rect 2317 2601 2329 2604
rect 2363 2601 2375 2635
rect 5166 2632 5172 2644
rect 5127 2604 5172 2632
rect 2317 2595 2375 2601
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 5442 2592 5448 2644
rect 5500 2632 5506 2644
rect 6273 2635 6331 2641
rect 6273 2632 6285 2635
rect 5500 2604 6285 2632
rect 5500 2592 5506 2604
rect 6273 2601 6285 2604
rect 6319 2632 6331 2635
rect 6549 2635 6607 2641
rect 6549 2632 6561 2635
rect 6319 2604 6561 2632
rect 6319 2601 6331 2604
rect 6273 2595 6331 2601
rect 6549 2601 6561 2604
rect 6595 2601 6607 2635
rect 6914 2632 6920 2644
rect 6875 2604 6920 2632
rect 6549 2595 6607 2601
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 8754 2592 8760 2644
rect 8812 2632 8818 2644
rect 9217 2635 9275 2641
rect 9217 2632 9229 2635
rect 8812 2604 9229 2632
rect 8812 2592 8818 2604
rect 9217 2601 9229 2604
rect 9263 2601 9275 2635
rect 9217 2595 9275 2601
rect 13633 2635 13691 2641
rect 13633 2601 13645 2635
rect 13679 2632 13691 2635
rect 13722 2632 13728 2644
rect 13679 2604 13728 2632
rect 13679 2601 13691 2604
rect 13633 2595 13691 2601
rect 5813 2567 5871 2573
rect 5813 2533 5825 2567
rect 5859 2564 5871 2567
rect 7742 2564 7748 2576
rect 5859 2536 7748 2564
rect 5859 2533 5871 2536
rect 5813 2527 5871 2533
rect 7742 2524 7748 2536
rect 7800 2524 7806 2576
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 1949 2499 2007 2505
rect 1949 2496 1961 2499
rect 1443 2468 1961 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 1949 2465 1961 2468
rect 1995 2496 2007 2499
rect 2222 2496 2228 2508
rect 1995 2468 2228 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 2222 2456 2228 2468
rect 2280 2456 2286 2508
rect 2501 2499 2559 2505
rect 2501 2465 2513 2499
rect 2547 2496 2559 2499
rect 3142 2496 3148 2508
rect 2547 2468 3148 2496
rect 2547 2465 2559 2468
rect 2501 2459 2559 2465
rect 3142 2456 3148 2468
rect 3200 2496 3206 2508
rect 3237 2499 3295 2505
rect 3237 2496 3249 2499
rect 3200 2468 3249 2496
rect 3200 2456 3206 2468
rect 3237 2465 3249 2468
rect 3283 2465 3295 2499
rect 3237 2459 3295 2465
rect 3881 2499 3939 2505
rect 3881 2465 3893 2499
rect 3927 2496 3939 2499
rect 4062 2496 4068 2508
rect 3927 2468 4068 2496
rect 3927 2465 3939 2468
rect 3881 2459 3939 2465
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 5537 2499 5595 2505
rect 5537 2465 5549 2499
rect 5583 2496 5595 2499
rect 5626 2496 5632 2508
rect 5583 2468 5632 2496
rect 5583 2465 5595 2468
rect 5537 2459 5595 2465
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 7282 2496 7288 2508
rect 7195 2468 7288 2496
rect 7282 2456 7288 2468
rect 7340 2496 7346 2508
rect 7929 2499 7987 2505
rect 7929 2496 7941 2499
rect 7340 2468 7941 2496
rect 7340 2456 7346 2468
rect 7929 2465 7941 2468
rect 7975 2465 7987 2499
rect 7929 2459 7987 2465
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9732 2468 9781 2496
rect 9732 2456 9738 2468
rect 9769 2465 9781 2468
rect 9815 2496 9827 2499
rect 10505 2499 10563 2505
rect 10505 2496 10517 2499
rect 9815 2468 10517 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 10505 2465 10517 2468
rect 10551 2465 10563 2499
rect 11054 2496 11060 2508
rect 11015 2468 11060 2496
rect 10505 2459 10563 2465
rect 11054 2456 11060 2468
rect 11112 2496 11118 2508
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 11112 2468 11805 2496
rect 11112 2456 11118 2468
rect 11793 2465 11805 2468
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 12805 2499 12863 2505
rect 12805 2465 12817 2499
rect 12851 2496 12863 2499
rect 13648 2496 13676 2595
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 16390 2632 16396 2644
rect 16351 2604 16396 2632
rect 16390 2592 16396 2604
rect 16448 2592 16454 2644
rect 18598 2632 18604 2644
rect 18559 2604 18604 2632
rect 18598 2592 18604 2604
rect 18656 2592 18662 2644
rect 19429 2635 19487 2641
rect 19429 2601 19441 2635
rect 19475 2632 19487 2635
rect 19978 2632 19984 2644
rect 19475 2604 19984 2632
rect 19475 2601 19487 2604
rect 19429 2595 19487 2601
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 20162 2592 20168 2644
rect 20220 2632 20226 2644
rect 20533 2635 20591 2641
rect 20533 2632 20545 2635
rect 20220 2604 20545 2632
rect 20220 2592 20226 2604
rect 20533 2601 20545 2604
rect 20579 2601 20591 2635
rect 20533 2595 20591 2601
rect 20806 2592 20812 2644
rect 20864 2632 20870 2644
rect 20901 2635 20959 2641
rect 20901 2632 20913 2635
rect 20864 2604 20913 2632
rect 20864 2592 20870 2604
rect 20901 2601 20913 2604
rect 20947 2601 20959 2635
rect 20901 2595 20959 2601
rect 21266 2592 21272 2644
rect 21324 2632 21330 2644
rect 21361 2635 21419 2641
rect 21361 2632 21373 2635
rect 21324 2604 21373 2632
rect 21324 2592 21330 2604
rect 21361 2601 21373 2604
rect 21407 2601 21419 2635
rect 21361 2595 21419 2601
rect 12851 2468 13676 2496
rect 15657 2499 15715 2505
rect 12851 2465 12863 2468
rect 12805 2459 12863 2465
rect 15657 2465 15669 2499
rect 15703 2496 15715 2499
rect 16408 2496 16436 2592
rect 18230 2524 18236 2576
rect 18288 2564 18294 2576
rect 18969 2567 19027 2573
rect 18969 2564 18981 2567
rect 18288 2536 18981 2564
rect 18288 2524 18294 2536
rect 18969 2533 18981 2536
rect 19015 2564 19027 2567
rect 19889 2567 19947 2573
rect 19889 2564 19901 2567
rect 19015 2536 19901 2564
rect 19015 2533 19027 2536
rect 18969 2527 19027 2533
rect 19889 2533 19901 2536
rect 19935 2533 19947 2567
rect 19889 2527 19947 2533
rect 24670 2524 24676 2576
rect 24728 2564 24734 2576
rect 24728 2536 25728 2564
rect 24728 2524 24734 2536
rect 15703 2468 16436 2496
rect 16945 2499 17003 2505
rect 15703 2465 15715 2468
rect 15657 2459 15715 2465
rect 16945 2465 16957 2499
rect 16991 2496 17003 2499
rect 17773 2499 17831 2505
rect 17773 2496 17785 2499
rect 16991 2468 17785 2496
rect 16991 2465 17003 2468
rect 16945 2459 17003 2465
rect 17773 2465 17785 2468
rect 17819 2496 17831 2499
rect 17862 2496 17868 2508
rect 17819 2468 17868 2496
rect 17819 2465 17831 2468
rect 17773 2459 17831 2465
rect 17862 2456 17868 2468
rect 17920 2456 17926 2508
rect 22278 2496 22284 2508
rect 22239 2468 22284 2496
rect 22278 2456 22284 2468
rect 22336 2496 22342 2508
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22336 2468 23029 2496
rect 22336 2456 22342 2468
rect 23017 2465 23029 2468
rect 23063 2465 23075 2499
rect 24026 2496 24032 2508
rect 23987 2468 24032 2496
rect 23017 2459 23075 2465
rect 24026 2456 24032 2468
rect 24084 2496 24090 2508
rect 25700 2505 25728 2536
rect 24765 2499 24823 2505
rect 24765 2496 24777 2499
rect 24084 2468 24777 2496
rect 24084 2456 24090 2468
rect 24765 2465 24777 2468
rect 24811 2465 24823 2499
rect 24765 2459 24823 2465
rect 25685 2499 25743 2505
rect 25685 2465 25697 2499
rect 25731 2496 25743 2499
rect 26237 2499 26295 2505
rect 26237 2496 26249 2499
rect 25731 2468 26249 2496
rect 25731 2465 25743 2468
rect 25685 2459 25743 2465
rect 26237 2465 26249 2468
rect 26283 2465 26295 2499
rect 26237 2459 26295 2465
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2428 2835 2431
rect 3510 2428 3516 2440
rect 2823 2400 3516 2428
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 4890 2428 4896 2440
rect 4387 2400 4896 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2428 6607 2431
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 6595 2400 7389 2428
rect 6595 2397 6607 2400
rect 6549 2391 6607 2397
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2397 7527 2431
rect 9950 2428 9956 2440
rect 9911 2400 9956 2428
rect 7469 2391 7527 2397
rect 6733 2363 6791 2369
rect 6733 2329 6745 2363
rect 6779 2360 6791 2363
rect 7190 2360 7196 2372
rect 6779 2332 7196 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 7190 2320 7196 2332
rect 7248 2360 7254 2372
rect 7484 2360 7512 2391
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 10594 2388 10600 2440
rect 10652 2428 10658 2440
rect 11241 2431 11299 2437
rect 11241 2428 11253 2431
rect 10652 2400 11253 2428
rect 10652 2388 10658 2400
rect 11241 2397 11253 2400
rect 11287 2397 11299 2431
rect 11241 2391 11299 2397
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2428 13139 2431
rect 13446 2428 13452 2440
rect 13127 2400 13452 2428
rect 13127 2397 13139 2400
rect 13081 2391 13139 2397
rect 13446 2388 13452 2400
rect 13504 2388 13510 2440
rect 15933 2431 15991 2437
rect 15933 2397 15945 2431
rect 15979 2428 15991 2431
rect 16298 2428 16304 2440
rect 15979 2400 16304 2428
rect 15979 2397 15991 2400
rect 15933 2391 15991 2397
rect 16298 2388 16304 2400
rect 16356 2388 16362 2440
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2428 17279 2431
rect 19150 2428 19156 2440
rect 17267 2400 19156 2428
rect 17267 2397 17279 2400
rect 17221 2391 17279 2397
rect 19150 2388 19156 2400
rect 19208 2388 19214 2440
rect 20070 2428 20076 2440
rect 20031 2400 20076 2428
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 22557 2431 22615 2437
rect 22557 2397 22569 2431
rect 22603 2428 22615 2431
rect 23474 2428 23480 2440
rect 22603 2400 23480 2428
rect 22603 2397 22615 2400
rect 22557 2391 22615 2397
rect 23474 2388 23480 2400
rect 23532 2388 23538 2440
rect 24210 2428 24216 2440
rect 24171 2400 24216 2428
rect 24210 2388 24216 2400
rect 24268 2388 24274 2440
rect 7248 2332 7512 2360
rect 19521 2363 19579 2369
rect 7248 2320 7254 2332
rect 19521 2329 19533 2363
rect 19567 2360 19579 2363
rect 20530 2360 20536 2372
rect 19567 2332 20536 2360
rect 19567 2329 19579 2332
rect 19521 2323 19579 2329
rect 20530 2320 20536 2332
rect 20588 2320 20594 2372
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 25866 2292 25872 2304
rect 25827 2264 25872 2292
rect 25866 2252 25872 2264
rect 25924 2252 25930 2304
rect 27065 2295 27123 2301
rect 27065 2261 27077 2295
rect 27111 2292 27123 2295
rect 29178 2292 29184 2304
rect 27111 2264 29184 2292
rect 27111 2261 27123 2264
rect 27065 2255 27123 2261
rect 29178 2252 29184 2264
rect 29236 2252 29242 2304
rect 1104 2202 28888 2224
rect 1104 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 15982 2202
rect 16034 2150 16046 2202
rect 16098 2150 16110 2202
rect 16162 2150 16174 2202
rect 16226 2150 25982 2202
rect 26034 2150 26046 2202
rect 26098 2150 26110 2202
rect 26162 2150 26174 2202
rect 26226 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 3332 22108 3384 22160
rect 12072 22108 12124 22160
rect 21824 22108 21876 22160
rect 24860 22108 24912 22160
rect 1676 22040 1728 22092
rect 2136 22040 2188 22092
rect 5982 21734 6034 21786
rect 6046 21734 6098 21786
rect 6110 21734 6162 21786
rect 6174 21734 6226 21786
rect 15982 21734 16034 21786
rect 16046 21734 16098 21786
rect 16110 21734 16162 21786
rect 16174 21734 16226 21786
rect 25982 21734 26034 21786
rect 26046 21734 26098 21786
rect 26110 21734 26162 21786
rect 26174 21734 26226 21786
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 20982 21190 21034 21242
rect 21046 21190 21098 21242
rect 21110 21190 21162 21242
rect 21174 21190 21226 21242
rect 3976 21088 4028 21140
rect 7288 21088 7340 21140
rect 17040 20927 17092 20936
rect 17040 20893 17049 20927
rect 17049 20893 17083 20927
rect 17083 20893 17092 20927
rect 17040 20884 17092 20893
rect 4068 20748 4120 20800
rect 7564 20748 7616 20800
rect 8392 20791 8444 20800
rect 8392 20757 8401 20791
rect 8401 20757 8435 20791
rect 8435 20757 8444 20791
rect 8392 20748 8444 20757
rect 13544 20791 13596 20800
rect 13544 20757 13553 20791
rect 13553 20757 13587 20791
rect 13587 20757 13596 20791
rect 13544 20748 13596 20757
rect 23664 20791 23716 20800
rect 23664 20757 23673 20791
rect 23673 20757 23707 20791
rect 23707 20757 23716 20791
rect 23664 20748 23716 20757
rect 5982 20646 6034 20698
rect 6046 20646 6098 20698
rect 6110 20646 6162 20698
rect 6174 20646 6226 20698
rect 15982 20646 16034 20698
rect 16046 20646 16098 20698
rect 16110 20646 16162 20698
rect 16174 20646 16226 20698
rect 25982 20646 26034 20698
rect 26046 20646 26098 20698
rect 26110 20646 26162 20698
rect 26174 20646 26226 20698
rect 8208 20544 8260 20596
rect 21640 20544 21692 20596
rect 20628 20519 20680 20528
rect 20628 20485 20637 20519
rect 20637 20485 20671 20519
rect 20671 20485 20680 20519
rect 20628 20476 20680 20485
rect 18328 20408 18380 20460
rect 3516 20383 3568 20392
rect 3516 20349 3525 20383
rect 3525 20349 3559 20383
rect 3559 20349 3568 20383
rect 3516 20340 3568 20349
rect 8392 20340 8444 20392
rect 12440 20340 12492 20392
rect 13544 20383 13596 20392
rect 13544 20349 13553 20383
rect 13553 20349 13587 20383
rect 13587 20349 13596 20383
rect 13544 20340 13596 20349
rect 16672 20383 16724 20392
rect 16672 20349 16681 20383
rect 16681 20349 16715 20383
rect 16715 20349 16724 20383
rect 16672 20340 16724 20349
rect 19248 20383 19300 20392
rect 19248 20349 19257 20383
rect 19257 20349 19291 20383
rect 19291 20349 19300 20383
rect 19248 20340 19300 20349
rect 23664 20383 23716 20392
rect 23664 20349 23673 20383
rect 23673 20349 23707 20383
rect 23707 20349 23716 20383
rect 23664 20340 23716 20349
rect 4068 20272 4120 20324
rect 4896 20247 4948 20256
rect 4896 20213 4905 20247
rect 4905 20213 4939 20247
rect 4939 20213 4948 20247
rect 4896 20204 4948 20213
rect 7840 20204 7892 20256
rect 20720 20272 20772 20324
rect 24676 20272 24728 20324
rect 9680 20247 9732 20256
rect 9680 20213 9689 20247
rect 9689 20213 9723 20247
rect 9723 20213 9732 20247
rect 9680 20204 9732 20213
rect 13452 20247 13504 20256
rect 13452 20213 13461 20247
rect 13461 20213 13495 20247
rect 13495 20213 13504 20247
rect 13452 20204 13504 20213
rect 15108 20204 15160 20256
rect 25044 20247 25096 20256
rect 25044 20213 25053 20247
rect 25053 20213 25087 20247
rect 25087 20213 25096 20247
rect 25044 20204 25096 20213
rect 26332 20247 26384 20256
rect 26332 20213 26341 20247
rect 26341 20213 26375 20247
rect 26375 20213 26384 20247
rect 26332 20204 26384 20213
rect 26884 20204 26936 20256
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 20982 20102 21034 20154
rect 21046 20102 21098 20154
rect 21110 20102 21162 20154
rect 21174 20102 21226 20154
rect 3516 20043 3568 20052
rect 3516 20009 3525 20043
rect 3525 20009 3559 20043
rect 3559 20009 3568 20043
rect 3516 20000 3568 20009
rect 6644 20043 6696 20052
rect 6644 20009 6653 20043
rect 6653 20009 6687 20043
rect 6687 20009 6696 20043
rect 6644 20000 6696 20009
rect 13084 20000 13136 20052
rect 17040 20000 17092 20052
rect 17684 20043 17736 20052
rect 17684 20009 17693 20043
rect 17693 20009 17727 20043
rect 17727 20009 17736 20043
rect 17684 20000 17736 20009
rect 19248 20043 19300 20052
rect 19248 20009 19257 20043
rect 19257 20009 19291 20043
rect 19291 20009 19300 20043
rect 19248 20000 19300 20009
rect 28264 20000 28316 20052
rect 8024 19932 8076 19984
rect 5264 19907 5316 19916
rect 5264 19873 5273 19907
rect 5273 19873 5307 19907
rect 5307 19873 5316 19907
rect 5264 19864 5316 19873
rect 5540 19907 5592 19916
rect 5540 19873 5574 19907
rect 5574 19873 5592 19907
rect 5540 19864 5592 19873
rect 6736 19864 6788 19916
rect 6920 19728 6972 19780
rect 8208 19839 8260 19848
rect 8208 19805 8217 19839
rect 8217 19805 8251 19839
rect 8251 19805 8260 19839
rect 8208 19796 8260 19805
rect 8392 19864 8444 19916
rect 10692 19864 10744 19916
rect 10968 19932 11020 19984
rect 17316 19932 17368 19984
rect 21548 19932 21600 19984
rect 11612 19864 11664 19916
rect 16396 19864 16448 19916
rect 14004 19839 14056 19848
rect 14004 19805 14013 19839
rect 14013 19805 14047 19839
rect 14047 19805 14056 19839
rect 14004 19796 14056 19805
rect 15108 19796 15160 19848
rect 15844 19796 15896 19848
rect 16304 19839 16356 19848
rect 16304 19805 16313 19839
rect 16313 19805 16347 19839
rect 16347 19805 16356 19839
rect 16304 19796 16356 19805
rect 7748 19771 7800 19780
rect 7748 19737 7757 19771
rect 7757 19737 7791 19771
rect 7791 19737 7800 19771
rect 7748 19728 7800 19737
rect 13728 19728 13780 19780
rect 21640 19864 21692 19916
rect 26792 19864 26844 19916
rect 17868 19839 17920 19848
rect 17868 19805 17877 19839
rect 17877 19805 17911 19839
rect 17911 19805 17920 19839
rect 17868 19796 17920 19805
rect 3148 19703 3200 19712
rect 3148 19669 3157 19703
rect 3157 19669 3191 19703
rect 3191 19669 3200 19703
rect 3148 19660 3200 19669
rect 7196 19703 7248 19712
rect 7196 19669 7205 19703
rect 7205 19669 7239 19703
rect 7239 19669 7248 19703
rect 7196 19660 7248 19669
rect 8852 19703 8904 19712
rect 8852 19669 8861 19703
rect 8861 19669 8895 19703
rect 8895 19669 8904 19703
rect 8852 19660 8904 19669
rect 11428 19660 11480 19712
rect 13176 19660 13228 19712
rect 15108 19660 15160 19712
rect 22928 19703 22980 19712
rect 22928 19669 22937 19703
rect 22937 19669 22971 19703
rect 22971 19669 22980 19703
rect 22928 19660 22980 19669
rect 23756 19703 23808 19712
rect 23756 19669 23765 19703
rect 23765 19669 23799 19703
rect 23799 19669 23808 19703
rect 23756 19660 23808 19669
rect 25596 19660 25648 19712
rect 5982 19558 6034 19610
rect 6046 19558 6098 19610
rect 6110 19558 6162 19610
rect 6174 19558 6226 19610
rect 15982 19558 16034 19610
rect 16046 19558 16098 19610
rect 16110 19558 16162 19610
rect 16174 19558 16226 19610
rect 25982 19558 26034 19610
rect 26046 19558 26098 19610
rect 26110 19558 26162 19610
rect 26174 19558 26226 19610
rect 5264 19456 5316 19508
rect 8024 19456 8076 19508
rect 13084 19499 13136 19508
rect 13084 19465 13093 19499
rect 13093 19465 13127 19499
rect 13127 19465 13136 19499
rect 13084 19456 13136 19465
rect 13728 19499 13780 19508
rect 13728 19465 13737 19499
rect 13737 19465 13771 19499
rect 13771 19465 13780 19499
rect 13728 19456 13780 19465
rect 17684 19499 17736 19508
rect 17684 19465 17693 19499
rect 17693 19465 17727 19499
rect 17727 19465 17736 19499
rect 17684 19456 17736 19465
rect 20812 19456 20864 19508
rect 21640 19456 21692 19508
rect 23480 19499 23532 19508
rect 23480 19465 23489 19499
rect 23489 19465 23523 19499
rect 23523 19465 23532 19499
rect 23480 19456 23532 19465
rect 14004 19388 14056 19440
rect 17132 19388 17184 19440
rect 17868 19388 17920 19440
rect 3700 19363 3752 19372
rect 3700 19329 3709 19363
rect 3709 19329 3743 19363
rect 3743 19329 3752 19363
rect 3700 19320 3752 19329
rect 3148 19252 3200 19304
rect 5540 19320 5592 19372
rect 7748 19363 7800 19372
rect 7748 19329 7757 19363
rect 7757 19329 7791 19363
rect 7791 19329 7800 19363
rect 7748 19320 7800 19329
rect 8760 19363 8812 19372
rect 8760 19329 8769 19363
rect 8769 19329 8803 19363
rect 8803 19329 8812 19363
rect 8760 19320 8812 19329
rect 9680 19320 9732 19372
rect 11796 19320 11848 19372
rect 13912 19320 13964 19372
rect 8392 19252 8444 19304
rect 8852 19252 8904 19304
rect 10968 19252 11020 19304
rect 15108 19252 15160 19304
rect 20720 19252 20772 19304
rect 22928 19320 22980 19372
rect 22468 19252 22520 19304
rect 23756 19320 23808 19372
rect 24676 19388 24728 19440
rect 25044 19320 25096 19372
rect 26148 19320 26200 19372
rect 24860 19252 24912 19304
rect 25596 19295 25648 19304
rect 3056 19159 3108 19168
rect 3056 19125 3065 19159
rect 3065 19125 3099 19159
rect 3099 19125 3108 19159
rect 3056 19116 3108 19125
rect 8116 19184 8168 19236
rect 8300 19184 8352 19236
rect 3608 19116 3660 19168
rect 6552 19159 6604 19168
rect 6552 19125 6561 19159
rect 6561 19125 6595 19159
rect 6595 19125 6604 19159
rect 6552 19116 6604 19125
rect 7104 19159 7156 19168
rect 7104 19125 7113 19159
rect 7113 19125 7147 19159
rect 7147 19125 7156 19159
rect 7104 19116 7156 19125
rect 7196 19116 7248 19168
rect 14740 19184 14792 19236
rect 25596 19261 25605 19295
rect 25605 19261 25639 19295
rect 25639 19261 25648 19295
rect 25596 19252 25648 19261
rect 9312 19159 9364 19168
rect 9312 19125 9321 19159
rect 9321 19125 9355 19159
rect 9355 19125 9364 19159
rect 9312 19116 9364 19125
rect 10600 19116 10652 19168
rect 10784 19116 10836 19168
rect 14280 19116 14332 19168
rect 16304 19159 16356 19168
rect 16304 19125 16313 19159
rect 16313 19125 16347 19159
rect 16347 19125 16356 19159
rect 16304 19116 16356 19125
rect 17316 19159 17368 19168
rect 17316 19125 17325 19159
rect 17325 19125 17359 19159
rect 17359 19125 17368 19159
rect 17316 19116 17368 19125
rect 21548 19159 21600 19168
rect 21548 19125 21557 19159
rect 21557 19125 21591 19159
rect 21591 19125 21600 19159
rect 21548 19116 21600 19125
rect 21916 19116 21968 19168
rect 22652 19116 22704 19168
rect 25872 19184 25924 19236
rect 26792 19116 26844 19168
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 20982 19014 21034 19066
rect 21046 19014 21098 19066
rect 21110 19014 21162 19066
rect 21174 19014 21226 19066
rect 3056 18912 3108 18964
rect 3424 18955 3476 18964
rect 3424 18921 3433 18955
rect 3433 18921 3467 18955
rect 3467 18921 3476 18955
rect 3424 18912 3476 18921
rect 7196 18912 7248 18964
rect 7564 18955 7616 18964
rect 7564 18921 7573 18955
rect 7573 18921 7607 18955
rect 7607 18921 7616 18955
rect 7564 18912 7616 18921
rect 8300 18955 8352 18964
rect 8300 18921 8309 18955
rect 8309 18921 8343 18955
rect 8343 18921 8352 18955
rect 8300 18912 8352 18921
rect 13728 18912 13780 18964
rect 15844 18955 15896 18964
rect 15844 18921 15853 18955
rect 15853 18921 15887 18955
rect 15887 18921 15896 18955
rect 15844 18912 15896 18921
rect 22652 18955 22704 18964
rect 22652 18921 22661 18955
rect 22661 18921 22695 18955
rect 22695 18921 22704 18955
rect 22652 18912 22704 18921
rect 23756 18912 23808 18964
rect 4160 18844 4212 18896
rect 4436 18887 4488 18896
rect 4436 18853 4445 18887
rect 4445 18853 4479 18887
rect 4479 18853 4488 18887
rect 4436 18844 4488 18853
rect 6736 18844 6788 18896
rect 7380 18844 7432 18896
rect 8760 18844 8812 18896
rect 10876 18887 10928 18896
rect 10876 18853 10910 18887
rect 10910 18853 10928 18887
rect 10876 18844 10928 18853
rect 11428 18844 11480 18896
rect 16396 18844 16448 18896
rect 1768 18819 1820 18828
rect 1768 18785 1802 18819
rect 1802 18785 1820 18819
rect 1768 18776 1820 18785
rect 3700 18776 3752 18828
rect 1492 18751 1544 18760
rect 1492 18717 1501 18751
rect 1501 18717 1535 18751
rect 1535 18717 1544 18751
rect 1492 18708 1544 18717
rect 4528 18751 4580 18760
rect 4528 18717 4537 18751
rect 4537 18717 4571 18751
rect 4571 18717 4580 18751
rect 4528 18708 4580 18717
rect 13636 18776 13688 18828
rect 13820 18776 13872 18828
rect 4804 18708 4856 18760
rect 7656 18751 7708 18760
rect 7656 18717 7665 18751
rect 7665 18717 7699 18751
rect 7699 18717 7708 18751
rect 7656 18708 7708 18717
rect 7748 18708 7800 18760
rect 8576 18708 8628 18760
rect 10600 18751 10652 18760
rect 10600 18717 10609 18751
rect 10609 18717 10643 18751
rect 10643 18717 10652 18751
rect 10600 18708 10652 18717
rect 14188 18751 14240 18760
rect 14188 18717 14197 18751
rect 14197 18717 14231 18751
rect 14231 18717 14240 18751
rect 14188 18708 14240 18717
rect 12348 18640 12400 18692
rect 16580 18640 16632 18692
rect 17040 18819 17092 18828
rect 17040 18785 17049 18819
rect 17049 18785 17083 18819
rect 17083 18785 17092 18819
rect 17040 18776 17092 18785
rect 17868 18776 17920 18828
rect 19248 18844 19300 18896
rect 22468 18887 22520 18896
rect 22468 18853 22477 18887
rect 22477 18853 22511 18887
rect 22511 18853 22520 18887
rect 22468 18844 22520 18853
rect 18420 18776 18472 18828
rect 23020 18819 23072 18828
rect 23020 18785 23029 18819
rect 23029 18785 23063 18819
rect 23063 18785 23072 18819
rect 23020 18776 23072 18785
rect 24768 18819 24820 18828
rect 24768 18785 24777 18819
rect 24777 18785 24811 18819
rect 24811 18785 24820 18819
rect 24768 18776 24820 18785
rect 25136 18776 25188 18828
rect 17132 18751 17184 18760
rect 17132 18717 17141 18751
rect 17141 18717 17175 18751
rect 17175 18717 17184 18751
rect 17132 18708 17184 18717
rect 21364 18708 21416 18760
rect 23112 18751 23164 18760
rect 23112 18717 23121 18751
rect 23121 18717 23155 18751
rect 23155 18717 23164 18751
rect 23112 18708 23164 18717
rect 23480 18708 23532 18760
rect 24676 18708 24728 18760
rect 2872 18615 2924 18624
rect 2872 18581 2881 18615
rect 2881 18581 2915 18615
rect 2915 18581 2924 18615
rect 2872 18572 2924 18581
rect 3516 18572 3568 18624
rect 7196 18615 7248 18624
rect 7196 18581 7205 18615
rect 7205 18581 7239 18615
rect 7239 18581 7248 18615
rect 7196 18572 7248 18581
rect 9312 18572 9364 18624
rect 9772 18572 9824 18624
rect 9956 18615 10008 18624
rect 9956 18581 9965 18615
rect 9965 18581 9999 18615
rect 9999 18581 10008 18615
rect 9956 18572 10008 18581
rect 10416 18572 10468 18624
rect 19708 18615 19760 18624
rect 19708 18581 19717 18615
rect 19717 18581 19751 18615
rect 19751 18581 19760 18615
rect 19708 18572 19760 18581
rect 21272 18572 21324 18624
rect 5982 18470 6034 18522
rect 6046 18470 6098 18522
rect 6110 18470 6162 18522
rect 6174 18470 6226 18522
rect 15982 18470 16034 18522
rect 16046 18470 16098 18522
rect 16110 18470 16162 18522
rect 16174 18470 16226 18522
rect 25982 18470 26034 18522
rect 26046 18470 26098 18522
rect 26110 18470 26162 18522
rect 26174 18470 26226 18522
rect 1768 18368 1820 18420
rect 4528 18411 4580 18420
rect 4528 18377 4537 18411
rect 4537 18377 4571 18411
rect 4571 18377 4580 18411
rect 4528 18368 4580 18377
rect 6828 18411 6880 18420
rect 6828 18377 6837 18411
rect 6837 18377 6871 18411
rect 6871 18377 6880 18411
rect 6828 18368 6880 18377
rect 7564 18368 7616 18420
rect 9772 18411 9824 18420
rect 9772 18377 9781 18411
rect 9781 18377 9815 18411
rect 9815 18377 9824 18411
rect 9772 18368 9824 18377
rect 10876 18411 10928 18420
rect 10876 18377 10885 18411
rect 10885 18377 10919 18411
rect 10919 18377 10928 18411
rect 10876 18368 10928 18377
rect 13452 18368 13504 18420
rect 14188 18368 14240 18420
rect 16580 18411 16632 18420
rect 16580 18377 16589 18411
rect 16589 18377 16623 18411
rect 16623 18377 16632 18411
rect 16580 18368 16632 18377
rect 17040 18411 17092 18420
rect 17040 18377 17049 18411
rect 17049 18377 17083 18411
rect 17083 18377 17092 18411
rect 17040 18368 17092 18377
rect 17132 18368 17184 18420
rect 17868 18411 17920 18420
rect 17868 18377 17877 18411
rect 17877 18377 17911 18411
rect 17911 18377 17920 18411
rect 17868 18368 17920 18377
rect 19340 18411 19392 18420
rect 19340 18377 19349 18411
rect 19349 18377 19383 18411
rect 19383 18377 19392 18411
rect 21180 18411 21232 18420
rect 19340 18368 19392 18377
rect 1492 18300 1544 18352
rect 2872 18300 2924 18352
rect 4436 18300 4488 18352
rect 7748 18300 7800 18352
rect 13820 18300 13872 18352
rect 3516 18275 3568 18284
rect 3516 18241 3525 18275
rect 3525 18241 3559 18275
rect 3559 18241 3568 18275
rect 3516 18232 3568 18241
rect 3700 18275 3752 18284
rect 3700 18241 3709 18275
rect 3709 18241 3743 18275
rect 3743 18241 3752 18275
rect 3700 18232 3752 18241
rect 7196 18232 7248 18284
rect 7380 18275 7432 18284
rect 7380 18241 7389 18275
rect 7389 18241 7423 18275
rect 7423 18241 7432 18275
rect 7380 18232 7432 18241
rect 9588 18232 9640 18284
rect 10416 18275 10468 18284
rect 10416 18241 10425 18275
rect 10425 18241 10459 18275
rect 10459 18241 10468 18275
rect 10416 18232 10468 18241
rect 13544 18232 13596 18284
rect 14740 18275 14792 18284
rect 14740 18241 14749 18275
rect 14749 18241 14783 18275
rect 14783 18241 14792 18275
rect 14740 18232 14792 18241
rect 3424 18207 3476 18216
rect 3424 18173 3433 18207
rect 3433 18173 3467 18207
rect 3467 18173 3476 18207
rect 3424 18164 3476 18173
rect 21180 18377 21189 18411
rect 21189 18377 21223 18411
rect 21223 18377 21232 18411
rect 21180 18368 21232 18377
rect 21548 18368 21600 18420
rect 23480 18368 23532 18420
rect 26332 18368 26384 18420
rect 20720 18300 20772 18352
rect 23020 18300 23072 18352
rect 25136 18343 25188 18352
rect 25136 18309 25145 18343
rect 25145 18309 25179 18343
rect 25179 18309 25188 18343
rect 25136 18300 25188 18309
rect 9956 18164 10008 18216
rect 20168 18207 20220 18216
rect 20168 18173 20177 18207
rect 20177 18173 20211 18207
rect 20211 18173 20220 18207
rect 20168 18164 20220 18173
rect 7104 18096 7156 18148
rect 10324 18096 10376 18148
rect 13636 18096 13688 18148
rect 21272 18232 21324 18284
rect 24676 18232 24728 18284
rect 21364 18164 21416 18216
rect 23572 18164 23624 18216
rect 24768 18207 24820 18216
rect 24768 18173 24777 18207
rect 24777 18173 24811 18207
rect 24811 18173 24820 18207
rect 24768 18164 24820 18173
rect 26148 18207 26200 18216
rect 26148 18173 26157 18207
rect 26157 18173 26191 18207
rect 26191 18173 26200 18207
rect 26148 18164 26200 18173
rect 3056 18071 3108 18080
rect 3056 18037 3065 18071
rect 3065 18037 3099 18071
rect 3099 18037 3108 18071
rect 3056 18028 3108 18037
rect 4804 18071 4856 18080
rect 4804 18037 4813 18071
rect 4813 18037 4847 18071
rect 4847 18037 4856 18071
rect 4804 18028 4856 18037
rect 10600 18028 10652 18080
rect 12348 18028 12400 18080
rect 13820 18028 13872 18080
rect 15292 18028 15344 18080
rect 18420 18071 18472 18080
rect 18420 18037 18429 18071
rect 18429 18037 18463 18071
rect 18463 18037 18472 18071
rect 21180 18096 21232 18148
rect 21824 18139 21876 18148
rect 21824 18105 21833 18139
rect 21833 18105 21867 18139
rect 21867 18105 21876 18139
rect 21824 18096 21876 18105
rect 23940 18096 23992 18148
rect 18420 18028 18472 18037
rect 19800 18071 19852 18080
rect 19800 18037 19809 18071
rect 19809 18037 19843 18071
rect 19843 18037 19852 18071
rect 19800 18028 19852 18037
rect 23480 18071 23532 18080
rect 23480 18037 23489 18071
rect 23489 18037 23523 18071
rect 23523 18037 23532 18071
rect 24032 18071 24084 18080
rect 23480 18028 23532 18037
rect 24032 18037 24041 18071
rect 24041 18037 24075 18071
rect 24075 18037 24084 18071
rect 24032 18028 24084 18037
rect 24860 18028 24912 18080
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 20982 17926 21034 17978
rect 21046 17926 21098 17978
rect 21110 17926 21162 17978
rect 21174 17926 21226 17978
rect 7104 17824 7156 17876
rect 8208 17824 8260 17876
rect 10324 17867 10376 17876
rect 10324 17833 10333 17867
rect 10333 17833 10367 17867
rect 10367 17833 10376 17867
rect 10324 17824 10376 17833
rect 13728 17824 13780 17876
rect 17132 17824 17184 17876
rect 19800 17824 19852 17876
rect 21364 17867 21416 17876
rect 21364 17833 21373 17867
rect 21373 17833 21407 17867
rect 21407 17833 21416 17867
rect 21364 17824 21416 17833
rect 23020 17867 23072 17876
rect 23020 17833 23029 17867
rect 23029 17833 23063 17867
rect 23063 17833 23072 17867
rect 23020 17824 23072 17833
rect 23112 17824 23164 17876
rect 24676 17824 24728 17876
rect 26240 17867 26292 17876
rect 26240 17833 26249 17867
rect 26249 17833 26283 17867
rect 26283 17833 26292 17867
rect 26240 17824 26292 17833
rect 7656 17756 7708 17808
rect 15108 17756 15160 17808
rect 1676 17688 1728 17740
rect 3608 17688 3660 17740
rect 5264 17731 5316 17740
rect 5264 17697 5273 17731
rect 5273 17697 5307 17731
rect 5307 17697 5316 17731
rect 5264 17688 5316 17697
rect 5356 17688 5408 17740
rect 8024 17688 8076 17740
rect 10692 17731 10744 17740
rect 10692 17697 10701 17731
rect 10701 17697 10735 17731
rect 10735 17697 10744 17731
rect 10692 17688 10744 17697
rect 14004 17731 14056 17740
rect 14004 17697 14013 17731
rect 14013 17697 14047 17731
rect 14047 17697 14056 17731
rect 14004 17688 14056 17697
rect 16304 17756 16356 17808
rect 17868 17756 17920 17808
rect 20076 17756 20128 17808
rect 20628 17756 20680 17808
rect 16488 17731 16540 17740
rect 16488 17697 16522 17731
rect 16522 17697 16540 17731
rect 16488 17688 16540 17697
rect 23756 17731 23808 17740
rect 23756 17697 23765 17731
rect 23765 17697 23799 17731
rect 23799 17697 23808 17731
rect 23756 17688 23808 17697
rect 24032 17688 24084 17740
rect 8484 17663 8536 17672
rect 8484 17629 8493 17663
rect 8493 17629 8527 17663
rect 8527 17629 8536 17663
rect 8484 17620 8536 17629
rect 8576 17620 8628 17672
rect 9588 17620 9640 17672
rect 10784 17663 10836 17672
rect 10784 17629 10793 17663
rect 10793 17629 10827 17663
rect 10827 17629 10836 17663
rect 10784 17620 10836 17629
rect 10876 17663 10928 17672
rect 10876 17629 10885 17663
rect 10885 17629 10919 17663
rect 10919 17629 10928 17663
rect 14096 17663 14148 17672
rect 10876 17620 10928 17629
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 14740 17620 14792 17672
rect 19708 17620 19760 17672
rect 23112 17620 23164 17672
rect 13636 17595 13688 17604
rect 13636 17561 13645 17595
rect 13645 17561 13679 17595
rect 13679 17561 13688 17595
rect 13636 17552 13688 17561
rect 18236 17595 18288 17604
rect 18236 17561 18245 17595
rect 18245 17561 18279 17595
rect 18279 17561 18288 17595
rect 18236 17552 18288 17561
rect 1584 17527 1636 17536
rect 1584 17493 1593 17527
rect 1593 17493 1627 17527
rect 1627 17493 1636 17527
rect 1584 17484 1636 17493
rect 2872 17527 2924 17536
rect 2872 17493 2881 17527
rect 2881 17493 2915 17527
rect 2915 17493 2924 17527
rect 2872 17484 2924 17493
rect 3148 17527 3200 17536
rect 3148 17493 3157 17527
rect 3157 17493 3191 17527
rect 3191 17493 3200 17527
rect 3148 17484 3200 17493
rect 7104 17484 7156 17536
rect 15752 17484 15804 17536
rect 16396 17484 16448 17536
rect 19248 17527 19300 17536
rect 19248 17493 19257 17527
rect 19257 17493 19291 17527
rect 19291 17493 19300 17527
rect 19248 17484 19300 17493
rect 24676 17484 24728 17536
rect 5982 17382 6034 17434
rect 6046 17382 6098 17434
rect 6110 17382 6162 17434
rect 6174 17382 6226 17434
rect 15982 17382 16034 17434
rect 16046 17382 16098 17434
rect 16110 17382 16162 17434
rect 16174 17382 16226 17434
rect 25982 17382 26034 17434
rect 26046 17382 26098 17434
rect 26110 17382 26162 17434
rect 26174 17382 26226 17434
rect 2044 17323 2096 17332
rect 2044 17289 2053 17323
rect 2053 17289 2087 17323
rect 2087 17289 2096 17323
rect 2044 17280 2096 17289
rect 5356 17323 5408 17332
rect 5356 17289 5365 17323
rect 5365 17289 5399 17323
rect 5399 17289 5408 17323
rect 5356 17280 5408 17289
rect 8484 17280 8536 17332
rect 10876 17280 10928 17332
rect 14004 17280 14056 17332
rect 17776 17323 17828 17332
rect 17776 17289 17785 17323
rect 17785 17289 17819 17323
rect 17819 17289 17828 17323
rect 17776 17280 17828 17289
rect 19800 17280 19852 17332
rect 20076 17323 20128 17332
rect 20076 17289 20085 17323
rect 20085 17289 20119 17323
rect 20119 17289 20128 17323
rect 20076 17280 20128 17289
rect 23112 17323 23164 17332
rect 23112 17289 23121 17323
rect 23121 17289 23155 17323
rect 23155 17289 23164 17323
rect 23112 17280 23164 17289
rect 2872 17144 2924 17196
rect 3240 17187 3292 17196
rect 3240 17153 3249 17187
rect 3249 17153 3283 17187
rect 3283 17153 3292 17187
rect 3240 17144 3292 17153
rect 3700 17144 3752 17196
rect 9496 17255 9548 17264
rect 9496 17221 9505 17255
rect 9505 17221 9539 17255
rect 9539 17221 9548 17255
rect 9496 17212 9548 17221
rect 10692 17212 10744 17264
rect 8576 17144 8628 17196
rect 14096 17212 14148 17264
rect 18420 17212 18472 17264
rect 13544 17187 13596 17196
rect 13544 17153 13553 17187
rect 13553 17153 13587 17187
rect 13587 17153 13596 17187
rect 13544 17144 13596 17153
rect 13912 17144 13964 17196
rect 15844 17144 15896 17196
rect 16488 17144 16540 17196
rect 18236 17144 18288 17196
rect 18880 17144 18932 17196
rect 19708 17144 19760 17196
rect 24676 17187 24728 17196
rect 24676 17153 24685 17187
rect 24685 17153 24719 17187
rect 24719 17153 24728 17187
rect 24676 17144 24728 17153
rect 2044 17076 2096 17128
rect 3148 17119 3200 17128
rect 3148 17085 3157 17119
rect 3157 17085 3191 17119
rect 3191 17085 3200 17119
rect 3148 17076 3200 17085
rect 5264 17076 5316 17128
rect 14832 17119 14884 17128
rect 14832 17085 14841 17119
rect 14841 17085 14875 17119
rect 14875 17085 14884 17119
rect 14832 17076 14884 17085
rect 16396 17119 16448 17128
rect 16396 17085 16405 17119
rect 16405 17085 16439 17119
rect 16439 17085 16448 17119
rect 16396 17076 16448 17085
rect 16764 17076 16816 17128
rect 17776 17076 17828 17128
rect 18512 17119 18564 17128
rect 18512 17085 18521 17119
rect 18521 17085 18555 17119
rect 18555 17085 18564 17119
rect 18512 17076 18564 17085
rect 23480 17119 23532 17128
rect 23480 17085 23489 17119
rect 23489 17085 23523 17119
rect 23523 17085 23532 17119
rect 26424 17119 26476 17128
rect 23480 17076 23532 17085
rect 10232 17008 10284 17060
rect 10784 17008 10836 17060
rect 18604 17008 18656 17060
rect 23756 17008 23808 17060
rect 26424 17085 26433 17119
rect 26433 17085 26467 17119
rect 26467 17085 26476 17119
rect 26424 17076 26476 17085
rect 1860 16940 1912 16992
rect 4068 16940 4120 16992
rect 8024 16983 8076 16992
rect 8024 16949 8033 16983
rect 8033 16949 8067 16983
rect 8067 16949 8076 16983
rect 8024 16940 8076 16949
rect 10324 16983 10376 16992
rect 10324 16949 10333 16983
rect 10333 16949 10367 16983
rect 10367 16949 10376 16983
rect 10324 16940 10376 16949
rect 13912 16983 13964 16992
rect 13912 16949 13921 16983
rect 13921 16949 13955 16983
rect 13955 16949 13964 16983
rect 13912 16940 13964 16949
rect 14924 16983 14976 16992
rect 14924 16949 14933 16983
rect 14933 16949 14967 16983
rect 14967 16949 14976 16983
rect 14924 16940 14976 16949
rect 17960 16940 18012 16992
rect 23848 16983 23900 16992
rect 23848 16949 23857 16983
rect 23857 16949 23891 16983
rect 23891 16949 23900 16983
rect 23848 16940 23900 16949
rect 24032 16983 24084 16992
rect 24032 16949 24041 16983
rect 24041 16949 24075 16983
rect 24075 16949 24084 16983
rect 24032 16940 24084 16949
rect 27344 17008 27396 17060
rect 25872 16940 25924 16992
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 20982 16838 21034 16890
rect 21046 16838 21098 16890
rect 21110 16838 21162 16890
rect 21174 16838 21226 16890
rect 1676 16779 1728 16788
rect 1676 16745 1685 16779
rect 1685 16745 1719 16779
rect 1719 16745 1728 16779
rect 1676 16736 1728 16745
rect 3148 16736 3200 16788
rect 4804 16736 4856 16788
rect 4988 16736 5040 16788
rect 5724 16779 5776 16788
rect 5724 16745 5733 16779
rect 5733 16745 5767 16779
rect 5767 16745 5776 16779
rect 5724 16736 5776 16745
rect 9956 16736 10008 16788
rect 13912 16736 13964 16788
rect 14832 16736 14884 16788
rect 15292 16779 15344 16788
rect 15292 16745 15301 16779
rect 15301 16745 15335 16779
rect 15335 16745 15344 16779
rect 15292 16736 15344 16745
rect 15752 16779 15804 16788
rect 15752 16745 15761 16779
rect 15761 16745 15795 16779
rect 15795 16745 15804 16779
rect 15752 16736 15804 16745
rect 16304 16779 16356 16788
rect 16304 16745 16313 16779
rect 16313 16745 16347 16779
rect 16347 16745 16356 16779
rect 16304 16736 16356 16745
rect 17960 16736 18012 16788
rect 19248 16779 19300 16788
rect 19248 16745 19257 16779
rect 19257 16745 19291 16779
rect 19291 16745 19300 16779
rect 19248 16736 19300 16745
rect 24032 16736 24084 16788
rect 2688 16668 2740 16720
rect 5632 16711 5684 16720
rect 5632 16677 5641 16711
rect 5641 16677 5675 16711
rect 5675 16677 5684 16711
rect 5632 16668 5684 16677
rect 9864 16668 9916 16720
rect 11060 16668 11112 16720
rect 15660 16711 15712 16720
rect 15660 16677 15669 16711
rect 15669 16677 15703 16711
rect 15703 16677 15712 16711
rect 15660 16668 15712 16677
rect 5264 16600 5316 16652
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 7104 16643 7156 16652
rect 7104 16609 7138 16643
rect 7138 16609 7156 16643
rect 7104 16600 7156 16609
rect 10968 16600 11020 16652
rect 12532 16600 12584 16652
rect 2872 16575 2924 16584
rect 2872 16541 2881 16575
rect 2881 16541 2915 16575
rect 2915 16541 2924 16575
rect 2872 16532 2924 16541
rect 3056 16575 3108 16584
rect 3056 16541 3065 16575
rect 3065 16541 3099 16575
rect 3099 16541 3108 16575
rect 3056 16532 3108 16541
rect 5816 16575 5868 16584
rect 5816 16541 5825 16575
rect 5825 16541 5859 16575
rect 5859 16541 5868 16575
rect 5816 16532 5868 16541
rect 10876 16575 10928 16584
rect 10876 16541 10885 16575
rect 10885 16541 10919 16575
rect 10919 16541 10928 16575
rect 10876 16532 10928 16541
rect 12348 16532 12400 16584
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 18696 16575 18748 16584
rect 18696 16541 18705 16575
rect 18705 16541 18739 16575
rect 18739 16541 18748 16575
rect 18696 16532 18748 16541
rect 18788 16575 18840 16584
rect 18788 16541 18797 16575
rect 18797 16541 18831 16575
rect 18831 16541 18840 16575
rect 19708 16600 19760 16652
rect 20996 16600 21048 16652
rect 23756 16600 23808 16652
rect 18788 16532 18840 16541
rect 20720 16532 20772 16584
rect 24308 16600 24360 16652
rect 24492 16575 24544 16584
rect 24492 16541 24501 16575
rect 24501 16541 24535 16575
rect 24535 16541 24544 16575
rect 24492 16532 24544 16541
rect 24676 16575 24728 16584
rect 24676 16541 24685 16575
rect 24685 16541 24719 16575
rect 24719 16541 24728 16575
rect 24676 16532 24728 16541
rect 24860 16532 24912 16584
rect 8208 16439 8260 16448
rect 8208 16405 8217 16439
rect 8217 16405 8251 16439
rect 8251 16405 8260 16439
rect 8208 16396 8260 16405
rect 10324 16396 10376 16448
rect 12716 16396 12768 16448
rect 19156 16396 19208 16448
rect 21824 16396 21876 16448
rect 5982 16294 6034 16346
rect 6046 16294 6098 16346
rect 6110 16294 6162 16346
rect 6174 16294 6226 16346
rect 15982 16294 16034 16346
rect 16046 16294 16098 16346
rect 16110 16294 16162 16346
rect 16174 16294 16226 16346
rect 25982 16294 26034 16346
rect 26046 16294 26098 16346
rect 26110 16294 26162 16346
rect 26174 16294 26226 16346
rect 3240 16192 3292 16244
rect 5816 16192 5868 16244
rect 7104 16192 7156 16244
rect 11060 16192 11112 16244
rect 15476 16192 15528 16244
rect 15752 16192 15804 16244
rect 15844 16192 15896 16244
rect 17868 16235 17920 16244
rect 17868 16201 17877 16235
rect 17877 16201 17911 16235
rect 17911 16201 17920 16235
rect 17868 16192 17920 16201
rect 18696 16235 18748 16244
rect 18696 16201 18705 16235
rect 18705 16201 18739 16235
rect 18739 16201 18748 16235
rect 18696 16192 18748 16201
rect 20996 16235 21048 16244
rect 20996 16201 21005 16235
rect 21005 16201 21039 16235
rect 21039 16201 21048 16235
rect 20996 16192 21048 16201
rect 23940 16235 23992 16244
rect 23940 16201 23949 16235
rect 23949 16201 23983 16235
rect 23983 16201 23992 16235
rect 23940 16192 23992 16201
rect 5724 16167 5776 16176
rect 5724 16133 5733 16167
rect 5733 16133 5767 16167
rect 5767 16133 5776 16167
rect 5724 16124 5776 16133
rect 6920 16124 6972 16176
rect 11336 16124 11388 16176
rect 15660 16167 15712 16176
rect 15660 16133 15669 16167
rect 15669 16133 15703 16167
rect 15703 16133 15712 16167
rect 15660 16124 15712 16133
rect 18788 16124 18840 16176
rect 3056 16056 3108 16108
rect 4804 16056 4856 16108
rect 5632 16056 5684 16108
rect 19156 16056 19208 16108
rect 20720 16124 20772 16176
rect 21732 16124 21784 16176
rect 21824 16056 21876 16108
rect 24860 16192 24912 16244
rect 1492 15988 1544 16040
rect 8852 16031 8904 16040
rect 8852 15997 8861 16031
rect 8861 15997 8895 16031
rect 8895 15997 8904 16031
rect 8852 15988 8904 15997
rect 19340 15988 19392 16040
rect 23112 16031 23164 16040
rect 23112 15997 23121 16031
rect 23121 15997 23155 16031
rect 23155 15997 23164 16031
rect 23112 15988 23164 15997
rect 24400 15988 24452 16040
rect 25964 15988 26016 16040
rect 1676 15963 1728 15972
rect 1676 15929 1710 15963
rect 1710 15929 1728 15963
rect 1676 15920 1728 15929
rect 3608 15920 3660 15972
rect 4252 15963 4304 15972
rect 4252 15929 4261 15963
rect 4261 15929 4295 15963
rect 4295 15929 4304 15963
rect 4252 15920 4304 15929
rect 9036 15920 9088 15972
rect 10968 15920 11020 15972
rect 4068 15852 4120 15904
rect 12440 15852 12492 15904
rect 12992 15895 13044 15904
rect 12992 15861 13001 15895
rect 13001 15861 13035 15895
rect 13035 15861 13044 15895
rect 12992 15852 13044 15861
rect 19064 15852 19116 15904
rect 23940 15852 23992 15904
rect 25228 15852 25280 15904
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 20982 15750 21034 15802
rect 21046 15750 21098 15802
rect 21110 15750 21162 15802
rect 21174 15750 21226 15802
rect 1492 15648 1544 15700
rect 1768 15648 1820 15700
rect 2688 15648 2740 15700
rect 2872 15691 2924 15700
rect 2872 15657 2881 15691
rect 2881 15657 2915 15691
rect 2915 15657 2924 15691
rect 2872 15648 2924 15657
rect 4068 15691 4120 15700
rect 4068 15657 4077 15691
rect 4077 15657 4111 15691
rect 4111 15657 4120 15691
rect 4068 15648 4120 15657
rect 10876 15648 10928 15700
rect 4436 15623 4488 15632
rect 4436 15589 4445 15623
rect 4445 15589 4479 15623
rect 4479 15589 4488 15623
rect 4436 15580 4488 15589
rect 11336 15580 11388 15632
rect 16304 15648 16356 15700
rect 18696 15648 18748 15700
rect 19156 15691 19208 15700
rect 19156 15657 19165 15691
rect 19165 15657 19199 15691
rect 19199 15657 19208 15691
rect 19156 15648 19208 15657
rect 24492 15648 24544 15700
rect 24860 15691 24912 15700
rect 24860 15657 24869 15691
rect 24869 15657 24903 15691
rect 24903 15657 24912 15691
rect 24860 15648 24912 15657
rect 25964 15691 26016 15700
rect 25964 15657 25973 15691
rect 25973 15657 26007 15691
rect 26007 15657 26016 15691
rect 25964 15648 26016 15657
rect 21824 15580 21876 15632
rect 8300 15512 8352 15564
rect 9588 15512 9640 15564
rect 15292 15555 15344 15564
rect 15292 15521 15301 15555
rect 15301 15521 15335 15555
rect 15335 15521 15344 15555
rect 15292 15512 15344 15521
rect 15384 15512 15436 15564
rect 17960 15555 18012 15564
rect 17960 15521 17969 15555
rect 17969 15521 18003 15555
rect 18003 15521 18012 15555
rect 17960 15512 18012 15521
rect 18420 15555 18472 15564
rect 18420 15521 18429 15555
rect 18429 15521 18463 15555
rect 18463 15521 18472 15555
rect 18420 15512 18472 15521
rect 21732 15555 21784 15564
rect 21732 15521 21741 15555
rect 21741 15521 21775 15555
rect 21775 15521 21784 15555
rect 21732 15512 21784 15521
rect 26516 15555 26568 15564
rect 26516 15521 26525 15555
rect 26525 15521 26559 15555
rect 26559 15521 26568 15555
rect 26516 15512 26568 15521
rect 4528 15487 4580 15496
rect 4528 15453 4537 15487
rect 4537 15453 4571 15487
rect 4571 15453 4580 15487
rect 4528 15444 4580 15453
rect 1676 15419 1728 15428
rect 1676 15385 1685 15419
rect 1685 15385 1719 15419
rect 1719 15385 1728 15419
rect 4896 15444 4948 15496
rect 1676 15376 1728 15385
rect 7656 15308 7708 15360
rect 8484 15308 8536 15360
rect 8852 15351 8904 15360
rect 8852 15317 8861 15351
rect 8861 15317 8895 15351
rect 8895 15317 8904 15351
rect 11244 15444 11296 15496
rect 18512 15487 18564 15496
rect 18512 15453 18521 15487
rect 18521 15453 18555 15487
rect 18555 15453 18564 15487
rect 18512 15444 18564 15453
rect 18052 15376 18104 15428
rect 18880 15376 18932 15428
rect 19248 15376 19300 15428
rect 8852 15308 8904 15317
rect 12440 15308 12492 15360
rect 16672 15351 16724 15360
rect 16672 15317 16681 15351
rect 16681 15317 16715 15351
rect 16715 15317 16724 15351
rect 16672 15308 16724 15317
rect 23112 15351 23164 15360
rect 23112 15317 23121 15351
rect 23121 15317 23155 15351
rect 23155 15317 23164 15351
rect 23112 15308 23164 15317
rect 24308 15308 24360 15360
rect 24768 15308 24820 15360
rect 27252 15308 27304 15360
rect 5982 15206 6034 15258
rect 6046 15206 6098 15258
rect 6110 15206 6162 15258
rect 6174 15206 6226 15258
rect 15982 15206 16034 15258
rect 16046 15206 16098 15258
rect 16110 15206 16162 15258
rect 16174 15206 16226 15258
rect 25982 15206 26034 15258
rect 26046 15206 26098 15258
rect 26110 15206 26162 15258
rect 26174 15206 26226 15258
rect 1400 15104 1452 15156
rect 1768 15104 1820 15156
rect 4436 15147 4488 15156
rect 4436 15113 4445 15147
rect 4445 15113 4479 15147
rect 4479 15113 4488 15147
rect 4436 15104 4488 15113
rect 5172 15104 5224 15156
rect 6828 15104 6880 15156
rect 7932 15104 7984 15156
rect 8300 15104 8352 15156
rect 9036 15147 9088 15156
rect 9036 15113 9045 15147
rect 9045 15113 9079 15147
rect 9079 15113 9088 15147
rect 9036 15104 9088 15113
rect 9680 15147 9732 15156
rect 9680 15113 9689 15147
rect 9689 15113 9723 15147
rect 9723 15113 9732 15147
rect 9680 15104 9732 15113
rect 11244 15104 11296 15156
rect 12348 15104 12400 15156
rect 12992 15104 13044 15156
rect 15384 15147 15436 15156
rect 15384 15113 15393 15147
rect 15393 15113 15427 15147
rect 15427 15113 15436 15147
rect 15384 15104 15436 15113
rect 16304 15104 16356 15156
rect 17960 15104 18012 15156
rect 18420 15104 18472 15156
rect 19340 15104 19392 15156
rect 21732 15104 21784 15156
rect 21824 15104 21876 15156
rect 26516 15147 26568 15156
rect 26516 15113 26525 15147
rect 26525 15113 26559 15147
rect 26559 15113 26568 15147
rect 26516 15104 26568 15113
rect 18052 15036 18104 15088
rect 7656 15011 7708 15020
rect 7656 14977 7665 15011
rect 7665 14977 7699 15011
rect 7699 14977 7708 15011
rect 7656 14968 7708 14977
rect 25228 15011 25280 15020
rect 25228 14977 25237 15011
rect 25237 14977 25271 15011
rect 25271 14977 25280 15011
rect 25228 14968 25280 14977
rect 8208 14900 8260 14952
rect 18972 14943 19024 14952
rect 18972 14909 18981 14943
rect 18981 14909 19015 14943
rect 19015 14909 19024 14943
rect 18972 14900 19024 14909
rect 19892 14832 19944 14884
rect 26148 14832 26200 14884
rect 4528 14764 4580 14816
rect 4896 14807 4948 14816
rect 4896 14773 4905 14807
rect 4905 14773 4939 14807
rect 4939 14773 4948 14807
rect 4896 14764 4948 14773
rect 11336 14807 11388 14816
rect 11336 14773 11345 14807
rect 11345 14773 11379 14807
rect 11379 14773 11388 14807
rect 11336 14764 11388 14773
rect 18880 14807 18932 14816
rect 18880 14773 18889 14807
rect 18889 14773 18923 14807
rect 18923 14773 18932 14807
rect 18880 14764 18932 14773
rect 24492 14764 24544 14816
rect 25044 14807 25096 14816
rect 25044 14773 25053 14807
rect 25053 14773 25087 14807
rect 25087 14773 25096 14807
rect 25044 14764 25096 14773
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 20982 14662 21034 14714
rect 21046 14662 21098 14714
rect 21110 14662 21162 14714
rect 21174 14662 21226 14714
rect 1400 14560 1452 14612
rect 1676 14492 1728 14544
rect 4896 14560 4948 14612
rect 18512 14560 18564 14612
rect 19892 14603 19944 14612
rect 19892 14569 19901 14603
rect 19901 14569 19935 14603
rect 19935 14569 19944 14603
rect 19892 14560 19944 14569
rect 25044 14560 25096 14612
rect 4252 14492 4304 14544
rect 11704 14535 11756 14544
rect 11704 14501 11713 14535
rect 11713 14501 11747 14535
rect 11747 14501 11756 14535
rect 11704 14492 11756 14501
rect 15384 14492 15436 14544
rect 16672 14492 16724 14544
rect 18972 14492 19024 14544
rect 20444 14492 20496 14544
rect 23112 14492 23164 14544
rect 24860 14492 24912 14544
rect 25412 14492 25464 14544
rect 5172 14467 5224 14476
rect 5172 14433 5181 14467
rect 5181 14433 5215 14467
rect 5215 14433 5224 14467
rect 5172 14424 5224 14433
rect 5448 14467 5500 14476
rect 5448 14433 5482 14467
rect 5482 14433 5500 14467
rect 5448 14424 5500 14433
rect 7840 14424 7892 14476
rect 11060 14424 11112 14476
rect 11612 14467 11664 14476
rect 11612 14433 11621 14467
rect 11621 14433 11655 14467
rect 11655 14433 11664 14467
rect 11612 14424 11664 14433
rect 15292 14467 15344 14476
rect 15292 14433 15301 14467
rect 15301 14433 15335 14467
rect 15335 14433 15344 14467
rect 15292 14424 15344 14433
rect 17776 14424 17828 14476
rect 18696 14467 18748 14476
rect 18696 14433 18705 14467
rect 18705 14433 18739 14467
rect 18739 14433 18748 14467
rect 18696 14424 18748 14433
rect 20536 14424 20588 14476
rect 21732 14424 21784 14476
rect 22560 14424 22612 14476
rect 1400 14356 1452 14408
rect 7472 14356 7524 14408
rect 8208 14399 8260 14408
rect 8208 14365 8217 14399
rect 8217 14365 8251 14399
rect 8251 14365 8260 14399
rect 8208 14356 8260 14365
rect 11336 14356 11388 14408
rect 12808 14399 12860 14408
rect 12808 14365 12817 14399
rect 12817 14365 12851 14399
rect 12851 14365 12860 14399
rect 12808 14356 12860 14365
rect 18512 14356 18564 14408
rect 18880 14399 18932 14408
rect 18880 14365 18889 14399
rect 18889 14365 18923 14399
rect 18923 14365 18932 14399
rect 18880 14356 18932 14365
rect 11152 14288 11204 14340
rect 2872 14263 2924 14272
rect 2872 14229 2881 14263
rect 2881 14229 2915 14263
rect 2915 14229 2924 14263
rect 2872 14220 2924 14229
rect 4344 14263 4396 14272
rect 4344 14229 4353 14263
rect 4353 14229 4387 14263
rect 4387 14229 4396 14263
rect 4344 14220 4396 14229
rect 8024 14220 8076 14272
rect 9220 14263 9272 14272
rect 9220 14229 9229 14263
rect 9229 14229 9263 14263
rect 9263 14229 9272 14263
rect 9220 14220 9272 14229
rect 14280 14263 14332 14272
rect 14280 14229 14289 14263
rect 14289 14229 14323 14263
rect 14323 14229 14332 14263
rect 14280 14220 14332 14229
rect 16672 14263 16724 14272
rect 16672 14229 16681 14263
rect 16681 14229 16715 14263
rect 16715 14229 16724 14263
rect 16672 14220 16724 14229
rect 23848 14263 23900 14272
rect 23848 14229 23857 14263
rect 23857 14229 23891 14263
rect 23891 14229 23900 14263
rect 23848 14220 23900 14229
rect 5982 14118 6034 14170
rect 6046 14118 6098 14170
rect 6110 14118 6162 14170
rect 6174 14118 6226 14170
rect 15982 14118 16034 14170
rect 16046 14118 16098 14170
rect 16110 14118 16162 14170
rect 16174 14118 16226 14170
rect 25982 14118 26034 14170
rect 26046 14118 26098 14170
rect 26110 14118 26162 14170
rect 26174 14118 26226 14170
rect 4068 14059 4120 14068
rect 4068 14025 4077 14059
rect 4077 14025 4111 14059
rect 4111 14025 4120 14059
rect 4068 14016 4120 14025
rect 4252 14016 4304 14068
rect 5172 14016 5224 14068
rect 8944 14016 8996 14068
rect 9588 14016 9640 14068
rect 5448 13948 5500 14000
rect 9036 13948 9088 14000
rect 2320 13923 2372 13932
rect 2320 13889 2329 13923
rect 2329 13889 2363 13923
rect 2363 13889 2372 13923
rect 2320 13880 2372 13889
rect 3516 13880 3568 13932
rect 4804 13923 4856 13932
rect 4804 13889 4813 13923
rect 4813 13889 4847 13923
rect 4847 13889 4856 13923
rect 4804 13880 4856 13889
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 8024 13923 8076 13932
rect 8024 13889 8033 13923
rect 8033 13889 8067 13923
rect 8067 13889 8076 13923
rect 8024 13880 8076 13889
rect 9680 13923 9732 13932
rect 9680 13889 9689 13923
rect 9689 13889 9723 13923
rect 9723 13889 9732 13923
rect 11612 14016 11664 14068
rect 15384 14059 15436 14068
rect 15384 14025 15393 14059
rect 15393 14025 15427 14059
rect 15427 14025 15436 14059
rect 15384 14016 15436 14025
rect 16764 14016 16816 14068
rect 17776 14059 17828 14068
rect 17776 14025 17785 14059
rect 17785 14025 17819 14059
rect 17819 14025 17828 14059
rect 17776 14016 17828 14025
rect 18880 14016 18932 14068
rect 20720 14016 20772 14068
rect 23112 14059 23164 14068
rect 12532 13948 12584 14000
rect 9680 13880 9732 13889
rect 12440 13880 12492 13932
rect 15016 13948 15068 14000
rect 15292 13948 15344 14000
rect 12992 13923 13044 13932
rect 12992 13889 13001 13923
rect 13001 13889 13035 13923
rect 13035 13889 13044 13923
rect 12992 13880 13044 13889
rect 14924 13923 14976 13932
rect 14924 13889 14933 13923
rect 14933 13889 14967 13923
rect 14967 13889 14976 13923
rect 14924 13880 14976 13889
rect 18236 13923 18288 13932
rect 18236 13889 18245 13923
rect 18245 13889 18279 13923
rect 18279 13889 18288 13923
rect 18236 13880 18288 13889
rect 756 13812 808 13864
rect 2688 13812 2740 13864
rect 4068 13812 4120 13864
rect 5172 13812 5224 13864
rect 7012 13812 7064 13864
rect 7840 13812 7892 13864
rect 1676 13744 1728 13796
rect 2320 13744 2372 13796
rect 4344 13744 4396 13796
rect 8576 13744 8628 13796
rect 9220 13812 9272 13864
rect 9772 13812 9824 13864
rect 11152 13855 11204 13864
rect 2044 13676 2096 13728
rect 2504 13676 2556 13728
rect 4252 13719 4304 13728
rect 4252 13685 4261 13719
rect 4261 13685 4295 13719
rect 4295 13685 4304 13719
rect 4252 13676 4304 13685
rect 7012 13676 7064 13728
rect 8116 13676 8168 13728
rect 11152 13821 11161 13855
rect 11161 13821 11195 13855
rect 11195 13821 11204 13855
rect 11152 13812 11204 13821
rect 11612 13744 11664 13796
rect 12808 13787 12860 13796
rect 12808 13753 12817 13787
rect 12817 13753 12851 13787
rect 12851 13753 12860 13787
rect 12808 13744 12860 13753
rect 13636 13744 13688 13796
rect 14280 13812 14332 13864
rect 20536 13812 20588 13864
rect 23112 14025 23121 14059
rect 23121 14025 23155 14059
rect 23155 14025 23164 14059
rect 23112 14016 23164 14025
rect 25228 14016 25280 14068
rect 23848 13880 23900 13932
rect 24032 13812 24084 13864
rect 26148 13855 26200 13864
rect 26148 13821 26157 13855
rect 26157 13821 26191 13855
rect 26191 13821 26200 13855
rect 26148 13812 26200 13821
rect 14648 13787 14700 13796
rect 14648 13753 14657 13787
rect 14657 13753 14691 13787
rect 14691 13753 14700 13787
rect 14648 13744 14700 13753
rect 17868 13744 17920 13796
rect 22100 13676 22152 13728
rect 23480 13719 23532 13728
rect 23480 13685 23489 13719
rect 23489 13685 23523 13719
rect 23523 13685 23532 13719
rect 23480 13676 23532 13685
rect 23664 13719 23716 13728
rect 23664 13685 23673 13719
rect 23673 13685 23707 13719
rect 23707 13685 23716 13719
rect 23664 13676 23716 13685
rect 26056 13719 26108 13728
rect 26056 13685 26065 13719
rect 26065 13685 26099 13719
rect 26099 13685 26108 13719
rect 26056 13676 26108 13685
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 20982 13574 21034 13626
rect 21046 13574 21098 13626
rect 21110 13574 21162 13626
rect 21174 13574 21226 13626
rect 1676 13515 1728 13524
rect 1676 13481 1685 13515
rect 1685 13481 1719 13515
rect 1719 13481 1728 13515
rect 1676 13472 1728 13481
rect 1860 13472 1912 13524
rect 2044 13472 2096 13524
rect 6828 13515 6880 13524
rect 6828 13481 6837 13515
rect 6837 13481 6871 13515
rect 6871 13481 6880 13515
rect 6828 13472 6880 13481
rect 7012 13472 7064 13524
rect 8208 13472 8260 13524
rect 9036 13472 9088 13524
rect 9220 13472 9272 13524
rect 10876 13515 10928 13524
rect 10876 13481 10885 13515
rect 10885 13481 10919 13515
rect 10919 13481 10928 13515
rect 10876 13472 10928 13481
rect 11336 13515 11388 13524
rect 11336 13481 11345 13515
rect 11345 13481 11379 13515
rect 11379 13481 11388 13515
rect 11336 13472 11388 13481
rect 11704 13515 11756 13524
rect 11704 13481 11713 13515
rect 11713 13481 11747 13515
rect 11747 13481 11756 13515
rect 11704 13472 11756 13481
rect 12164 13515 12216 13524
rect 12164 13481 12173 13515
rect 12173 13481 12207 13515
rect 12207 13481 12216 13515
rect 12164 13472 12216 13481
rect 13636 13515 13688 13524
rect 13636 13481 13645 13515
rect 13645 13481 13679 13515
rect 13679 13481 13688 13515
rect 13636 13472 13688 13481
rect 14648 13472 14700 13524
rect 16304 13472 16356 13524
rect 18880 13472 18932 13524
rect 22560 13515 22612 13524
rect 22560 13481 22569 13515
rect 22569 13481 22603 13515
rect 22603 13481 22612 13515
rect 22560 13472 22612 13481
rect 24032 13515 24084 13524
rect 24032 13481 24041 13515
rect 24041 13481 24075 13515
rect 24075 13481 24084 13515
rect 24032 13472 24084 13481
rect 25044 13472 25096 13524
rect 26240 13515 26292 13524
rect 26240 13481 26249 13515
rect 26249 13481 26283 13515
rect 26283 13481 26292 13515
rect 26240 13472 26292 13481
rect 26424 13472 26476 13524
rect 4712 13447 4764 13456
rect 4712 13413 4721 13447
rect 4721 13413 4755 13447
rect 4755 13413 4764 13447
rect 4712 13404 4764 13413
rect 12072 13447 12124 13456
rect 12072 13413 12081 13447
rect 12081 13413 12115 13447
rect 12115 13413 12124 13447
rect 12072 13404 12124 13413
rect 15384 13404 15436 13456
rect 15844 13404 15896 13456
rect 1676 13336 1728 13388
rect 1860 13336 1912 13388
rect 5080 13336 5132 13388
rect 8392 13379 8444 13388
rect 8392 13345 8401 13379
rect 8401 13345 8435 13379
rect 8435 13345 8444 13379
rect 8392 13336 8444 13345
rect 2596 13268 2648 13320
rect 2872 13268 2924 13320
rect 4804 13311 4856 13320
rect 4804 13277 4813 13311
rect 4813 13277 4847 13311
rect 4847 13277 4856 13311
rect 4804 13268 4856 13277
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 7932 13200 7984 13252
rect 9680 13200 9732 13252
rect 13636 13336 13688 13388
rect 14004 13379 14056 13388
rect 14004 13345 14013 13379
rect 14013 13345 14047 13379
rect 14047 13345 14056 13379
rect 14004 13336 14056 13345
rect 11612 13268 11664 13320
rect 12992 13268 13044 13320
rect 13728 13268 13780 13320
rect 15200 13268 15252 13320
rect 17960 13404 18012 13456
rect 18236 13404 18288 13456
rect 23664 13404 23716 13456
rect 25228 13379 25280 13388
rect 25228 13345 25237 13379
rect 25237 13345 25271 13379
rect 25271 13345 25280 13379
rect 25228 13336 25280 13345
rect 25320 13268 25372 13320
rect 26056 13268 26108 13320
rect 26516 13268 26568 13320
rect 10416 13200 10468 13252
rect 10784 13200 10836 13252
rect 19156 13200 19208 13252
rect 2412 13132 2464 13184
rect 4068 13132 4120 13184
rect 4344 13132 4396 13184
rect 4528 13132 4580 13184
rect 18512 13132 18564 13184
rect 22100 13175 22152 13184
rect 22100 13141 22109 13175
rect 22109 13141 22143 13175
rect 22143 13141 22152 13175
rect 22100 13132 22152 13141
rect 23848 13132 23900 13184
rect 24676 13132 24728 13184
rect 25504 13132 25556 13184
rect 5982 13030 6034 13082
rect 6046 13030 6098 13082
rect 6110 13030 6162 13082
rect 6174 13030 6226 13082
rect 15982 13030 16034 13082
rect 16046 13030 16098 13082
rect 16110 13030 16162 13082
rect 16174 13030 16226 13082
rect 25982 13030 26034 13082
rect 26046 13030 26098 13082
rect 26110 13030 26162 13082
rect 26174 13030 26226 13082
rect 3516 12971 3568 12980
rect 3516 12937 3525 12971
rect 3525 12937 3559 12971
rect 3559 12937 3568 12971
rect 3516 12928 3568 12937
rect 4712 12971 4764 12980
rect 4712 12937 4721 12971
rect 4721 12937 4755 12971
rect 4755 12937 4764 12971
rect 4712 12928 4764 12937
rect 8392 12928 8444 12980
rect 8852 12928 8904 12980
rect 10416 12971 10468 12980
rect 10416 12937 10425 12971
rect 10425 12937 10459 12971
rect 10459 12937 10468 12971
rect 10416 12928 10468 12937
rect 11612 12928 11664 12980
rect 12164 12971 12216 12980
rect 12164 12937 12173 12971
rect 12173 12937 12207 12971
rect 12207 12937 12216 12971
rect 12164 12928 12216 12937
rect 13636 12971 13688 12980
rect 13636 12937 13645 12971
rect 13645 12937 13679 12971
rect 13679 12937 13688 12971
rect 13636 12928 13688 12937
rect 15844 12928 15896 12980
rect 17868 12971 17920 12980
rect 17868 12937 17877 12971
rect 17877 12937 17911 12971
rect 17911 12937 17920 12971
rect 17868 12928 17920 12937
rect 23664 12928 23716 12980
rect 25228 12928 25280 12980
rect 5080 12903 5132 12912
rect 5080 12869 5089 12903
rect 5089 12869 5123 12903
rect 5123 12869 5132 12903
rect 5080 12860 5132 12869
rect 12072 12860 12124 12912
rect 14280 12903 14332 12912
rect 14280 12869 14289 12903
rect 14289 12869 14323 12903
rect 14323 12869 14332 12903
rect 14280 12860 14332 12869
rect 3148 12792 3200 12844
rect 3516 12792 3568 12844
rect 6828 12835 6880 12844
rect 6828 12801 6837 12835
rect 6837 12801 6871 12835
rect 6871 12801 6880 12835
rect 6828 12792 6880 12801
rect 10140 12835 10192 12844
rect 10140 12801 10149 12835
rect 10149 12801 10183 12835
rect 10183 12801 10192 12835
rect 16304 12860 16356 12912
rect 14924 12835 14976 12844
rect 10140 12792 10192 12801
rect 14924 12801 14933 12835
rect 14933 12801 14967 12835
rect 14967 12801 14976 12835
rect 14924 12792 14976 12801
rect 25320 12860 25372 12912
rect 18604 12835 18656 12844
rect 18604 12801 18613 12835
rect 18613 12801 18647 12835
rect 18647 12801 18656 12835
rect 18604 12792 18656 12801
rect 20444 12835 20496 12844
rect 20444 12801 20453 12835
rect 20453 12801 20487 12835
rect 20487 12801 20496 12835
rect 20444 12792 20496 12801
rect 26056 12835 26108 12844
rect 26056 12801 26065 12835
rect 26065 12801 26099 12835
rect 26099 12801 26108 12835
rect 26056 12792 26108 12801
rect 2412 12767 2464 12776
rect 2412 12733 2421 12767
rect 2421 12733 2455 12767
rect 2455 12733 2464 12767
rect 2412 12724 2464 12733
rect 4068 12767 4120 12776
rect 4068 12733 4077 12767
rect 4077 12733 4111 12767
rect 4111 12733 4120 12767
rect 4068 12724 4120 12733
rect 10048 12724 10100 12776
rect 14004 12724 14056 12776
rect 25044 12767 25096 12776
rect 25044 12733 25053 12767
rect 25053 12733 25087 12767
rect 25087 12733 25096 12767
rect 25044 12724 25096 12733
rect 25780 12724 25832 12776
rect 4252 12656 4304 12708
rect 6736 12656 6788 12708
rect 16764 12656 16816 12708
rect 20812 12656 20864 12708
rect 21732 12656 21784 12708
rect 25320 12699 25372 12708
rect 25320 12665 25329 12699
rect 25329 12665 25363 12699
rect 25363 12665 25372 12699
rect 25320 12656 25372 12665
rect 1860 12631 1912 12640
rect 1860 12597 1869 12631
rect 1869 12597 1903 12631
rect 1903 12597 1912 12631
rect 1860 12588 1912 12597
rect 2044 12631 2096 12640
rect 2044 12597 2053 12631
rect 2053 12597 2087 12631
rect 2087 12597 2096 12631
rect 2044 12588 2096 12597
rect 3608 12631 3660 12640
rect 3608 12597 3617 12631
rect 3617 12597 3651 12631
rect 3651 12597 3660 12631
rect 3608 12588 3660 12597
rect 8208 12631 8260 12640
rect 8208 12597 8217 12631
rect 8217 12597 8251 12631
rect 8251 12597 8260 12631
rect 8208 12588 8260 12597
rect 9680 12631 9732 12640
rect 9680 12597 9689 12631
rect 9689 12597 9723 12631
rect 9723 12597 9732 12631
rect 9680 12588 9732 12597
rect 14648 12631 14700 12640
rect 14648 12597 14657 12631
rect 14657 12597 14691 12631
rect 14691 12597 14700 12631
rect 14648 12588 14700 12597
rect 14740 12631 14792 12640
rect 14740 12597 14749 12631
rect 14749 12597 14783 12631
rect 14783 12597 14792 12631
rect 14740 12588 14792 12597
rect 15200 12588 15252 12640
rect 15476 12588 15528 12640
rect 18052 12631 18104 12640
rect 18052 12597 18061 12631
rect 18061 12597 18095 12631
rect 18095 12597 18104 12631
rect 18052 12588 18104 12597
rect 19156 12631 19208 12640
rect 19156 12597 19165 12631
rect 19165 12597 19199 12631
rect 19199 12597 19208 12631
rect 19156 12588 19208 12597
rect 21548 12588 21600 12640
rect 24860 12588 24912 12640
rect 25044 12588 25096 12640
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 20982 12486 21034 12538
rect 21046 12486 21098 12538
rect 21110 12486 21162 12538
rect 21174 12486 21226 12538
rect 3608 12384 3660 12436
rect 4068 12384 4120 12436
rect 4344 12384 4396 12436
rect 13728 12427 13780 12436
rect 13728 12393 13737 12427
rect 13737 12393 13771 12427
rect 13771 12393 13780 12427
rect 13728 12384 13780 12393
rect 18604 12384 18656 12436
rect 20444 12427 20496 12436
rect 20444 12393 20453 12427
rect 20453 12393 20487 12427
rect 20487 12393 20496 12427
rect 20444 12384 20496 12393
rect 20720 12384 20772 12436
rect 24768 12384 24820 12436
rect 24952 12384 25004 12436
rect 26516 12384 26568 12436
rect 26700 12384 26752 12436
rect 26976 12427 27028 12436
rect 26976 12393 26985 12427
rect 26985 12393 27019 12427
rect 27019 12393 27028 12427
rect 26976 12384 27028 12393
rect 2688 12316 2740 12368
rect 2872 12316 2924 12368
rect 17960 12316 18012 12368
rect 24308 12316 24360 12368
rect 24492 12316 24544 12368
rect 24584 12316 24636 12368
rect 25412 12316 25464 12368
rect 26424 12316 26476 12368
rect 2320 12291 2372 12300
rect 2320 12257 2329 12291
rect 2329 12257 2363 12291
rect 2363 12257 2372 12291
rect 2320 12248 2372 12257
rect 2964 12248 3016 12300
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 3516 12180 3568 12232
rect 10600 12291 10652 12300
rect 10600 12257 10609 12291
rect 10609 12257 10643 12291
rect 10643 12257 10652 12291
rect 10600 12248 10652 12257
rect 15660 12291 15712 12300
rect 15660 12257 15669 12291
rect 15669 12257 15703 12291
rect 15703 12257 15712 12291
rect 15660 12248 15712 12257
rect 17868 12248 17920 12300
rect 21640 12248 21692 12300
rect 25228 12291 25280 12300
rect 25228 12257 25237 12291
rect 25237 12257 25271 12291
rect 25271 12257 25280 12291
rect 25228 12248 25280 12257
rect 25596 12248 25648 12300
rect 26516 12248 26568 12300
rect 4252 12223 4304 12232
rect 4252 12189 4261 12223
rect 4261 12189 4295 12223
rect 4295 12189 4304 12223
rect 4252 12180 4304 12189
rect 10416 12180 10468 12232
rect 10784 12223 10836 12232
rect 10784 12189 10793 12223
rect 10793 12189 10827 12223
rect 10827 12189 10836 12223
rect 10784 12180 10836 12189
rect 15844 12180 15896 12232
rect 15936 12223 15988 12232
rect 15936 12189 15945 12223
rect 15945 12189 15979 12223
rect 15979 12189 15988 12223
rect 15936 12180 15988 12189
rect 16672 12180 16724 12232
rect 21364 12223 21416 12232
rect 21364 12189 21373 12223
rect 21373 12189 21407 12223
rect 21407 12189 21416 12223
rect 21364 12180 21416 12189
rect 21548 12223 21600 12232
rect 21548 12189 21557 12223
rect 21557 12189 21591 12223
rect 21591 12189 21600 12223
rect 21548 12180 21600 12189
rect 22468 12223 22520 12232
rect 22468 12189 22477 12223
rect 22477 12189 22511 12223
rect 22511 12189 22520 12223
rect 22468 12180 22520 12189
rect 23940 12180 23992 12232
rect 24492 12180 24544 12232
rect 27068 12223 27120 12232
rect 5632 12155 5684 12164
rect 5632 12121 5641 12155
rect 5641 12121 5675 12155
rect 5675 12121 5684 12155
rect 5632 12112 5684 12121
rect 14740 12155 14792 12164
rect 14740 12121 14749 12155
rect 14749 12121 14783 12155
rect 14783 12121 14792 12155
rect 14740 12112 14792 12121
rect 23848 12112 23900 12164
rect 24768 12155 24820 12164
rect 24768 12121 24777 12155
rect 24777 12121 24811 12155
rect 24811 12121 24820 12155
rect 27068 12189 27077 12223
rect 27077 12189 27111 12223
rect 27111 12189 27120 12223
rect 27068 12180 27120 12189
rect 24768 12112 24820 12121
rect 26056 12112 26108 12164
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 6920 12087 6972 12096
rect 6920 12053 6929 12087
rect 6929 12053 6963 12087
rect 6963 12053 6972 12087
rect 6920 12044 6972 12053
rect 10324 12044 10376 12096
rect 12716 12044 12768 12096
rect 14924 12044 14976 12096
rect 15384 12044 15436 12096
rect 16304 12087 16356 12096
rect 16304 12053 16313 12087
rect 16313 12053 16347 12087
rect 16347 12053 16356 12087
rect 16304 12044 16356 12053
rect 24216 12087 24268 12096
rect 24216 12053 24225 12087
rect 24225 12053 24259 12087
rect 24259 12053 24268 12087
rect 24216 12044 24268 12053
rect 24860 12087 24912 12096
rect 24860 12053 24869 12087
rect 24869 12053 24903 12087
rect 24903 12053 24912 12087
rect 24860 12044 24912 12053
rect 27160 12044 27212 12096
rect 27528 12087 27580 12096
rect 27528 12053 27537 12087
rect 27537 12053 27571 12087
rect 27571 12053 27580 12087
rect 27528 12044 27580 12053
rect 5982 11942 6034 11994
rect 6046 11942 6098 11994
rect 6110 11942 6162 11994
rect 6174 11942 6226 11994
rect 15982 11942 16034 11994
rect 16046 11942 16098 11994
rect 16110 11942 16162 11994
rect 16174 11942 16226 11994
rect 25982 11942 26034 11994
rect 26046 11942 26098 11994
rect 26110 11942 26162 11994
rect 26174 11942 26226 11994
rect 2320 11840 2372 11892
rect 2596 11840 2648 11892
rect 3976 11883 4028 11892
rect 3976 11849 3985 11883
rect 3985 11849 4019 11883
rect 4019 11849 4028 11883
rect 3976 11840 4028 11849
rect 4252 11840 4304 11892
rect 5448 11840 5500 11892
rect 10600 11840 10652 11892
rect 15108 11883 15160 11892
rect 3148 11704 3200 11756
rect 4436 11747 4488 11756
rect 4436 11713 4445 11747
rect 4445 11713 4479 11747
rect 4479 11713 4488 11747
rect 4436 11704 4488 11713
rect 6920 11704 6972 11756
rect 8208 11772 8260 11824
rect 8484 11747 8536 11756
rect 8484 11713 8493 11747
rect 8493 11713 8527 11747
rect 8527 11713 8536 11747
rect 8484 11704 8536 11713
rect 15108 11849 15117 11883
rect 15117 11849 15151 11883
rect 15151 11849 15160 11883
rect 15108 11840 15160 11849
rect 16672 11883 16724 11892
rect 16672 11849 16681 11883
rect 16681 11849 16715 11883
rect 16715 11849 16724 11883
rect 16672 11840 16724 11849
rect 21364 11840 21416 11892
rect 25228 11840 25280 11892
rect 26332 11840 26384 11892
rect 14924 11772 14976 11824
rect 17408 11772 17460 11824
rect 17960 11772 18012 11824
rect 21548 11772 21600 11824
rect 13636 11747 13688 11756
rect 13636 11713 13645 11747
rect 13645 11713 13679 11747
rect 13679 11713 13688 11747
rect 13636 11704 13688 11713
rect 3976 11636 4028 11688
rect 15016 11704 15068 11756
rect 16120 11747 16172 11756
rect 16120 11713 16129 11747
rect 16129 11713 16163 11747
rect 16163 11713 16172 11747
rect 16120 11704 16172 11713
rect 16304 11747 16356 11756
rect 16304 11713 16313 11747
rect 16313 11713 16347 11747
rect 16347 11713 16356 11747
rect 16304 11704 16356 11713
rect 19156 11704 19208 11756
rect 20812 11704 20864 11756
rect 22284 11704 22336 11756
rect 26424 11772 26476 11824
rect 26700 11704 26752 11756
rect 27160 11747 27212 11756
rect 27160 11713 27169 11747
rect 27169 11713 27203 11747
rect 27203 11713 27212 11747
rect 27160 11704 27212 11713
rect 14280 11636 14332 11688
rect 21272 11679 21324 11688
rect 21272 11645 21281 11679
rect 21281 11645 21315 11679
rect 21315 11645 21324 11679
rect 21272 11636 21324 11645
rect 23848 11636 23900 11688
rect 24216 11679 24268 11688
rect 24216 11645 24225 11679
rect 24225 11645 24259 11679
rect 24259 11645 24268 11679
rect 24216 11636 24268 11645
rect 24768 11636 24820 11688
rect 24860 11636 24912 11688
rect 27528 11636 27580 11688
rect 18144 11568 18196 11620
rect 19064 11568 19116 11620
rect 21640 11568 21692 11620
rect 25780 11568 25832 11620
rect 27252 11568 27304 11620
rect 1768 11543 1820 11552
rect 1768 11509 1777 11543
rect 1777 11509 1811 11543
rect 1811 11509 1820 11543
rect 1768 11500 1820 11509
rect 1952 11500 2004 11552
rect 2136 11543 2188 11552
rect 2136 11509 2145 11543
rect 2145 11509 2179 11543
rect 2179 11509 2188 11543
rect 2136 11500 2188 11509
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 2964 11500 3016 11552
rect 3516 11543 3568 11552
rect 3516 11509 3525 11543
rect 3525 11509 3559 11543
rect 3559 11509 3568 11543
rect 3516 11500 3568 11509
rect 6828 11543 6880 11552
rect 6828 11509 6837 11543
rect 6837 11509 6871 11543
rect 6871 11509 6880 11543
rect 6828 11500 6880 11509
rect 7196 11543 7248 11552
rect 7196 11509 7205 11543
rect 7205 11509 7239 11543
rect 7239 11509 7248 11543
rect 7196 11500 7248 11509
rect 8300 11543 8352 11552
rect 8300 11509 8309 11543
rect 8309 11509 8343 11543
rect 8343 11509 8352 11543
rect 8300 11500 8352 11509
rect 9588 11500 9640 11552
rect 10416 11543 10468 11552
rect 10416 11509 10425 11543
rect 10425 11509 10459 11543
rect 10459 11509 10468 11543
rect 10416 11500 10468 11509
rect 15200 11500 15252 11552
rect 18420 11543 18472 11552
rect 18420 11509 18429 11543
rect 18429 11509 18463 11543
rect 18463 11509 18472 11543
rect 18420 11500 18472 11509
rect 18880 11543 18932 11552
rect 18880 11509 18889 11543
rect 18889 11509 18923 11543
rect 18923 11509 18932 11543
rect 18880 11500 18932 11509
rect 21456 11500 21508 11552
rect 22008 11500 22060 11552
rect 26516 11543 26568 11552
rect 26516 11509 26525 11543
rect 26525 11509 26559 11543
rect 26559 11509 26568 11543
rect 26516 11500 26568 11509
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 20982 11398 21034 11450
rect 21046 11398 21098 11450
rect 21110 11398 21162 11450
rect 21174 11398 21226 11450
rect 2228 11296 2280 11348
rect 6920 11296 6972 11348
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 9680 11339 9732 11348
rect 9680 11305 9689 11339
rect 9689 11305 9723 11339
rect 9723 11305 9732 11339
rect 9680 11296 9732 11305
rect 16120 11296 16172 11348
rect 16764 11339 16816 11348
rect 16764 11305 16773 11339
rect 16773 11305 16807 11339
rect 16807 11305 16816 11339
rect 16764 11296 16816 11305
rect 17868 11339 17920 11348
rect 17868 11305 17877 11339
rect 17877 11305 17911 11339
rect 17911 11305 17920 11339
rect 17868 11296 17920 11305
rect 21364 11296 21416 11348
rect 21640 11339 21692 11348
rect 21640 11305 21649 11339
rect 21649 11305 21683 11339
rect 21683 11305 21692 11339
rect 21640 11296 21692 11305
rect 22100 11296 22152 11348
rect 22468 11296 22520 11348
rect 24768 11296 24820 11348
rect 1400 11228 1452 11280
rect 2964 11228 3016 11280
rect 3148 11228 3200 11280
rect 17224 11228 17276 11280
rect 18420 11228 18472 11280
rect 2228 11160 2280 11212
rect 2688 11160 2740 11212
rect 6920 11203 6972 11212
rect 6920 11169 6929 11203
rect 6929 11169 6963 11203
rect 6963 11169 6972 11203
rect 6920 11160 6972 11169
rect 10324 11160 10376 11212
rect 10968 11160 11020 11212
rect 12716 11203 12768 11212
rect 12716 11169 12750 11203
rect 12750 11169 12768 11203
rect 12716 11160 12768 11169
rect 15660 11160 15712 11212
rect 17960 11160 18012 11212
rect 18696 11203 18748 11212
rect 18696 11169 18705 11203
rect 18705 11169 18739 11203
rect 18739 11169 18748 11203
rect 18696 11160 18748 11169
rect 21732 11160 21784 11212
rect 25688 11296 25740 11348
rect 26700 11339 26752 11348
rect 26700 11305 26709 11339
rect 26709 11305 26743 11339
rect 26743 11305 26752 11339
rect 26700 11296 26752 11305
rect 27068 11339 27120 11348
rect 27068 11305 27077 11339
rect 27077 11305 27111 11339
rect 27111 11305 27120 11339
rect 27068 11296 27120 11305
rect 27160 11296 27212 11348
rect 27620 11339 27672 11348
rect 27620 11305 27629 11339
rect 27629 11305 27663 11339
rect 27663 11305 27672 11339
rect 27620 11296 27672 11305
rect 25504 11228 25556 11280
rect 25596 11228 25648 11280
rect 27344 11228 27396 11280
rect 25320 11203 25372 11212
rect 25320 11169 25329 11203
rect 25329 11169 25363 11203
rect 25363 11169 25372 11203
rect 25320 11160 25372 11169
rect 26516 11203 26568 11212
rect 26516 11169 26525 11203
rect 26525 11169 26559 11203
rect 26559 11169 26568 11203
rect 26516 11160 26568 11169
rect 2504 11135 2556 11144
rect 2504 11101 2513 11135
rect 2513 11101 2547 11135
rect 2547 11101 2556 11135
rect 7012 11135 7064 11144
rect 2504 11092 2556 11101
rect 7012 11101 7021 11135
rect 7021 11101 7055 11135
rect 7055 11101 7064 11135
rect 7012 11092 7064 11101
rect 10140 11135 10192 11144
rect 2780 11024 2832 11076
rect 6736 11024 6788 11076
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 9680 11024 9732 11076
rect 12440 11135 12492 11144
rect 12440 11101 12449 11135
rect 12449 11101 12483 11135
rect 12483 11101 12492 11135
rect 15292 11135 15344 11144
rect 12440 11092 12492 11101
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 17408 11135 17460 11144
rect 15844 11067 15896 11076
rect 15844 11033 15853 11067
rect 15853 11033 15887 11067
rect 15887 11033 15896 11067
rect 15844 11024 15896 11033
rect 16856 11024 16908 11076
rect 17408 11101 17417 11135
rect 17417 11101 17451 11135
rect 17451 11101 17460 11135
rect 17408 11092 17460 11101
rect 18788 11135 18840 11144
rect 18788 11101 18797 11135
rect 18797 11101 18831 11135
rect 18831 11101 18840 11135
rect 18788 11092 18840 11101
rect 18420 11024 18472 11076
rect 19156 11092 19208 11144
rect 22284 11135 22336 11144
rect 22284 11101 22293 11135
rect 22293 11101 22327 11135
rect 22327 11101 22336 11135
rect 22284 11092 22336 11101
rect 22468 11092 22520 11144
rect 19432 11067 19484 11076
rect 19432 11033 19441 11067
rect 19441 11033 19475 11067
rect 19475 11033 19484 11067
rect 19432 11024 19484 11033
rect 21456 11067 21508 11076
rect 21456 11033 21465 11067
rect 21465 11033 21499 11067
rect 21499 11033 21508 11067
rect 21456 11024 21508 11033
rect 25504 11067 25556 11076
rect 25504 11033 25513 11067
rect 25513 11033 25547 11067
rect 25547 11033 25556 11067
rect 25504 11024 25556 11033
rect 7840 10956 7892 11008
rect 10692 10999 10744 11008
rect 10692 10965 10701 10999
rect 10701 10965 10735 10999
rect 10735 10965 10744 10999
rect 10692 10956 10744 10965
rect 13544 10956 13596 11008
rect 14188 10956 14240 11008
rect 14464 10999 14516 11008
rect 14464 10965 14473 10999
rect 14473 10965 14507 10999
rect 14507 10965 14516 10999
rect 14464 10956 14516 10965
rect 5982 10854 6034 10906
rect 6046 10854 6098 10906
rect 6110 10854 6162 10906
rect 6174 10854 6226 10906
rect 15982 10854 16034 10906
rect 16046 10854 16098 10906
rect 16110 10854 16162 10906
rect 16174 10854 16226 10906
rect 25982 10854 26034 10906
rect 26046 10854 26098 10906
rect 26110 10854 26162 10906
rect 26174 10854 26226 10906
rect 2228 10752 2280 10804
rect 2320 10752 2372 10804
rect 2780 10752 2832 10804
rect 6920 10752 6972 10804
rect 10140 10752 10192 10804
rect 11060 10795 11112 10804
rect 11060 10761 11069 10795
rect 11069 10761 11103 10795
rect 11103 10761 11112 10795
rect 11060 10752 11112 10761
rect 12716 10795 12768 10804
rect 12716 10761 12725 10795
rect 12725 10761 12759 10795
rect 12759 10761 12768 10795
rect 12716 10752 12768 10761
rect 14188 10795 14240 10804
rect 14188 10761 14197 10795
rect 14197 10761 14231 10795
rect 14231 10761 14240 10795
rect 14188 10752 14240 10761
rect 14924 10752 14976 10804
rect 15292 10795 15344 10804
rect 15292 10761 15301 10795
rect 15301 10761 15335 10795
rect 15335 10761 15344 10795
rect 15292 10752 15344 10761
rect 17408 10752 17460 10804
rect 17868 10752 17920 10804
rect 18880 10795 18932 10804
rect 18880 10761 18889 10795
rect 18889 10761 18923 10795
rect 18923 10761 18932 10795
rect 18880 10752 18932 10761
rect 21732 10795 21784 10804
rect 21732 10761 21741 10795
rect 21741 10761 21775 10795
rect 21775 10761 21784 10795
rect 21732 10752 21784 10761
rect 22100 10795 22152 10804
rect 22100 10761 22109 10795
rect 22109 10761 22143 10795
rect 22143 10761 22152 10795
rect 25320 10795 25372 10804
rect 22100 10752 22152 10761
rect 25320 10761 25329 10795
rect 25329 10761 25363 10795
rect 25363 10761 25372 10795
rect 25320 10752 25372 10761
rect 26516 10752 26568 10804
rect 2504 10684 2556 10736
rect 6736 10684 6788 10736
rect 9588 10684 9640 10736
rect 13820 10684 13872 10736
rect 7564 10616 7616 10668
rect 8300 10616 8352 10668
rect 10692 10616 10744 10668
rect 11888 10616 11940 10668
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 3056 10591 3108 10600
rect 3056 10557 3065 10591
rect 3065 10557 3099 10591
rect 3099 10557 3108 10591
rect 3056 10548 3108 10557
rect 3148 10548 3200 10600
rect 7472 10591 7524 10600
rect 7472 10557 7481 10591
rect 7481 10557 7515 10591
rect 7515 10557 7524 10591
rect 7472 10548 7524 10557
rect 14464 10548 14516 10600
rect 14924 10659 14976 10668
rect 14924 10625 14933 10659
rect 14933 10625 14967 10659
rect 14967 10625 14976 10659
rect 14924 10616 14976 10625
rect 15384 10616 15436 10668
rect 16304 10616 16356 10668
rect 19432 10659 19484 10668
rect 19432 10625 19441 10659
rect 19441 10625 19475 10659
rect 19475 10625 19484 10659
rect 19432 10616 19484 10625
rect 15292 10548 15344 10600
rect 7012 10480 7064 10532
rect 10048 10480 10100 10532
rect 10600 10480 10652 10532
rect 14740 10523 14792 10532
rect 14740 10489 14749 10523
rect 14749 10489 14783 10523
rect 14783 10489 14792 10523
rect 14740 10480 14792 10489
rect 16396 10480 16448 10532
rect 18788 10480 18840 10532
rect 23848 10548 23900 10600
rect 27528 10591 27580 10600
rect 27528 10557 27537 10591
rect 27537 10557 27571 10591
rect 27571 10557 27580 10591
rect 27528 10548 27580 10557
rect 19524 10480 19576 10532
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 4436 10455 4488 10464
rect 4436 10421 4445 10455
rect 4445 10421 4479 10455
rect 4479 10421 4488 10455
rect 4436 10412 4488 10421
rect 6276 10455 6328 10464
rect 6276 10421 6285 10455
rect 6285 10421 6319 10455
rect 6319 10421 6328 10455
rect 6276 10412 6328 10421
rect 7840 10412 7892 10464
rect 9864 10455 9916 10464
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 9864 10412 9916 10421
rect 13268 10412 13320 10464
rect 19156 10412 19208 10464
rect 22468 10455 22520 10464
rect 22468 10421 22477 10455
rect 22477 10421 22511 10455
rect 22511 10421 22520 10455
rect 22468 10412 22520 10421
rect 23480 10412 23532 10464
rect 26608 10455 26660 10464
rect 26608 10421 26617 10455
rect 26617 10421 26651 10455
rect 26651 10421 26660 10455
rect 26608 10412 26660 10421
rect 27712 10455 27764 10464
rect 27712 10421 27721 10455
rect 27721 10421 27755 10455
rect 27755 10421 27764 10455
rect 27712 10412 27764 10421
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 20982 10310 21034 10362
rect 21046 10310 21098 10362
rect 21110 10310 21162 10362
rect 21174 10310 21226 10362
rect 2044 10251 2096 10260
rect 2044 10217 2053 10251
rect 2053 10217 2087 10251
rect 2087 10217 2096 10251
rect 2044 10208 2096 10217
rect 2136 10208 2188 10260
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 6736 10208 6788 10260
rect 6920 10251 6972 10260
rect 6920 10217 6929 10251
rect 6929 10217 6963 10251
rect 6963 10217 6972 10251
rect 6920 10208 6972 10217
rect 7012 10208 7064 10260
rect 11888 10251 11940 10260
rect 11888 10217 11897 10251
rect 11897 10217 11931 10251
rect 11931 10217 11940 10251
rect 11888 10208 11940 10217
rect 14740 10208 14792 10260
rect 16304 10251 16356 10260
rect 16304 10217 16313 10251
rect 16313 10217 16347 10251
rect 16347 10217 16356 10251
rect 16304 10208 16356 10217
rect 16856 10251 16908 10260
rect 16856 10217 16865 10251
rect 16865 10217 16899 10251
rect 16899 10217 16908 10251
rect 16856 10208 16908 10217
rect 17224 10251 17276 10260
rect 17224 10217 17233 10251
rect 17233 10217 17267 10251
rect 17267 10217 17276 10251
rect 17224 10208 17276 10217
rect 18420 10251 18472 10260
rect 18420 10217 18429 10251
rect 18429 10217 18463 10251
rect 18463 10217 18472 10251
rect 18420 10208 18472 10217
rect 18788 10251 18840 10260
rect 18788 10217 18797 10251
rect 18797 10217 18831 10251
rect 18831 10217 18840 10251
rect 18788 10208 18840 10217
rect 19064 10208 19116 10260
rect 22468 10208 22520 10260
rect 23480 10208 23532 10260
rect 1768 10140 1820 10192
rect 3056 10140 3108 10192
rect 3608 10140 3660 10192
rect 5540 10140 5592 10192
rect 7472 10140 7524 10192
rect 7748 10140 7800 10192
rect 10692 10140 10744 10192
rect 13636 10140 13688 10192
rect 15108 10140 15160 10192
rect 18236 10140 18288 10192
rect 24124 10140 24176 10192
rect 24860 10140 24912 10192
rect 27436 10140 27488 10192
rect 8852 10072 8904 10124
rect 13820 10115 13872 10124
rect 13820 10081 13829 10115
rect 13829 10081 13863 10115
rect 13863 10081 13872 10115
rect 13820 10072 13872 10081
rect 15660 10115 15712 10124
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 2320 10004 2372 10056
rect 7656 10047 7708 10056
rect 7656 10013 7665 10047
rect 7665 10013 7699 10047
rect 7699 10013 7708 10047
rect 7656 10004 7708 10013
rect 6276 9936 6328 9988
rect 7564 9936 7616 9988
rect 10416 10004 10468 10056
rect 14004 10047 14056 10056
rect 14004 10013 14013 10047
rect 14013 10013 14047 10047
rect 14047 10013 14056 10047
rect 14004 10004 14056 10013
rect 15568 10004 15620 10056
rect 16488 10072 16540 10124
rect 18604 10072 18656 10124
rect 18788 10072 18840 10124
rect 20536 10115 20588 10124
rect 20536 10081 20545 10115
rect 20545 10081 20579 10115
rect 20579 10081 20588 10115
rect 20536 10072 20588 10081
rect 21456 10072 21508 10124
rect 26424 10072 26476 10124
rect 16304 10004 16356 10056
rect 19432 10047 19484 10056
rect 19432 10013 19441 10047
rect 19441 10013 19475 10047
rect 19475 10013 19484 10047
rect 19432 10004 19484 10013
rect 20812 10004 20864 10056
rect 21364 10047 21416 10056
rect 21364 10013 21373 10047
rect 21373 10013 21407 10047
rect 21407 10013 21416 10047
rect 21364 10004 21416 10013
rect 24216 10004 24268 10056
rect 23296 9936 23348 9988
rect 1676 9868 1728 9920
rect 5172 9868 5224 9920
rect 8116 9868 8168 9920
rect 8392 9868 8444 9920
rect 8484 9868 8536 9920
rect 9588 9868 9640 9920
rect 10048 9911 10100 9920
rect 10048 9877 10057 9911
rect 10057 9877 10091 9911
rect 10091 9877 10100 9911
rect 10048 9868 10100 9877
rect 13268 9911 13320 9920
rect 13268 9877 13277 9911
rect 13277 9877 13311 9911
rect 13311 9877 13320 9911
rect 13268 9868 13320 9877
rect 13728 9868 13780 9920
rect 20352 9911 20404 9920
rect 20352 9877 20361 9911
rect 20361 9877 20395 9911
rect 20395 9877 20404 9911
rect 20352 9868 20404 9877
rect 24032 9868 24084 9920
rect 24400 9868 24452 9920
rect 26700 9911 26752 9920
rect 26700 9877 26709 9911
rect 26709 9877 26743 9911
rect 26743 9877 26752 9911
rect 26700 9868 26752 9877
rect 5982 9766 6034 9818
rect 6046 9766 6098 9818
rect 6110 9766 6162 9818
rect 6174 9766 6226 9818
rect 15982 9766 16034 9818
rect 16046 9766 16098 9818
rect 16110 9766 16162 9818
rect 16174 9766 16226 9818
rect 25982 9766 26034 9818
rect 26046 9766 26098 9818
rect 26110 9766 26162 9818
rect 26174 9766 26226 9818
rect 2320 9707 2372 9716
rect 2320 9673 2329 9707
rect 2329 9673 2363 9707
rect 2363 9673 2372 9707
rect 2320 9664 2372 9673
rect 3608 9707 3660 9716
rect 3608 9673 3617 9707
rect 3617 9673 3651 9707
rect 3651 9673 3660 9707
rect 3608 9664 3660 9673
rect 6276 9664 6328 9716
rect 7656 9664 7708 9716
rect 7840 9664 7892 9716
rect 2872 9596 2924 9648
rect 2964 9596 3016 9648
rect 3148 9639 3200 9648
rect 3148 9605 3157 9639
rect 3157 9605 3191 9639
rect 3191 9605 3200 9639
rect 3148 9596 3200 9605
rect 13820 9664 13872 9716
rect 15660 9664 15712 9716
rect 16304 9664 16356 9716
rect 20536 9664 20588 9716
rect 24124 9664 24176 9716
rect 26516 9664 26568 9716
rect 18696 9596 18748 9648
rect 3148 9460 3200 9512
rect 3608 9460 3660 9512
rect 7196 9528 7248 9580
rect 8024 9528 8076 9580
rect 8300 9571 8352 9580
rect 8300 9537 8309 9571
rect 8309 9537 8343 9571
rect 8343 9537 8352 9571
rect 8300 9528 8352 9537
rect 10692 9528 10744 9580
rect 19432 9571 19484 9580
rect 19432 9537 19441 9571
rect 19441 9537 19475 9571
rect 19475 9537 19484 9571
rect 19432 9528 19484 9537
rect 4436 9503 4488 9512
rect 4436 9469 4470 9503
rect 4470 9469 4488 9503
rect 2964 9392 3016 9444
rect 4436 9460 4488 9469
rect 7380 9460 7432 9512
rect 5356 9392 5408 9444
rect 9864 9460 9916 9512
rect 12440 9460 12492 9512
rect 13268 9460 13320 9512
rect 19248 9460 19300 9512
rect 22192 9528 22244 9580
rect 23940 9596 23992 9648
rect 24308 9596 24360 9648
rect 24492 9639 24544 9648
rect 24492 9605 24501 9639
rect 24501 9605 24535 9639
rect 24535 9605 24544 9639
rect 24492 9596 24544 9605
rect 24584 9596 24636 9648
rect 24952 9596 25004 9648
rect 26976 9639 27028 9648
rect 26976 9605 26985 9639
rect 26985 9605 27019 9639
rect 27019 9605 27028 9639
rect 26976 9596 27028 9605
rect 22560 9571 22612 9580
rect 22560 9537 22569 9571
rect 22569 9537 22603 9571
rect 22603 9537 22612 9571
rect 22560 9528 22612 9537
rect 23388 9528 23440 9580
rect 23572 9528 23624 9580
rect 24216 9571 24268 9580
rect 20628 9460 20680 9512
rect 7748 9392 7800 9444
rect 9956 9392 10008 9444
rect 10416 9392 10468 9444
rect 13544 9392 13596 9444
rect 19616 9392 19668 9444
rect 22652 9460 22704 9512
rect 23296 9460 23348 9512
rect 24216 9537 24225 9571
rect 24225 9537 24259 9571
rect 24259 9537 24268 9571
rect 24216 9528 24268 9537
rect 22560 9392 22612 9444
rect 23848 9392 23900 9444
rect 25688 9460 25740 9512
rect 27528 9392 27580 9444
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 2688 9367 2740 9376
rect 2688 9333 2697 9367
rect 2697 9333 2731 9367
rect 2731 9333 2740 9367
rect 2688 9324 2740 9333
rect 5540 9367 5592 9376
rect 5540 9333 5549 9367
rect 5549 9333 5583 9367
rect 5583 9333 5592 9367
rect 5540 9324 5592 9333
rect 7564 9367 7616 9376
rect 7564 9333 7573 9367
rect 7573 9333 7607 9367
rect 7607 9333 7616 9367
rect 7564 9324 7616 9333
rect 8024 9324 8076 9376
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 9864 9324 9916 9376
rect 10692 9324 10744 9376
rect 14004 9324 14056 9376
rect 14464 9324 14516 9376
rect 15568 9324 15620 9376
rect 18236 9367 18288 9376
rect 18236 9333 18245 9367
rect 18245 9333 18279 9367
rect 18279 9333 18288 9367
rect 18236 9324 18288 9333
rect 18788 9324 18840 9376
rect 19156 9324 19208 9376
rect 20812 9324 20864 9376
rect 21272 9324 21324 9376
rect 21456 9367 21508 9376
rect 21456 9333 21465 9367
rect 21465 9333 21499 9367
rect 21499 9333 21508 9367
rect 21456 9324 21508 9333
rect 22008 9367 22060 9376
rect 22008 9333 22017 9367
rect 22017 9333 22051 9367
rect 22051 9333 22060 9367
rect 22008 9324 22060 9333
rect 24124 9367 24176 9376
rect 24124 9333 24133 9367
rect 24133 9333 24167 9367
rect 24167 9333 24176 9367
rect 24124 9324 24176 9333
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 20982 9222 21034 9274
rect 21046 9222 21098 9274
rect 21110 9222 21162 9274
rect 21174 9222 21226 9274
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 4528 9163 4580 9172
rect 4528 9129 4537 9163
rect 4537 9129 4571 9163
rect 4571 9129 4580 9163
rect 4528 9120 4580 9129
rect 7656 9120 7708 9172
rect 7748 9163 7800 9172
rect 7748 9129 7757 9163
rect 7757 9129 7791 9163
rect 7791 9129 7800 9163
rect 7748 9120 7800 9129
rect 8116 9120 8168 9172
rect 8852 9163 8904 9172
rect 8852 9129 8861 9163
rect 8861 9129 8895 9163
rect 8895 9129 8904 9163
rect 8852 9120 8904 9129
rect 13636 9163 13688 9172
rect 13636 9129 13645 9163
rect 13645 9129 13679 9163
rect 13679 9129 13688 9163
rect 13636 9120 13688 9129
rect 19156 9120 19208 9172
rect 19616 9163 19668 9172
rect 19616 9129 19625 9163
rect 19625 9129 19659 9163
rect 19659 9129 19668 9163
rect 19616 9120 19668 9129
rect 22192 9163 22244 9172
rect 22192 9129 22201 9163
rect 22201 9129 22235 9163
rect 22235 9129 22244 9163
rect 22192 9120 22244 9129
rect 22652 9120 22704 9172
rect 26700 9163 26752 9172
rect 26700 9129 26709 9163
rect 26709 9129 26743 9163
rect 26743 9129 26752 9163
rect 26700 9120 26752 9129
rect 1768 9052 1820 9104
rect 8484 9052 8536 9104
rect 13544 9052 13596 9104
rect 19340 9052 19392 9104
rect 20444 9052 20496 9104
rect 25044 9052 25096 9104
rect 2044 8984 2096 9036
rect 7104 9027 7156 9036
rect 7104 8993 7113 9027
rect 7113 8993 7147 9027
rect 7147 8993 7156 9027
rect 7104 8984 7156 8993
rect 8024 8984 8076 9036
rect 8576 8984 8628 9036
rect 9588 8984 9640 9036
rect 10508 8984 10560 9036
rect 16856 8984 16908 9036
rect 20352 8984 20404 9036
rect 21824 9027 21876 9036
rect 21824 8993 21833 9027
rect 21833 8993 21867 9027
rect 21867 8993 21876 9027
rect 21824 8984 21876 8993
rect 23296 8984 23348 9036
rect 26424 8984 26476 9036
rect 8392 8959 8444 8968
rect 8392 8925 8401 8959
rect 8401 8925 8435 8959
rect 8435 8925 8444 8959
rect 8392 8916 8444 8925
rect 16764 8959 16816 8968
rect 16764 8925 16773 8959
rect 16773 8925 16807 8959
rect 16807 8925 16816 8959
rect 16764 8916 16816 8925
rect 23664 8959 23716 8968
rect 23664 8925 23673 8959
rect 23673 8925 23707 8959
rect 23707 8925 23716 8959
rect 23664 8916 23716 8925
rect 24216 8916 24268 8968
rect 2412 8848 2464 8900
rect 2596 8848 2648 8900
rect 9680 8848 9732 8900
rect 1400 8780 1452 8832
rect 5356 8780 5408 8832
rect 10416 8823 10468 8832
rect 10416 8789 10425 8823
rect 10425 8789 10459 8823
rect 10459 8789 10468 8823
rect 10416 8780 10468 8789
rect 14648 8823 14700 8832
rect 14648 8789 14657 8823
rect 14657 8789 14691 8823
rect 14691 8789 14700 8823
rect 14648 8780 14700 8789
rect 18144 8823 18196 8832
rect 18144 8789 18153 8823
rect 18153 8789 18187 8823
rect 18187 8789 18196 8823
rect 18144 8780 18196 8789
rect 19248 8823 19300 8832
rect 19248 8789 19257 8823
rect 19257 8789 19291 8823
rect 19291 8789 19300 8823
rect 19248 8780 19300 8789
rect 20168 8780 20220 8832
rect 21272 8780 21324 8832
rect 21916 8780 21968 8832
rect 22284 8780 22336 8832
rect 23204 8823 23256 8832
rect 23204 8789 23213 8823
rect 23213 8789 23247 8823
rect 23247 8789 23256 8823
rect 23204 8780 23256 8789
rect 24216 8823 24268 8832
rect 24216 8789 24225 8823
rect 24225 8789 24259 8823
rect 24259 8789 24268 8823
rect 24216 8780 24268 8789
rect 25688 8823 25740 8832
rect 25688 8789 25697 8823
rect 25697 8789 25731 8823
rect 25731 8789 25740 8823
rect 25688 8780 25740 8789
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 15982 8678 16034 8730
rect 16046 8678 16098 8730
rect 16110 8678 16162 8730
rect 16174 8678 16226 8730
rect 25982 8678 26034 8730
rect 26046 8678 26098 8730
rect 26110 8678 26162 8730
rect 26174 8678 26226 8730
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 4252 8619 4304 8628
rect 4252 8585 4261 8619
rect 4261 8585 4295 8619
rect 4295 8585 4304 8619
rect 4252 8576 4304 8585
rect 7104 8619 7156 8628
rect 7104 8585 7113 8619
rect 7113 8585 7147 8619
rect 7147 8585 7156 8619
rect 7104 8576 7156 8585
rect 8116 8576 8168 8628
rect 8392 8576 8444 8628
rect 10692 8576 10744 8628
rect 14464 8619 14516 8628
rect 14464 8585 14473 8619
rect 14473 8585 14507 8619
rect 14507 8585 14516 8619
rect 14464 8576 14516 8585
rect 16856 8619 16908 8628
rect 16856 8585 16865 8619
rect 16865 8585 16899 8619
rect 16899 8585 16908 8619
rect 16856 8576 16908 8585
rect 1584 8551 1636 8560
rect 1584 8517 1593 8551
rect 1593 8517 1627 8551
rect 1627 8517 1636 8551
rect 1584 8508 1636 8517
rect 2412 8483 2464 8492
rect 2412 8449 2421 8483
rect 2421 8449 2455 8483
rect 2455 8449 2464 8483
rect 2412 8440 2464 8449
rect 5540 8440 5592 8492
rect 16764 8508 16816 8560
rect 19248 8508 19300 8560
rect 4252 8372 4304 8424
rect 4528 8304 4580 8356
rect 10416 8372 10468 8424
rect 14648 8415 14700 8424
rect 14648 8381 14657 8415
rect 14657 8381 14691 8415
rect 14691 8381 14700 8415
rect 14648 8372 14700 8381
rect 20352 8576 20404 8628
rect 21456 8619 21508 8628
rect 21456 8585 21465 8619
rect 21465 8585 21499 8619
rect 21499 8585 21508 8619
rect 21456 8576 21508 8585
rect 21824 8576 21876 8628
rect 21916 8508 21968 8560
rect 23296 8508 23348 8560
rect 23388 8508 23440 8560
rect 24216 8483 24268 8492
rect 24216 8449 24225 8483
rect 24225 8449 24259 8483
rect 24259 8449 24268 8483
rect 24216 8440 24268 8449
rect 20168 8372 20220 8424
rect 10140 8304 10192 8356
rect 20812 8304 20864 8356
rect 24492 8304 24544 8356
rect 26424 8304 26476 8356
rect 4436 8279 4488 8288
rect 4436 8245 4445 8279
rect 4445 8245 4479 8279
rect 4479 8245 4488 8279
rect 4436 8236 4488 8245
rect 8024 8236 8076 8288
rect 9312 8279 9364 8288
rect 9312 8245 9321 8279
rect 9321 8245 9355 8279
rect 9355 8245 9364 8279
rect 9312 8236 9364 8245
rect 24400 8236 24452 8288
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 20982 8134 21034 8186
rect 21046 8134 21098 8186
rect 21110 8134 21162 8186
rect 21174 8134 21226 8186
rect 1492 8032 1544 8084
rect 4436 8032 4488 8084
rect 10508 8075 10560 8084
rect 10508 8041 10517 8075
rect 10517 8041 10551 8075
rect 10551 8041 10560 8075
rect 10508 8032 10560 8041
rect 21548 8075 21600 8084
rect 21548 8041 21557 8075
rect 21557 8041 21591 8075
rect 21591 8041 21600 8075
rect 21548 8032 21600 8041
rect 22008 8032 22060 8084
rect 23664 8032 23716 8084
rect 24124 8032 24176 8084
rect 24768 8032 24820 8084
rect 26700 8075 26752 8084
rect 26700 8041 26709 8075
rect 26709 8041 26743 8075
rect 26743 8041 26752 8075
rect 26700 8032 26752 8041
rect 5540 7964 5592 8016
rect 5724 7964 5776 8016
rect 24216 7964 24268 8016
rect 1952 7896 2004 7948
rect 4344 7896 4396 7948
rect 11520 7896 11572 7948
rect 15568 7896 15620 7948
rect 21640 7939 21692 7948
rect 21640 7905 21649 7939
rect 21649 7905 21683 7939
rect 21683 7905 21692 7939
rect 21640 7896 21692 7905
rect 25872 7896 25924 7948
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 5356 7828 5408 7880
rect 11428 7871 11480 7880
rect 11428 7837 11437 7871
rect 11437 7837 11471 7871
rect 11471 7837 11480 7871
rect 11428 7828 11480 7837
rect 16396 7871 16448 7880
rect 16396 7837 16405 7871
rect 16405 7837 16439 7871
rect 16439 7837 16448 7871
rect 16396 7828 16448 7837
rect 16580 7871 16632 7880
rect 16580 7837 16589 7871
rect 16589 7837 16623 7871
rect 16623 7837 16632 7871
rect 16580 7828 16632 7837
rect 21732 7871 21784 7880
rect 21732 7837 21741 7871
rect 21741 7837 21775 7871
rect 21775 7837 21784 7871
rect 21732 7828 21784 7837
rect 23940 7828 23992 7880
rect 1768 7692 1820 7744
rect 4068 7735 4120 7744
rect 4068 7701 4077 7735
rect 4077 7701 4111 7735
rect 4111 7701 4120 7735
rect 4068 7692 4120 7701
rect 6368 7692 6420 7744
rect 7380 7692 7432 7744
rect 12808 7735 12860 7744
rect 12808 7701 12817 7735
rect 12817 7701 12851 7735
rect 12851 7701 12860 7735
rect 12808 7692 12860 7701
rect 14648 7692 14700 7744
rect 16304 7692 16356 7744
rect 20168 7735 20220 7744
rect 20168 7701 20177 7735
rect 20177 7701 20211 7735
rect 20211 7701 20220 7735
rect 20168 7692 20220 7701
rect 20720 7692 20772 7744
rect 25044 7735 25096 7744
rect 25044 7701 25053 7735
rect 25053 7701 25087 7735
rect 25087 7701 25096 7735
rect 25044 7692 25096 7701
rect 25688 7692 25740 7744
rect 26792 7692 26844 7744
rect 27068 7692 27120 7744
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 15982 7590 16034 7642
rect 16046 7590 16098 7642
rect 16110 7590 16162 7642
rect 16174 7590 16226 7642
rect 25982 7590 26034 7642
rect 26046 7590 26098 7642
rect 26110 7590 26162 7642
rect 26174 7590 26226 7642
rect 4344 7488 4396 7540
rect 4436 7488 4488 7540
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 10140 7531 10192 7540
rect 10140 7497 10149 7531
rect 10149 7497 10183 7531
rect 10183 7497 10192 7531
rect 10140 7488 10192 7497
rect 11520 7531 11572 7540
rect 11520 7497 11529 7531
rect 11529 7497 11563 7531
rect 11563 7497 11572 7531
rect 11520 7488 11572 7497
rect 5540 7420 5592 7472
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 2688 7284 2740 7336
rect 5356 7327 5408 7336
rect 5356 7293 5365 7327
rect 5365 7293 5399 7327
rect 5399 7293 5408 7327
rect 5356 7284 5408 7293
rect 6644 7327 6696 7336
rect 6644 7293 6653 7327
rect 6653 7293 6687 7327
rect 6687 7293 6696 7327
rect 7288 7327 7340 7336
rect 6644 7284 6696 7293
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 8760 7327 8812 7336
rect 8760 7293 8769 7327
rect 8769 7293 8803 7327
rect 8803 7293 8812 7327
rect 8760 7284 8812 7293
rect 9312 7284 9364 7336
rect 11428 7284 11480 7336
rect 12440 7488 12492 7540
rect 20812 7488 20864 7540
rect 21732 7488 21784 7540
rect 24400 7531 24452 7540
rect 24400 7497 24409 7531
rect 24409 7497 24443 7531
rect 24443 7497 24452 7531
rect 24400 7488 24452 7497
rect 25596 7488 25648 7540
rect 27528 7531 27580 7540
rect 27528 7497 27537 7531
rect 27537 7497 27571 7531
rect 27571 7497 27580 7531
rect 27528 7488 27580 7497
rect 13084 7420 13136 7472
rect 16396 7420 16448 7472
rect 24216 7463 24268 7472
rect 24216 7429 24225 7463
rect 24225 7429 24259 7463
rect 24259 7429 24268 7463
rect 24216 7420 24268 7429
rect 13268 7352 13320 7404
rect 14648 7352 14700 7404
rect 16856 7352 16908 7404
rect 1768 7259 1820 7268
rect 1768 7225 1802 7259
rect 1802 7225 1820 7259
rect 1768 7216 1820 7225
rect 4620 7216 4672 7268
rect 6368 7216 6420 7268
rect 9588 7216 9640 7268
rect 13452 7216 13504 7268
rect 2872 7191 2924 7200
rect 2872 7157 2881 7191
rect 2881 7157 2915 7191
rect 2915 7157 2924 7191
rect 2872 7148 2924 7157
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 12164 7191 12216 7200
rect 12164 7157 12173 7191
rect 12173 7157 12207 7191
rect 12207 7157 12216 7191
rect 12164 7148 12216 7157
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 13360 7191 13412 7200
rect 13360 7157 13369 7191
rect 13369 7157 13403 7191
rect 13403 7157 13412 7191
rect 15752 7284 15804 7336
rect 16580 7284 16632 7336
rect 18144 7284 18196 7336
rect 19340 7284 19392 7336
rect 19892 7327 19944 7336
rect 19892 7293 19901 7327
rect 19901 7293 19935 7327
rect 19935 7293 19944 7327
rect 19892 7284 19944 7293
rect 25044 7395 25096 7404
rect 25044 7361 25053 7395
rect 25053 7361 25087 7395
rect 25087 7361 25096 7395
rect 25044 7352 25096 7361
rect 25688 7352 25740 7404
rect 20628 7284 20680 7336
rect 24216 7284 24268 7336
rect 25964 7327 26016 7336
rect 25964 7293 25973 7327
rect 25973 7293 26007 7327
rect 26007 7293 26016 7327
rect 25964 7284 26016 7293
rect 14372 7259 14424 7268
rect 14372 7225 14381 7259
rect 14381 7225 14415 7259
rect 14415 7225 14424 7259
rect 14372 7216 14424 7225
rect 15384 7216 15436 7268
rect 13360 7148 13412 7157
rect 14556 7148 14608 7200
rect 14924 7191 14976 7200
rect 14924 7157 14933 7191
rect 14933 7157 14967 7191
rect 14967 7157 14976 7191
rect 15568 7191 15620 7200
rect 14924 7148 14976 7157
rect 15568 7157 15577 7191
rect 15577 7157 15611 7191
rect 15611 7157 15620 7191
rect 15568 7148 15620 7157
rect 16120 7148 16172 7200
rect 16672 7216 16724 7268
rect 25596 7216 25648 7268
rect 26792 7216 26844 7268
rect 18972 7148 19024 7200
rect 23940 7191 23992 7200
rect 23940 7157 23949 7191
rect 23949 7157 23983 7191
rect 23983 7157 23992 7191
rect 23940 7148 23992 7157
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 20982 7046 21034 7098
rect 21046 7046 21098 7098
rect 21110 7046 21162 7098
rect 21174 7046 21226 7098
rect 1952 6987 2004 6996
rect 1952 6953 1961 6987
rect 1961 6953 1995 6987
rect 1995 6953 2004 6987
rect 1952 6944 2004 6953
rect 3700 6944 3752 6996
rect 4068 6944 4120 6996
rect 6184 6987 6236 6996
rect 6184 6953 6193 6987
rect 6193 6953 6227 6987
rect 6227 6953 6236 6987
rect 6184 6944 6236 6953
rect 12900 6944 12952 6996
rect 13268 6987 13320 6996
rect 13268 6953 13277 6987
rect 13277 6953 13311 6987
rect 13311 6953 13320 6987
rect 13268 6944 13320 6953
rect 14556 6987 14608 6996
rect 14556 6953 14565 6987
rect 14565 6953 14599 6987
rect 14599 6953 14608 6987
rect 14556 6944 14608 6953
rect 18972 6987 19024 6996
rect 18972 6953 18981 6987
rect 18981 6953 19015 6987
rect 19015 6953 19024 6987
rect 18972 6944 19024 6953
rect 19340 6944 19392 6996
rect 19892 6987 19944 6996
rect 19892 6953 19901 6987
rect 19901 6953 19935 6987
rect 19935 6953 19944 6987
rect 19892 6944 19944 6953
rect 21640 6944 21692 6996
rect 23204 6944 23256 6996
rect 24124 6987 24176 6996
rect 24124 6953 24133 6987
rect 24133 6953 24167 6987
rect 24167 6953 24176 6987
rect 24124 6944 24176 6953
rect 24768 6987 24820 6996
rect 24768 6953 24777 6987
rect 24777 6953 24811 6987
rect 24811 6953 24820 6987
rect 24768 6944 24820 6953
rect 24952 6944 25004 6996
rect 3884 6876 3936 6928
rect 11520 6876 11572 6928
rect 21548 6919 21600 6928
rect 21548 6885 21557 6919
rect 21557 6885 21591 6919
rect 21591 6885 21600 6919
rect 21548 6876 21600 6885
rect 23296 6876 23348 6928
rect 2136 6808 2188 6860
rect 4344 6808 4396 6860
rect 4712 6808 4764 6860
rect 7196 6808 7248 6860
rect 11060 6808 11112 6860
rect 13084 6808 13136 6860
rect 16856 6808 16908 6860
rect 19064 6851 19116 6860
rect 4620 6783 4672 6792
rect 4620 6749 4629 6783
rect 4629 6749 4663 6783
rect 4663 6749 4672 6783
rect 4620 6740 4672 6749
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 10140 6783 10192 6792
rect 6368 6740 6420 6749
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 12808 6783 12860 6792
rect 10232 6740 10284 6749
rect 12808 6749 12817 6783
rect 12817 6749 12851 6783
rect 12851 6749 12860 6783
rect 12808 6740 12860 6749
rect 16120 6783 16172 6792
rect 16120 6749 16129 6783
rect 16129 6749 16163 6783
rect 16163 6749 16172 6783
rect 16120 6740 16172 6749
rect 17500 6783 17552 6792
rect 17500 6749 17509 6783
rect 17509 6749 17543 6783
rect 17543 6749 17552 6783
rect 17500 6740 17552 6749
rect 17592 6783 17644 6792
rect 17592 6749 17601 6783
rect 17601 6749 17635 6783
rect 17635 6749 17644 6783
rect 18144 6783 18196 6792
rect 17592 6740 17644 6749
rect 18144 6749 18153 6783
rect 18153 6749 18187 6783
rect 18187 6749 18196 6783
rect 18144 6740 18196 6749
rect 1584 6715 1636 6724
rect 1584 6681 1593 6715
rect 1593 6681 1627 6715
rect 1627 6681 1636 6715
rect 1584 6672 1636 6681
rect 19064 6817 19073 6851
rect 19073 6817 19107 6851
rect 19107 6817 19116 6851
rect 19064 6808 19116 6817
rect 22928 6851 22980 6860
rect 22928 6817 22937 6851
rect 22937 6817 22971 6851
rect 22971 6817 22980 6851
rect 22928 6808 22980 6817
rect 23388 6808 23440 6860
rect 23756 6808 23808 6860
rect 24400 6808 24452 6860
rect 26976 6808 27028 6860
rect 18696 6672 18748 6724
rect 22560 6740 22612 6792
rect 25044 6783 25096 6792
rect 25044 6749 25053 6783
rect 25053 6749 25087 6783
rect 25087 6749 25096 6783
rect 25044 6740 25096 6749
rect 21640 6672 21692 6724
rect 24492 6672 24544 6724
rect 26700 6715 26752 6724
rect 26700 6681 26709 6715
rect 26709 6681 26743 6715
rect 26743 6681 26752 6715
rect 26700 6672 26752 6681
rect 2688 6604 2740 6656
rect 3608 6604 3660 6656
rect 5448 6604 5500 6656
rect 7288 6647 7340 6656
rect 7288 6613 7297 6647
rect 7297 6613 7331 6647
rect 7331 6613 7340 6647
rect 7288 6604 7340 6613
rect 8760 6647 8812 6656
rect 8760 6613 8769 6647
rect 8769 6613 8803 6647
rect 8803 6613 8812 6647
rect 8760 6604 8812 6613
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 9680 6604 9732 6613
rect 11060 6604 11112 6656
rect 16396 6604 16448 6656
rect 21088 6604 21140 6656
rect 26792 6604 26844 6656
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 15982 6502 16034 6554
rect 16046 6502 16098 6554
rect 16110 6502 16162 6554
rect 16174 6502 16226 6554
rect 25982 6502 26034 6554
rect 26046 6502 26098 6554
rect 26110 6502 26162 6554
rect 26174 6502 26226 6554
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 2136 6400 2188 6452
rect 5816 6400 5868 6452
rect 10140 6400 10192 6452
rect 11060 6443 11112 6452
rect 11060 6409 11069 6443
rect 11069 6409 11103 6443
rect 11103 6409 11112 6443
rect 11060 6400 11112 6409
rect 12900 6400 12952 6452
rect 13084 6443 13136 6452
rect 13084 6409 13093 6443
rect 13093 6409 13127 6443
rect 13127 6409 13136 6443
rect 13084 6400 13136 6409
rect 17500 6443 17552 6452
rect 17500 6409 17509 6443
rect 17509 6409 17543 6443
rect 17543 6409 17552 6443
rect 17500 6400 17552 6409
rect 19064 6443 19116 6452
rect 19064 6409 19073 6443
rect 19073 6409 19107 6443
rect 19107 6409 19116 6443
rect 19064 6400 19116 6409
rect 19340 6400 19392 6452
rect 20444 6443 20496 6452
rect 20444 6409 20453 6443
rect 20453 6409 20487 6443
rect 20487 6409 20496 6443
rect 20444 6400 20496 6409
rect 22560 6443 22612 6452
rect 22560 6409 22569 6443
rect 22569 6409 22603 6443
rect 22603 6409 22612 6443
rect 22560 6400 22612 6409
rect 22928 6443 22980 6452
rect 22928 6409 22937 6443
rect 22937 6409 22971 6443
rect 22971 6409 22980 6443
rect 22928 6400 22980 6409
rect 23204 6443 23256 6452
rect 23204 6409 23213 6443
rect 23213 6409 23247 6443
rect 23247 6409 23256 6443
rect 23204 6400 23256 6409
rect 24400 6443 24452 6452
rect 24400 6409 24409 6443
rect 24409 6409 24443 6443
rect 24443 6409 24452 6443
rect 24400 6400 24452 6409
rect 24676 6400 24728 6452
rect 25044 6400 25096 6452
rect 26792 6400 26844 6452
rect 26976 6443 27028 6452
rect 26976 6409 26985 6443
rect 26985 6409 27019 6443
rect 27019 6409 27028 6443
rect 26976 6400 27028 6409
rect 4068 6332 4120 6384
rect 10232 6332 10284 6384
rect 3700 6307 3752 6316
rect 3700 6273 3709 6307
rect 3709 6273 3743 6307
rect 3743 6273 3752 6307
rect 3700 6264 3752 6273
rect 5448 6307 5500 6316
rect 2044 6196 2096 6248
rect 3608 6239 3660 6248
rect 3608 6205 3617 6239
rect 3617 6205 3651 6239
rect 3651 6205 3660 6239
rect 3608 6196 3660 6205
rect 5448 6273 5457 6307
rect 5457 6273 5491 6307
rect 5491 6273 5500 6307
rect 5448 6264 5500 6273
rect 7656 6307 7708 6316
rect 2872 6128 2924 6180
rect 5080 6196 5132 6248
rect 7288 6196 7340 6248
rect 7656 6273 7665 6307
rect 7665 6273 7699 6307
rect 7699 6273 7708 6307
rect 7656 6264 7708 6273
rect 9588 6264 9640 6316
rect 12808 6264 12860 6316
rect 16304 6307 16356 6316
rect 16304 6273 16313 6307
rect 16313 6273 16347 6307
rect 16347 6273 16356 6307
rect 16304 6264 16356 6273
rect 17224 6332 17276 6384
rect 17592 6332 17644 6384
rect 18144 6264 18196 6316
rect 18604 6307 18656 6316
rect 18604 6273 18613 6307
rect 18613 6273 18647 6307
rect 18647 6273 18656 6307
rect 18604 6264 18656 6273
rect 21088 6307 21140 6316
rect 21088 6273 21097 6307
rect 21097 6273 21131 6307
rect 21131 6273 21140 6307
rect 21088 6264 21140 6273
rect 26240 6307 26292 6316
rect 26240 6273 26249 6307
rect 26249 6273 26283 6307
rect 26283 6273 26292 6307
rect 26240 6264 26292 6273
rect 7840 6196 7892 6248
rect 18420 6239 18472 6248
rect 18420 6205 18429 6239
rect 18429 6205 18463 6239
rect 18463 6205 18472 6239
rect 18420 6196 18472 6205
rect 20444 6196 20496 6248
rect 5448 6128 5500 6180
rect 10784 6128 10836 6180
rect 15752 6128 15804 6180
rect 1400 6060 1452 6112
rect 3240 6103 3292 6112
rect 3240 6069 3249 6103
rect 3249 6069 3283 6103
rect 3283 6069 3292 6103
rect 3240 6060 3292 6069
rect 4344 6103 4396 6112
rect 4344 6069 4353 6103
rect 4353 6069 4387 6103
rect 4387 6069 4396 6103
rect 4344 6060 4396 6069
rect 4712 6103 4764 6112
rect 4712 6069 4721 6103
rect 4721 6069 4755 6103
rect 4755 6069 4764 6103
rect 4712 6060 4764 6069
rect 7380 6060 7432 6112
rect 7656 6060 7708 6112
rect 10324 6103 10376 6112
rect 10324 6069 10333 6103
rect 10333 6069 10367 6103
rect 10367 6069 10376 6103
rect 10324 6060 10376 6069
rect 15844 6103 15896 6112
rect 15844 6069 15853 6103
rect 15853 6069 15887 6103
rect 15887 6069 15896 6103
rect 15844 6060 15896 6069
rect 17960 6060 18012 6112
rect 18512 6103 18564 6112
rect 18512 6069 18521 6103
rect 18521 6069 18555 6103
rect 18555 6069 18564 6103
rect 18512 6060 18564 6069
rect 20536 6103 20588 6112
rect 20536 6069 20545 6103
rect 20545 6069 20579 6103
rect 20579 6069 20588 6103
rect 20536 6060 20588 6069
rect 20812 6060 20864 6112
rect 24768 6103 24820 6112
rect 24768 6069 24777 6103
rect 24777 6069 24811 6103
rect 24811 6069 24820 6103
rect 24768 6060 24820 6069
rect 26608 6103 26660 6112
rect 26608 6069 26617 6103
rect 26617 6069 26651 6103
rect 26651 6069 26660 6103
rect 26608 6060 26660 6069
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 20982 5958 21034 6010
rect 21046 5958 21098 6010
rect 21110 5958 21162 6010
rect 21174 5958 21226 6010
rect 4620 5856 4672 5908
rect 5080 5899 5132 5908
rect 5080 5865 5089 5899
rect 5089 5865 5123 5899
rect 5123 5865 5132 5899
rect 5080 5856 5132 5865
rect 5448 5899 5500 5908
rect 5448 5865 5457 5899
rect 5457 5865 5491 5899
rect 5491 5865 5500 5899
rect 5448 5856 5500 5865
rect 6276 5856 6328 5908
rect 9588 5856 9640 5908
rect 10324 5899 10376 5908
rect 10324 5865 10333 5899
rect 10333 5865 10367 5899
rect 10367 5865 10376 5899
rect 10324 5856 10376 5865
rect 10692 5856 10744 5908
rect 12348 5856 12400 5908
rect 12716 5856 12768 5908
rect 17224 5899 17276 5908
rect 17224 5865 17233 5899
rect 17233 5865 17267 5899
rect 17267 5865 17276 5899
rect 17224 5856 17276 5865
rect 17960 5856 18012 5908
rect 18604 5899 18656 5908
rect 18604 5865 18613 5899
rect 18613 5865 18647 5899
rect 18647 5865 18656 5899
rect 18604 5856 18656 5865
rect 19248 5856 19300 5908
rect 20536 5856 20588 5908
rect 20812 5856 20864 5908
rect 2780 5788 2832 5840
rect 7748 5788 7800 5840
rect 12532 5831 12584 5840
rect 12532 5797 12541 5831
rect 12541 5797 12575 5831
rect 12575 5797 12584 5831
rect 12532 5788 12584 5797
rect 16304 5788 16356 5840
rect 16488 5788 16540 5840
rect 2688 5720 2740 5772
rect 7472 5763 7524 5772
rect 7472 5729 7481 5763
rect 7481 5729 7515 5763
rect 7515 5729 7524 5763
rect 10968 5763 11020 5772
rect 7472 5720 7524 5729
rect 10968 5729 10977 5763
rect 10977 5729 11011 5763
rect 11011 5729 11020 5763
rect 10968 5720 11020 5729
rect 12440 5720 12492 5772
rect 13268 5720 13320 5772
rect 15660 5720 15712 5772
rect 22468 5720 22520 5772
rect 26516 5763 26568 5772
rect 26516 5729 26525 5763
rect 26525 5729 26559 5763
rect 26559 5729 26568 5763
rect 26516 5720 26568 5729
rect 6920 5652 6972 5704
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 11520 5652 11572 5704
rect 19708 5695 19760 5704
rect 2872 5559 2924 5568
rect 2872 5525 2881 5559
rect 2881 5525 2915 5559
rect 2915 5525 2924 5559
rect 2872 5516 2924 5525
rect 7012 5559 7064 5568
rect 7012 5525 7021 5559
rect 7021 5525 7055 5559
rect 7055 5525 7064 5559
rect 7012 5516 7064 5525
rect 19708 5661 19717 5695
rect 19717 5661 19751 5695
rect 19751 5661 19760 5695
rect 19708 5652 19760 5661
rect 19432 5584 19484 5636
rect 22376 5695 22428 5704
rect 22376 5661 22385 5695
rect 22385 5661 22419 5695
rect 22419 5661 22428 5695
rect 22376 5652 22428 5661
rect 23848 5652 23900 5704
rect 27436 5652 27488 5704
rect 13636 5516 13688 5568
rect 19340 5516 19392 5568
rect 23848 5516 23900 5568
rect 25504 5559 25556 5568
rect 25504 5525 25513 5559
rect 25513 5525 25547 5559
rect 25547 5525 25556 5559
rect 25504 5516 25556 5525
rect 26700 5559 26752 5568
rect 26700 5525 26709 5559
rect 26709 5525 26743 5559
rect 26743 5525 26752 5559
rect 26700 5516 26752 5525
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 15982 5414 16034 5466
rect 16046 5414 16098 5466
rect 16110 5414 16162 5466
rect 16174 5414 16226 5466
rect 25982 5414 26034 5466
rect 26046 5414 26098 5466
rect 26110 5414 26162 5466
rect 26174 5414 26226 5466
rect 1584 5355 1636 5364
rect 1584 5321 1593 5355
rect 1593 5321 1627 5355
rect 1627 5321 1636 5355
rect 1584 5312 1636 5321
rect 2872 5312 2924 5364
rect 4068 5312 4120 5364
rect 6644 5355 6696 5364
rect 6644 5321 6653 5355
rect 6653 5321 6687 5355
rect 6687 5321 6696 5355
rect 6644 5312 6696 5321
rect 6920 5312 6972 5364
rect 7748 5312 7800 5364
rect 10784 5355 10836 5364
rect 10784 5321 10793 5355
rect 10793 5321 10827 5355
rect 10827 5321 10836 5355
rect 10784 5312 10836 5321
rect 12348 5312 12400 5364
rect 12532 5312 12584 5364
rect 14648 5355 14700 5364
rect 14648 5321 14657 5355
rect 14657 5321 14691 5355
rect 14691 5321 14700 5355
rect 14648 5312 14700 5321
rect 15752 5312 15804 5364
rect 16304 5312 16356 5364
rect 2780 5176 2832 5228
rect 3240 5176 3292 5228
rect 10968 5244 11020 5296
rect 7288 5176 7340 5228
rect 11520 5176 11572 5228
rect 13268 5219 13320 5228
rect 13268 5185 13277 5219
rect 13277 5185 13311 5219
rect 13311 5185 13320 5219
rect 13268 5176 13320 5185
rect 19248 5312 19300 5364
rect 19708 5355 19760 5364
rect 19708 5321 19717 5355
rect 19717 5321 19751 5355
rect 19751 5321 19760 5355
rect 19708 5312 19760 5321
rect 26516 5312 26568 5364
rect 22468 5287 22520 5296
rect 20352 5219 20404 5228
rect 20352 5185 20361 5219
rect 20361 5185 20395 5219
rect 20395 5185 20404 5219
rect 22468 5253 22477 5287
rect 22477 5253 22511 5287
rect 22511 5253 22520 5287
rect 22468 5244 22520 5253
rect 26792 5287 26844 5296
rect 26792 5253 26801 5287
rect 26801 5253 26835 5287
rect 26835 5253 26844 5287
rect 26792 5244 26844 5253
rect 20352 5176 20404 5185
rect 8116 5151 8168 5160
rect 8116 5117 8125 5151
rect 8125 5117 8159 5151
rect 8159 5117 8168 5151
rect 8116 5108 8168 5117
rect 15200 5108 15252 5160
rect 16488 5108 16540 5160
rect 21272 5176 21324 5228
rect 4068 5040 4120 5092
rect 2136 4972 2188 5024
rect 3148 4972 3200 5024
rect 5816 4972 5868 5024
rect 7656 5040 7708 5092
rect 12072 5040 12124 5092
rect 13636 5040 13688 5092
rect 15660 5040 15712 5092
rect 16212 5040 16264 5092
rect 20536 5040 20588 5092
rect 25504 5108 25556 5160
rect 9496 5015 9548 5024
rect 9496 4981 9505 5015
rect 9505 4981 9539 5015
rect 9539 4981 9548 5015
rect 9496 4972 9548 4981
rect 11336 4972 11388 5024
rect 11888 5015 11940 5024
rect 11888 4981 11897 5015
rect 11897 4981 11931 5015
rect 11931 4981 11940 5015
rect 11888 4972 11940 4981
rect 16120 4972 16172 5024
rect 16672 4972 16724 5024
rect 19432 4972 19484 5024
rect 20168 4972 20220 5024
rect 22376 4972 22428 5024
rect 23572 4972 23624 5024
rect 24952 4972 25004 5024
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 20982 4870 21034 4922
rect 21046 4870 21098 4922
rect 21110 4870 21162 4922
rect 21174 4870 21226 4922
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 3240 4768 3292 4820
rect 7012 4768 7064 4820
rect 7472 4768 7524 4820
rect 8116 4811 8168 4820
rect 8116 4777 8125 4811
rect 8125 4777 8159 4811
rect 8159 4777 8168 4811
rect 8116 4768 8168 4777
rect 10692 4768 10744 4820
rect 11336 4768 11388 4820
rect 11796 4811 11848 4820
rect 11796 4777 11805 4811
rect 11805 4777 11839 4811
rect 11839 4777 11848 4811
rect 11796 4768 11848 4777
rect 11888 4768 11940 4820
rect 13452 4768 13504 4820
rect 16120 4811 16172 4820
rect 16120 4777 16129 4811
rect 16129 4777 16163 4811
rect 16163 4777 16172 4811
rect 16120 4768 16172 4777
rect 19340 4768 19392 4820
rect 20536 4811 20588 4820
rect 20536 4777 20545 4811
rect 20545 4777 20579 4811
rect 20579 4777 20588 4811
rect 20536 4768 20588 4777
rect 11520 4700 11572 4752
rect 2044 4675 2096 4684
rect 2044 4641 2053 4675
rect 2053 4641 2087 4675
rect 2087 4641 2096 4675
rect 2044 4632 2096 4641
rect 2596 4632 2648 4684
rect 4896 4675 4948 4684
rect 4896 4641 4930 4675
rect 4930 4641 4948 4675
rect 4896 4632 4948 4641
rect 7380 4632 7432 4684
rect 2688 4564 2740 4616
rect 4620 4607 4672 4616
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 7196 4564 7248 4616
rect 9496 4564 9548 4616
rect 11520 4564 11572 4616
rect 15384 4700 15436 4752
rect 17224 4700 17276 4752
rect 13544 4632 13596 4684
rect 16212 4675 16264 4684
rect 16212 4641 16221 4675
rect 16221 4641 16255 4675
rect 16255 4641 16264 4675
rect 16212 4632 16264 4641
rect 23572 4675 23624 4684
rect 23572 4641 23581 4675
rect 23581 4641 23615 4675
rect 23615 4641 23624 4675
rect 23572 4632 23624 4641
rect 23848 4675 23900 4684
rect 23848 4641 23882 4675
rect 23882 4641 23900 4675
rect 23848 4632 23900 4641
rect 26516 4675 26568 4684
rect 26516 4641 26525 4675
rect 26525 4641 26559 4675
rect 26559 4641 26568 4675
rect 26516 4632 26568 4641
rect 27160 4632 27212 4684
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 13636 4607 13688 4616
rect 13636 4573 13645 4607
rect 13645 4573 13679 4607
rect 13679 4573 13688 4607
rect 13636 4564 13688 4573
rect 19708 4607 19760 4616
rect 19708 4573 19717 4607
rect 19717 4573 19751 4607
rect 19751 4573 19760 4607
rect 19708 4564 19760 4573
rect 19892 4607 19944 4616
rect 19892 4573 19901 4607
rect 19901 4573 19935 4607
rect 19935 4573 19944 4607
rect 19892 4564 19944 4573
rect 24952 4539 25004 4548
rect 24952 4505 24961 4539
rect 24961 4505 24995 4539
rect 24995 4505 25004 4539
rect 24952 4496 25004 4505
rect 2780 4428 2832 4480
rect 5816 4428 5868 4480
rect 7104 4471 7156 4480
rect 7104 4437 7113 4471
rect 7113 4437 7147 4471
rect 7147 4437 7156 4471
rect 7104 4428 7156 4437
rect 17592 4471 17644 4480
rect 17592 4437 17601 4471
rect 17601 4437 17635 4471
rect 17635 4437 17644 4471
rect 17592 4428 17644 4437
rect 19248 4471 19300 4480
rect 19248 4437 19257 4471
rect 19257 4437 19291 4471
rect 19291 4437 19300 4471
rect 19248 4428 19300 4437
rect 21364 4428 21416 4480
rect 21640 4471 21692 4480
rect 21640 4437 21649 4471
rect 21649 4437 21683 4471
rect 21683 4437 21692 4471
rect 21640 4428 21692 4437
rect 26700 4471 26752 4480
rect 26700 4437 26709 4471
rect 26709 4437 26743 4471
rect 26743 4437 26752 4471
rect 26700 4428 26752 4437
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 15982 4326 16034 4378
rect 16046 4326 16098 4378
rect 16110 4326 16162 4378
rect 16174 4326 16226 4378
rect 25982 4326 26034 4378
rect 26046 4326 26098 4378
rect 26110 4326 26162 4378
rect 26174 4326 26226 4378
rect 2596 4267 2648 4276
rect 2596 4233 2605 4267
rect 2605 4233 2639 4267
rect 2639 4233 2648 4267
rect 2596 4224 2648 4233
rect 4344 4224 4396 4276
rect 4896 4224 4948 4276
rect 7196 4267 7248 4276
rect 7196 4233 7205 4267
rect 7205 4233 7239 4267
rect 7239 4233 7248 4267
rect 7196 4224 7248 4233
rect 7472 4267 7524 4276
rect 7472 4233 7481 4267
rect 7481 4233 7515 4267
rect 7515 4233 7524 4267
rect 7472 4224 7524 4233
rect 11520 4267 11572 4276
rect 11520 4233 11529 4267
rect 11529 4233 11563 4267
rect 11563 4233 11572 4267
rect 11520 4224 11572 4233
rect 12072 4224 12124 4276
rect 13452 4267 13504 4276
rect 13452 4233 13461 4267
rect 13461 4233 13495 4267
rect 13495 4233 13504 4267
rect 13452 4224 13504 4233
rect 13636 4224 13688 4276
rect 17224 4224 17276 4276
rect 19892 4224 19944 4276
rect 21272 4224 21324 4276
rect 23572 4224 23624 4276
rect 27160 4267 27212 4276
rect 27160 4233 27169 4267
rect 27169 4233 27203 4267
rect 27203 4233 27212 4267
rect 27160 4224 27212 4233
rect 4620 4156 4672 4208
rect 7012 4088 7064 4140
rect 7380 4156 7432 4208
rect 11796 4199 11848 4208
rect 11796 4165 11805 4199
rect 11805 4165 11839 4199
rect 11839 4165 11848 4199
rect 11796 4156 11848 4165
rect 13544 4156 13596 4208
rect 8116 4088 8168 4140
rect 15936 4088 15988 4140
rect 16488 4131 16540 4140
rect 16488 4097 16497 4131
rect 16497 4097 16531 4131
rect 16531 4097 16540 4131
rect 16488 4088 16540 4097
rect 19708 4088 19760 4140
rect 21456 4156 21508 4208
rect 20628 4131 20680 4140
rect 20628 4097 20637 4131
rect 20637 4097 20671 4131
rect 20671 4097 20680 4131
rect 20628 4088 20680 4097
rect 21364 4131 21416 4140
rect 21364 4097 21373 4131
rect 21373 4097 21407 4131
rect 21407 4097 21416 4131
rect 21364 4088 21416 4097
rect 21640 4088 21692 4140
rect 2688 4020 2740 4072
rect 2872 4020 2924 4072
rect 5264 4063 5316 4072
rect 5264 4029 5273 4063
rect 5273 4029 5307 4063
rect 5307 4029 5316 4063
rect 5264 4020 5316 4029
rect 19432 4020 19484 4072
rect 23848 4063 23900 4072
rect 2044 3995 2096 4004
rect 2044 3961 2053 3995
rect 2053 3961 2087 3995
rect 2087 3961 2096 3995
rect 2044 3952 2096 3961
rect 3976 3952 4028 4004
rect 1492 3884 1544 3936
rect 16304 3995 16356 4004
rect 16304 3961 16313 3995
rect 16313 3961 16347 3995
rect 16347 3961 16356 3995
rect 16304 3952 16356 3961
rect 20352 3995 20404 4004
rect 20352 3961 20361 3995
rect 20361 3961 20395 3995
rect 20395 3961 20404 3995
rect 23848 4029 23857 4063
rect 23857 4029 23891 4063
rect 23891 4029 23900 4063
rect 23848 4020 23900 4029
rect 26332 4020 26384 4072
rect 26608 4020 26660 4072
rect 20352 3952 20404 3961
rect 15844 3884 15896 3936
rect 20444 3927 20496 3936
rect 20444 3893 20453 3927
rect 20453 3893 20487 3927
rect 20487 3893 20496 3927
rect 22008 3952 22060 4004
rect 20444 3884 20496 3893
rect 26700 3884 26752 3936
rect 27528 3927 27580 3936
rect 27528 3893 27537 3927
rect 27537 3893 27571 3927
rect 27571 3893 27580 3927
rect 27528 3884 27580 3893
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 20982 3782 21034 3834
rect 21046 3782 21098 3834
rect 21110 3782 21162 3834
rect 21174 3782 21226 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 2872 3680 2924 3732
rect 4344 3723 4396 3732
rect 4344 3689 4353 3723
rect 4353 3689 4387 3723
rect 4387 3689 4396 3723
rect 4344 3680 4396 3689
rect 5172 3680 5224 3732
rect 5632 3680 5684 3732
rect 6828 3680 6880 3732
rect 7564 3680 7616 3732
rect 12072 3680 12124 3732
rect 15936 3723 15988 3732
rect 15936 3689 15945 3723
rect 15945 3689 15979 3723
rect 15979 3689 15988 3723
rect 15936 3680 15988 3689
rect 19340 3723 19392 3732
rect 19340 3689 19349 3723
rect 19349 3689 19383 3723
rect 19383 3689 19392 3723
rect 19340 3680 19392 3689
rect 20444 3680 20496 3732
rect 2688 3612 2740 3664
rect 4620 3612 4672 3664
rect 4988 3612 5040 3664
rect 15660 3612 15712 3664
rect 2596 3544 2648 3596
rect 6276 3544 6328 3596
rect 5816 3476 5868 3528
rect 6552 3476 6604 3528
rect 8024 3544 8076 3596
rect 11060 3587 11112 3596
rect 11060 3553 11094 3587
rect 11094 3553 11112 3587
rect 11060 3544 11112 3553
rect 16488 3612 16540 3664
rect 17592 3612 17644 3664
rect 20352 3655 20404 3664
rect 20352 3621 20361 3655
rect 20361 3621 20395 3655
rect 20395 3621 20404 3655
rect 20352 3612 20404 3621
rect 20812 3612 20864 3664
rect 21824 3680 21876 3732
rect 17776 3544 17828 3596
rect 25320 3587 25372 3596
rect 25320 3553 25329 3587
rect 25329 3553 25363 3587
rect 25363 3553 25372 3587
rect 25320 3544 25372 3553
rect 27344 3544 27396 3596
rect 8760 3476 8812 3528
rect 10784 3519 10836 3528
rect 10784 3485 10793 3519
rect 10793 3485 10827 3519
rect 10827 3485 10836 3519
rect 10784 3476 10836 3485
rect 20720 3476 20772 3528
rect 21364 3519 21416 3528
rect 21364 3485 21373 3519
rect 21373 3485 21407 3519
rect 21407 3485 21416 3519
rect 21364 3476 21416 3485
rect 21456 3519 21508 3528
rect 21456 3485 21465 3519
rect 21465 3485 21499 3519
rect 21499 3485 21508 3519
rect 21456 3476 21508 3485
rect 25504 3451 25556 3460
rect 25504 3417 25513 3451
rect 25513 3417 25547 3451
rect 25547 3417 25556 3451
rect 25504 3408 25556 3417
rect 2688 3383 2740 3392
rect 2688 3349 2697 3383
rect 2697 3349 2731 3383
rect 2731 3349 2740 3383
rect 2688 3340 2740 3349
rect 4896 3383 4948 3392
rect 4896 3349 4905 3383
rect 4905 3349 4939 3383
rect 4939 3349 4948 3383
rect 4896 3340 4948 3349
rect 5448 3340 5500 3392
rect 6920 3383 6972 3392
rect 6920 3349 6929 3383
rect 6929 3349 6963 3383
rect 6963 3349 6972 3383
rect 6920 3340 6972 3349
rect 7288 3340 7340 3392
rect 18604 3383 18656 3392
rect 18604 3349 18613 3383
rect 18613 3349 18647 3383
rect 18647 3349 18656 3383
rect 18604 3340 18656 3349
rect 26700 3383 26752 3392
rect 26700 3349 26709 3383
rect 26709 3349 26743 3383
rect 26743 3349 26752 3383
rect 26700 3340 26752 3349
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 15982 3238 16034 3290
rect 16046 3238 16098 3290
rect 16110 3238 16162 3290
rect 16174 3238 16226 3290
rect 25982 3238 26034 3290
rect 26046 3238 26098 3290
rect 26110 3238 26162 3290
rect 26174 3238 26226 3290
rect 2596 3179 2648 3188
rect 2596 3145 2605 3179
rect 2605 3145 2639 3179
rect 2639 3145 2648 3179
rect 2596 3136 2648 3145
rect 4896 3136 4948 3188
rect 5172 3179 5224 3188
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 6552 3111 6604 3120
rect 6552 3077 6561 3111
rect 6561 3077 6595 3111
rect 6595 3077 6604 3111
rect 6552 3068 6604 3077
rect 1676 3000 1728 3052
rect 4344 3000 4396 3052
rect 1860 2932 1912 2984
rect 2504 2932 2556 2984
rect 5264 3000 5316 3052
rect 6920 3000 6972 3052
rect 11060 3136 11112 3188
rect 13176 3179 13228 3188
rect 13176 3145 13185 3179
rect 13185 3145 13219 3179
rect 13219 3145 13228 3179
rect 13176 3136 13228 3145
rect 7564 3068 7616 3120
rect 10784 3068 10836 3120
rect 4988 2932 5040 2984
rect 5724 2975 5776 2984
rect 5724 2941 5733 2975
rect 5733 2941 5767 2975
rect 5767 2941 5776 2975
rect 5724 2932 5776 2941
rect 7104 2932 7156 2984
rect 8760 2932 8812 2984
rect 9496 2975 9548 2984
rect 9496 2941 9530 2975
rect 9530 2941 9548 2975
rect 9496 2932 9548 2941
rect 13176 2932 13228 2984
rect 15844 3136 15896 3188
rect 16672 3136 16724 3188
rect 17592 3136 17644 3188
rect 17776 3179 17828 3188
rect 17776 3145 17785 3179
rect 17785 3145 17819 3179
rect 17819 3145 17828 3179
rect 17776 3136 17828 3145
rect 21364 3136 21416 3188
rect 21456 3068 21508 3120
rect 18604 3000 18656 3052
rect 20076 3000 20128 3052
rect 16672 2975 16724 2984
rect 16672 2941 16681 2975
rect 16681 2941 16715 2975
rect 16715 2941 16724 2975
rect 16672 2932 16724 2941
rect 17776 2932 17828 2984
rect 18880 2975 18932 2984
rect 18880 2941 18889 2975
rect 18889 2941 18923 2975
rect 18923 2941 18932 2975
rect 18880 2932 18932 2941
rect 20168 2975 20220 2984
rect 20168 2941 20177 2975
rect 20177 2941 20211 2975
rect 20211 2941 20220 2975
rect 20168 2932 20220 2941
rect 25412 3136 25464 3188
rect 27344 3179 27396 3188
rect 27344 3145 27353 3179
rect 27353 3145 27387 3179
rect 27387 3145 27396 3179
rect 27344 3136 27396 3145
rect 26332 3068 26384 3120
rect 25320 3043 25372 3052
rect 25320 3009 25329 3043
rect 25329 3009 25363 3043
rect 25363 3009 25372 3043
rect 25320 3000 25372 3009
rect 26424 2975 26476 2984
rect 26424 2941 26433 2975
rect 26433 2941 26467 2975
rect 26467 2941 26476 2975
rect 26424 2932 26476 2941
rect 27436 2932 27488 2984
rect 2044 2864 2096 2916
rect 5540 2864 5592 2916
rect 6920 2864 6972 2916
rect 12072 2864 12124 2916
rect 14924 2864 14976 2916
rect 19156 2907 19208 2916
rect 19156 2873 19165 2907
rect 19165 2873 19199 2907
rect 19199 2873 19208 2907
rect 19156 2864 19208 2873
rect 2872 2839 2924 2848
rect 2872 2805 2881 2839
rect 2881 2805 2915 2839
rect 2915 2805 2924 2839
rect 2872 2796 2924 2805
rect 5172 2796 5224 2848
rect 5816 2796 5868 2848
rect 6828 2839 6880 2848
rect 6828 2805 6837 2839
rect 6837 2805 6871 2839
rect 6871 2805 6880 2839
rect 6828 2796 6880 2805
rect 23848 2839 23900 2848
rect 23848 2805 23857 2839
rect 23857 2805 23891 2839
rect 23891 2805 23900 2839
rect 23848 2796 23900 2805
rect 26608 2839 26660 2848
rect 26608 2805 26617 2839
rect 26617 2805 26651 2839
rect 26651 2805 26660 2839
rect 26608 2796 26660 2805
rect 27712 2839 27764 2848
rect 27712 2805 27721 2839
rect 27721 2805 27755 2839
rect 27755 2805 27764 2839
rect 27712 2796 27764 2805
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 20982 2694 21034 2746
rect 21046 2694 21098 2746
rect 21110 2694 21162 2746
rect 21174 2694 21226 2746
rect 1860 2592 1912 2644
rect 5172 2635 5224 2644
rect 5172 2601 5181 2635
rect 5181 2601 5215 2635
rect 5215 2601 5224 2635
rect 5172 2592 5224 2601
rect 5448 2592 5500 2644
rect 6920 2635 6972 2644
rect 6920 2601 6929 2635
rect 6929 2601 6963 2635
rect 6963 2601 6972 2635
rect 6920 2592 6972 2601
rect 8760 2592 8812 2644
rect 7748 2524 7800 2576
rect 2228 2456 2280 2508
rect 3148 2456 3200 2508
rect 4068 2499 4120 2508
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4068 2456 4120 2465
rect 5632 2456 5684 2508
rect 7288 2499 7340 2508
rect 7288 2465 7297 2499
rect 7297 2465 7331 2499
rect 7331 2465 7340 2499
rect 7288 2456 7340 2465
rect 9680 2456 9732 2508
rect 11060 2499 11112 2508
rect 11060 2465 11069 2499
rect 11069 2465 11103 2499
rect 11103 2465 11112 2499
rect 11060 2456 11112 2465
rect 13728 2592 13780 2644
rect 16396 2635 16448 2644
rect 16396 2601 16405 2635
rect 16405 2601 16439 2635
rect 16439 2601 16448 2635
rect 16396 2592 16448 2601
rect 18604 2635 18656 2644
rect 18604 2601 18613 2635
rect 18613 2601 18647 2635
rect 18647 2601 18656 2635
rect 18604 2592 18656 2601
rect 19984 2635 20036 2644
rect 19984 2601 19993 2635
rect 19993 2601 20027 2635
rect 20027 2601 20036 2635
rect 19984 2592 20036 2601
rect 20168 2592 20220 2644
rect 20812 2592 20864 2644
rect 21272 2592 21324 2644
rect 18236 2524 18288 2576
rect 24676 2524 24728 2576
rect 17868 2456 17920 2508
rect 22284 2499 22336 2508
rect 22284 2465 22293 2499
rect 22293 2465 22327 2499
rect 22327 2465 22336 2499
rect 22284 2456 22336 2465
rect 24032 2499 24084 2508
rect 24032 2465 24041 2499
rect 24041 2465 24075 2499
rect 24075 2465 24084 2499
rect 24032 2456 24084 2465
rect 3516 2388 3568 2440
rect 4896 2388 4948 2440
rect 9956 2431 10008 2440
rect 7196 2320 7248 2372
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 10600 2388 10652 2440
rect 13452 2388 13504 2440
rect 16304 2388 16356 2440
rect 19156 2388 19208 2440
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 23480 2388 23532 2440
rect 24216 2431 24268 2440
rect 24216 2397 24225 2431
rect 24225 2397 24259 2431
rect 24259 2397 24268 2431
rect 24216 2388 24268 2397
rect 20536 2320 20588 2372
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 25872 2295 25924 2304
rect 25872 2261 25881 2295
rect 25881 2261 25915 2295
rect 25915 2261 25924 2295
rect 25872 2252 25924 2261
rect 29184 2252 29236 2304
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 15982 2150 16034 2202
rect 16046 2150 16098 2202
rect 16110 2150 16162 2202
rect 16174 2150 16226 2202
rect 25982 2150 26034 2202
rect 26046 2150 26098 2202
rect 26110 2150 26162 2202
rect 26174 2150 26226 2202
<< metal2 >>
rect 1674 23520 1730 24000
rect 3330 23624 3386 23633
rect 3330 23559 3386 23568
rect 1688 22098 1716 23520
rect 2778 22400 2834 22409
rect 2778 22335 2834 22344
rect 1676 22092 1728 22098
rect 1676 22034 1728 22040
rect 2136 22092 2188 22098
rect 2136 22034 2188 22040
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1492 18760 1544 18766
rect 1492 18702 1544 18708
rect 1504 18358 1532 18702
rect 1780 18426 1808 18770
rect 2042 18728 2098 18737
rect 2042 18663 2098 18672
rect 1768 18420 1820 18426
rect 1768 18362 1820 18368
rect 1492 18352 1544 18358
rect 1492 18294 1544 18300
rect 1504 16046 1532 18294
rect 1676 17740 1728 17746
rect 1676 17682 1728 17688
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 1492 16040 1544 16046
rect 1492 15982 1544 15988
rect 1504 15706 1532 15982
rect 1492 15700 1544 15706
rect 1492 15642 1544 15648
rect 754 15328 810 15337
rect 754 15263 810 15272
rect 768 13870 796 15263
rect 1400 15156 1452 15162
rect 1400 15098 1452 15104
rect 1412 14618 1440 15098
rect 1400 14612 1452 14618
rect 1400 14554 1452 14560
rect 1412 14414 1440 14554
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 756 13864 808 13870
rect 756 13806 808 13812
rect 1400 11280 1452 11286
rect 1400 11222 1452 11228
rect 1412 10606 1440 11222
rect 1596 11121 1624 17478
rect 1688 16794 1716 17682
rect 2056 17338 2084 18663
rect 2044 17332 2096 17338
rect 2044 17274 2096 17280
rect 2056 17134 2084 17274
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1676 15972 1728 15978
rect 1676 15914 1728 15920
rect 1688 15434 1716 15914
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 1676 15428 1728 15434
rect 1676 15370 1728 15376
rect 1780 15162 1808 15642
rect 1768 15156 1820 15162
rect 1768 15098 1820 15104
rect 1676 14544 1728 14550
rect 1676 14486 1728 14492
rect 1688 13802 1716 14486
rect 1676 13796 1728 13802
rect 1676 13738 1728 13744
rect 1688 13530 1716 13738
rect 1872 13530 1900 16934
rect 2044 13728 2096 13734
rect 2044 13670 2096 13676
rect 2056 13530 2084 13670
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 2044 13524 2096 13530
rect 2044 13466 2096 13472
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1860 13388 1912 13394
rect 1860 13330 1912 13336
rect 1688 11778 1716 13330
rect 1872 12646 1900 13330
rect 1860 12640 1912 12646
rect 1858 12608 1860 12617
rect 2044 12640 2096 12646
rect 1912 12608 1914 12617
rect 2044 12582 2096 12588
rect 1858 12543 1914 12552
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1688 11750 1900 11778
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1582 11112 1638 11121
rect 1582 11047 1638 11056
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1584 10464 1636 10470
rect 1582 10432 1584 10441
rect 1636 10432 1638 10441
rect 1582 10367 1638 10376
rect 1780 10198 1808 11494
rect 1768 10192 1820 10198
rect 1768 10134 1820 10140
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1584 9376 1636 9382
rect 1582 9344 1584 9353
rect 1636 9344 1638 9353
rect 1582 9279 1638 9288
rect 1400 8832 1452 8838
rect 1400 8774 1452 8780
rect 1412 7449 1440 8774
rect 1490 8664 1546 8673
rect 1490 8599 1546 8608
rect 1504 8090 1532 8599
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 1596 8129 1624 8502
rect 1582 8120 1638 8129
rect 1492 8084 1544 8090
rect 1582 8055 1638 8064
rect 1492 8026 1544 8032
rect 1398 7440 1454 7449
rect 1398 7375 1454 7384
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1596 6730 1624 6831
rect 1584 6724 1636 6730
rect 1584 6666 1636 6672
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 662 3632 718 3641
rect 662 3567 718 3576
rect 676 480 704 3567
rect 662 0 718 480
rect 1412 377 1440 6054
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 1596 5370 1624 5607
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1582 5128 1638 5137
rect 1582 5063 1638 5072
rect 1596 4826 1624 5063
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1490 4448 1546 4457
rect 1490 4383 1546 4392
rect 1504 3942 1532 4383
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1582 3904 1638 3913
rect 1582 3839 1638 3848
rect 1596 3738 1624 3839
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1688 3058 1716 9862
rect 1780 9110 1808 10134
rect 1768 9104 1820 9110
rect 1768 9046 1820 9052
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1780 7274 1808 7686
rect 1768 7268 1820 7274
rect 1768 7210 1820 7216
rect 1872 6361 1900 11750
rect 1964 11558 1992 12038
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 2056 10282 2084 12582
rect 2148 11801 2176 22034
rect 2318 17912 2374 17921
rect 2318 17847 2374 17856
rect 2332 16969 2360 17847
rect 2318 16960 2374 16969
rect 2318 16895 2374 16904
rect 2686 16960 2742 16969
rect 2686 16895 2742 16904
rect 2700 16726 2728 16895
rect 2688 16720 2740 16726
rect 2688 16662 2740 16668
rect 2700 15706 2728 16662
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2332 13802 2360 13874
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2320 13796 2372 13802
rect 2320 13738 2372 13744
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2424 12782 2452 13126
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2332 12073 2360 12242
rect 2318 12064 2374 12073
rect 2516 12050 2544 13670
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2608 12238 2636 13262
rect 2700 12374 2728 13806
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2318 11999 2374 12008
rect 2424 12022 2544 12050
rect 2332 11898 2360 11999
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2134 11792 2190 11801
rect 2134 11727 2190 11736
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 1964 10266 2084 10282
rect 2148 10266 2176 11494
rect 2240 11354 2268 11494
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2240 10810 2268 11154
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 1964 10260 2096 10266
rect 1964 10254 2044 10260
rect 1964 9178 1992 10254
rect 2044 10202 2096 10208
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2332 10146 2360 10746
rect 2148 10118 2360 10146
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2042 9072 2098 9081
rect 2042 9007 2044 9016
rect 2096 9007 2098 9016
rect 2044 8978 2096 8984
rect 2056 8634 2084 8978
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1964 7449 1992 7890
rect 1950 7440 2006 7449
rect 1950 7375 2006 7384
rect 1964 7002 1992 7375
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 2148 6866 2176 10118
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2332 9722 2360 9998
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 2424 8906 2452 12022
rect 2608 11898 2636 12174
rect 2596 11892 2648 11898
rect 2516 11852 2596 11880
rect 2516 11150 2544 11852
rect 2596 11834 2648 11840
rect 2792 11540 2820 22335
rect 3344 22166 3372 23559
rect 4986 23520 5042 24000
rect 8298 23520 8354 24000
rect 11610 23520 11666 24000
rect 14922 23520 14978 24000
rect 18326 23520 18382 24000
rect 21638 23520 21694 24000
rect 24950 23520 25006 24000
rect 25410 23624 25466 23633
rect 25410 23559 25466 23568
rect 4158 23080 4214 23089
rect 4158 23015 4214 23024
rect 3332 22160 3384 22166
rect 3332 22102 3384 22108
rect 4066 21856 4122 21865
rect 4066 21791 4122 21800
rect 3974 21312 4030 21321
rect 3974 21247 4030 21256
rect 3988 21146 4016 21247
rect 3976 21140 4028 21146
rect 3976 21082 4028 21088
rect 4080 20806 4108 21791
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 3790 20632 3846 20641
rect 3790 20567 3846 20576
rect 3516 20392 3568 20398
rect 3516 20334 3568 20340
rect 3330 20088 3386 20097
rect 3528 20058 3556 20334
rect 3330 20023 3386 20032
rect 3516 20052 3568 20058
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3160 19310 3188 19654
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 3068 18970 3096 19110
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 2962 18864 3018 18873
rect 2962 18799 3018 18808
rect 2872 18624 2924 18630
rect 2872 18566 2924 18572
rect 2884 18358 2912 18566
rect 2872 18352 2924 18358
rect 2872 18294 2924 18300
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2884 17202 2912 17478
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2870 16688 2926 16697
rect 2870 16623 2926 16632
rect 2884 16590 2912 16623
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2884 15706 2912 16526
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2884 13326 2912 14214
rect 2976 13988 3004 18799
rect 3056 18080 3108 18086
rect 3054 18048 3056 18057
rect 3108 18048 3110 18057
rect 3054 17983 3110 17992
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 3160 17134 3188 17478
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 3148 17128 3200 17134
rect 3148 17070 3200 17076
rect 3160 16794 3188 17070
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 3068 16114 3096 16526
rect 3252 16250 3280 17138
rect 3240 16244 3292 16250
rect 3240 16186 3292 16192
rect 3056 16108 3108 16114
rect 3056 16050 3108 16056
rect 2976 13960 3096 13988
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 3068 12617 3096 13960
rect 3344 13569 3372 20023
rect 3516 19994 3568 20000
rect 3700 19372 3752 19378
rect 3700 19314 3752 19320
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3424 18964 3476 18970
rect 3424 18906 3476 18912
rect 3436 18222 3464 18906
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3528 18290 3556 18566
rect 3620 18329 3648 19110
rect 3712 18834 3740 19314
rect 3700 18828 3752 18834
rect 3700 18770 3752 18776
rect 3606 18320 3662 18329
rect 3516 18284 3568 18290
rect 3606 18255 3662 18264
rect 3700 18284 3752 18290
rect 3516 18226 3568 18232
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 3620 17746 3648 18255
rect 3700 18226 3752 18232
rect 3608 17740 3660 17746
rect 3608 17682 3660 17688
rect 3606 17640 3662 17649
rect 3606 17575 3662 17584
rect 3620 17082 3648 17575
rect 3712 17202 3740 18226
rect 3700 17196 3752 17202
rect 3700 17138 3752 17144
rect 3620 17054 3740 17082
rect 3608 15972 3660 15978
rect 3608 15914 3660 15920
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3330 13560 3386 13569
rect 3330 13495 3386 13504
rect 3528 12986 3556 13874
rect 3620 13433 3648 15914
rect 3606 13424 3662 13433
rect 3606 13359 3662 13368
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3054 12608 3110 12617
rect 3054 12543 3110 12552
rect 2872 12368 2924 12374
rect 3160 12345 3188 12786
rect 2872 12310 2924 12316
rect 3146 12336 3202 12345
rect 2700 11529 2820 11540
rect 2700 11520 2834 11529
rect 2700 11512 2778 11520
rect 2700 11218 2728 11512
rect 2778 11455 2834 11464
rect 2778 11248 2834 11257
rect 2688 11212 2740 11218
rect 2778 11183 2834 11192
rect 2688 11154 2740 11160
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2516 10742 2544 11086
rect 2792 11082 2820 11183
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2792 10810 2820 11018
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2504 10736 2556 10742
rect 2504 10678 2556 10684
rect 2686 9888 2742 9897
rect 2686 9823 2742 9832
rect 2700 9382 2728 9823
rect 2884 9654 2912 12310
rect 2964 12300 3016 12306
rect 3146 12271 3202 12280
rect 2964 12242 3016 12248
rect 2976 11558 3004 12242
rect 3160 11762 3188 12271
rect 3528 12238 3556 12786
rect 3620 12753 3648 13359
rect 3606 12744 3662 12753
rect 3606 12679 3662 12688
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3620 12442 3648 12582
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2976 11286 3004 11494
rect 3160 11286 3188 11698
rect 3514 11656 3570 11665
rect 3514 11591 3570 11600
rect 3528 11558 3556 11591
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 2964 11280 3016 11286
rect 2964 11222 3016 11228
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 2976 11121 3004 11222
rect 2962 11112 3018 11121
rect 2962 11047 3018 11056
rect 3160 10606 3188 11222
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3148 10600 3200 10606
rect 3712 10577 3740 17054
rect 3148 10542 3200 10548
rect 3698 10568 3754 10577
rect 3068 10198 3096 10542
rect 3160 10266 3188 10542
rect 3698 10503 3754 10512
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3056 10192 3108 10198
rect 3056 10134 3108 10140
rect 3608 10192 3660 10198
rect 3608 10134 3660 10140
rect 3620 9722 3648 10134
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2964 9648 3016 9654
rect 3148 9648 3200 9654
rect 3016 9608 3096 9636
rect 2964 9590 3016 9596
rect 2962 9480 3018 9489
rect 2962 9415 2964 9424
rect 3016 9415 3018 9424
rect 2964 9386 3016 9392
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 3068 8945 3096 9608
rect 3146 9616 3148 9625
rect 3200 9616 3202 9625
rect 3146 9551 3202 9560
rect 3160 9518 3188 9551
rect 3620 9518 3648 9658
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3054 8936 3110 8945
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2596 8900 2648 8906
rect 3054 8871 3110 8880
rect 2596 8842 2648 8848
rect 2410 8528 2466 8537
rect 2410 8463 2412 8472
rect 2464 8463 2466 8472
rect 2412 8434 2464 8440
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2042 6760 2098 6769
rect 2042 6695 2098 6704
rect 2056 6458 2084 6695
rect 2148 6458 2176 6802
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 1858 6352 1914 6361
rect 1858 6287 1914 6296
rect 2056 6254 2084 6394
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 2226 5536 2282 5545
rect 2226 5471 2282 5480
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2042 4720 2098 4729
rect 2042 4655 2044 4664
rect 2096 4655 2098 4664
rect 2044 4626 2096 4632
rect 2148 4185 2176 4966
rect 2134 4176 2190 4185
rect 2134 4111 2190 4120
rect 2042 4040 2098 4049
rect 2042 3975 2044 3984
rect 2096 3975 2098 3984
rect 2044 3946 2096 3952
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1860 2984 1912 2990
rect 1860 2926 1912 2932
rect 1872 2650 1900 2926
rect 2044 2916 2096 2922
rect 2044 2858 2096 2864
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 1596 1465 1624 2246
rect 1582 1456 1638 1465
rect 1582 1391 1638 1400
rect 2056 480 2084 2858
rect 2240 2514 2268 5471
rect 2608 4690 2636 8842
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2700 6662 2728 7278
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 5778 2728 6598
rect 2884 6186 2912 7142
rect 3804 7041 3832 20567
rect 4068 20324 4120 20330
rect 4068 20266 4120 20272
rect 4080 20097 4108 20266
rect 4066 20088 4122 20097
rect 4066 20023 4122 20032
rect 4172 18902 4200 23015
rect 5000 20369 5028 23520
rect 5956 21788 6252 21808
rect 6012 21786 6036 21788
rect 6092 21786 6116 21788
rect 6172 21786 6196 21788
rect 6034 21734 6036 21786
rect 6098 21734 6110 21786
rect 6172 21734 6174 21786
rect 6012 21732 6036 21734
rect 6092 21732 6116 21734
rect 6172 21732 6196 21734
rect 5956 21712 6252 21732
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 5956 20700 6252 20720
rect 6012 20698 6036 20700
rect 6092 20698 6116 20700
rect 6172 20698 6196 20700
rect 6034 20646 6036 20698
rect 6098 20646 6110 20698
rect 6172 20646 6174 20698
rect 6012 20644 6036 20646
rect 6092 20644 6116 20646
rect 6172 20644 6196 20646
rect 5956 20624 6252 20644
rect 4986 20360 5042 20369
rect 4986 20295 5042 20304
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 4160 18896 4212 18902
rect 4436 18896 4488 18902
rect 4160 18838 4212 18844
rect 4434 18864 4436 18873
rect 4488 18864 4490 18873
rect 4434 18799 4490 18808
rect 4448 18358 4476 18799
rect 4540 18766 4568 18797
rect 4528 18760 4580 18766
rect 4526 18728 4528 18737
rect 4804 18760 4856 18766
rect 4580 18728 4582 18737
rect 4804 18702 4856 18708
rect 4526 18663 4582 18672
rect 4540 18426 4568 18663
rect 4528 18420 4580 18426
rect 4528 18362 4580 18368
rect 4436 18352 4488 18358
rect 4436 18294 4488 18300
rect 4816 18086 4844 18702
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4526 17640 4582 17649
rect 4526 17575 4582 17584
rect 4434 17096 4490 17105
rect 4434 17031 4490 17040
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 4080 16833 4108 16934
rect 4066 16824 4122 16833
rect 4066 16759 4122 16768
rect 4250 16008 4306 16017
rect 4250 15943 4252 15952
rect 4304 15943 4306 15952
rect 4252 15914 4304 15920
rect 4068 15904 4120 15910
rect 3882 15872 3938 15881
rect 4068 15846 4120 15852
rect 3882 15807 3938 15816
rect 3790 7032 3846 7041
rect 3700 6996 3752 7002
rect 3790 6967 3846 6976
rect 3700 6938 3752 6944
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 6254 3648 6598
rect 3712 6322 3740 6938
rect 3896 6934 3924 15807
rect 4080 15706 4108 15846
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4448 15638 4476 17031
rect 4436 15632 4488 15638
rect 4436 15574 4488 15580
rect 4448 15162 4476 15574
rect 4540 15502 4568 17575
rect 4816 16794 4844 18022
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4816 16114 4844 16730
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 4908 15586 4936 20198
rect 6642 20088 6698 20097
rect 6642 20023 6644 20032
rect 6696 20023 6698 20032
rect 6644 19994 6696 20000
rect 5264 19916 5316 19922
rect 5264 19858 5316 19864
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 6736 19916 6788 19922
rect 6736 19858 6788 19864
rect 5276 19514 5304 19858
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 5276 17746 5304 19450
rect 5552 19378 5580 19858
rect 5956 19612 6252 19632
rect 6012 19610 6036 19612
rect 6092 19610 6116 19612
rect 6172 19610 6196 19612
rect 6034 19558 6036 19610
rect 6098 19558 6110 19610
rect 6172 19558 6174 19610
rect 6012 19556 6036 19558
rect 6092 19556 6116 19558
rect 6172 19556 6196 19558
rect 5956 19536 6252 19556
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 5956 18524 6252 18544
rect 6012 18522 6036 18524
rect 6092 18522 6116 18524
rect 6172 18522 6196 18524
rect 6034 18470 6036 18522
rect 6098 18470 6110 18522
rect 6172 18470 6174 18522
rect 6012 18468 6036 18470
rect 6092 18468 6116 18470
rect 6172 18468 6196 18470
rect 5956 18448 6252 18468
rect 5630 18048 5686 18057
rect 5630 17983 5686 17992
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 5276 17134 5304 17682
rect 5368 17338 5396 17682
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 4816 15558 4936 15586
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4252 14544 4304 14550
rect 4252 14486 4304 14492
rect 4066 14104 4122 14113
rect 4264 14074 4292 14486
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4066 14039 4068 14048
rect 4120 14039 4122 14048
rect 4252 14068 4304 14074
rect 4068 14010 4120 14016
rect 4252 14010 4304 14016
rect 4080 13870 4108 14010
rect 4068 13864 4120 13870
rect 4264 13818 4292 14010
rect 4068 13806 4120 13812
rect 4172 13790 4292 13818
rect 4356 13802 4384 14214
rect 4344 13796 4396 13802
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 4080 12782 4108 13126
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 3974 12200 4030 12209
rect 3974 12135 4030 12144
rect 3988 11898 4016 12135
rect 4080 12084 4108 12378
rect 4172 12220 4200 13790
rect 4344 13738 4396 13744
rect 4252 13728 4304 13734
rect 4252 13670 4304 13676
rect 4264 12714 4292 13670
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4250 12608 4306 12617
rect 4250 12543 4306 12552
rect 4264 12322 4292 12543
rect 4356 12442 4384 13126
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4264 12294 4384 12322
rect 4252 12232 4304 12238
rect 4172 12192 4252 12220
rect 4252 12174 4304 12180
rect 4080 12056 4200 12084
rect 4172 11937 4200 12056
rect 4158 11928 4214 11937
rect 3976 11892 4028 11898
rect 4264 11898 4292 12174
rect 4158 11863 4214 11872
rect 4252 11892 4304 11898
rect 3976 11834 4028 11840
rect 3988 11694 4016 11834
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 4172 10282 4200 11863
rect 4252 11834 4304 11840
rect 4172 10254 4292 10282
rect 4264 8634 4292 10254
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4264 8430 4292 8570
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4356 7954 4384 12294
rect 4448 12186 4476 15098
rect 4540 14822 4568 15438
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4540 13190 4568 14758
rect 4816 13938 4844 15558
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 4908 14822 4936 15438
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4908 14618 4936 14758
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 4724 13462 4752 13493
rect 4712 13456 4764 13462
rect 4710 13424 4712 13433
rect 4764 13424 4766 13433
rect 4710 13359 4766 13368
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4724 12986 4752 13359
rect 4816 13326 4844 13874
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4724 12889 4752 12922
rect 4710 12880 4766 12889
rect 4710 12815 4766 12824
rect 4448 12158 4568 12186
rect 4434 12064 4490 12073
rect 4434 11999 4490 12008
rect 4448 11762 4476 11999
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4448 9518 4476 10406
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4540 9178 4568 12158
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4540 8362 4568 9114
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4448 8090 4476 8230
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4080 7002 4108 7686
rect 4356 7546 4384 7890
rect 4448 7546 4476 8026
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 3884 6928 3936 6934
rect 3884 6870 3936 6876
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 2872 6180 2924 6186
rect 2792 6140 2872 6168
rect 2792 5846 2820 6140
rect 2872 6122 2924 6128
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2596 4684 2648 4690
rect 2596 4626 2648 4632
rect 2608 4282 2636 4626
rect 2700 4622 2728 5714
rect 2792 5234 2820 5782
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2884 5370 2912 5510
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2596 4276 2648 4282
rect 2596 4218 2648 4224
rect 2700 4078 2728 4558
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2700 3670 2728 4014
rect 2688 3664 2740 3670
rect 2688 3606 2740 3612
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2502 3496 2558 3505
rect 2502 3431 2558 3440
rect 2516 2990 2544 3431
rect 2608 3194 2636 3538
rect 2688 3392 2740 3398
rect 2792 3369 2820 4422
rect 2884 4078 2912 5306
rect 3252 5234 3280 6054
rect 4080 5370 4108 6326
rect 4356 6118 4384 6802
rect 4540 6769 4568 8298
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4632 7274 4660 7822
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4632 6798 4660 7210
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4620 6792 4672 6798
rect 4526 6760 4582 6769
rect 4620 6734 4672 6740
rect 4526 6695 4582 6704
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2884 3738 2912 4014
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2688 3334 2740 3340
rect 2778 3360 2834 3369
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 2700 2802 2728 3334
rect 2778 3295 2834 3304
rect 2872 2848 2924 2854
rect 2700 2774 2820 2802
rect 2872 2790 2924 2796
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 2792 2145 2820 2774
rect 2884 2689 2912 2790
rect 2870 2680 2926 2689
rect 2870 2615 2926 2624
rect 3160 2514 3188 4966
rect 3252 4826 3280 5170
rect 4080 5098 4108 5306
rect 4356 5273 4384 6054
rect 4632 5914 4660 6734
rect 4724 6118 4752 6802
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4724 5545 4752 6054
rect 4710 5536 4766 5545
rect 4710 5471 4766 5480
rect 4342 5264 4398 5273
rect 4342 5199 4398 5208
rect 4724 5137 4752 5471
rect 4710 5128 4766 5137
rect 4068 5092 4120 5098
rect 4710 5063 4766 5072
rect 4068 5034 4120 5040
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 3976 4004 4028 4010
rect 3976 3946 4028 3952
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 2778 2136 2834 2145
rect 2778 2071 2834 2080
rect 3528 480 3556 2382
rect 3988 921 4016 3946
rect 4356 3738 4384 4218
rect 4632 4214 4660 4558
rect 4908 4282 4936 4626
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4356 3058 4384 3674
rect 4632 3670 4660 4150
rect 5000 3670 5028 16730
rect 5276 16658 5304 17070
rect 5644 16726 5672 17983
rect 5956 17436 6252 17456
rect 6012 17434 6036 17436
rect 6092 17434 6116 17436
rect 6172 17434 6196 17436
rect 6034 17382 6036 17434
rect 6098 17382 6110 17434
rect 6172 17382 6174 17434
rect 6012 17380 6036 17382
rect 6092 17380 6116 17382
rect 6172 17380 6196 17382
rect 5956 17360 6252 17380
rect 5722 16824 5778 16833
rect 5722 16759 5724 16768
rect 5776 16759 5778 16768
rect 5724 16730 5776 16736
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5538 16416 5594 16425
rect 5538 16351 5594 16360
rect 5172 15156 5224 15162
rect 5172 15098 5224 15104
rect 5184 14482 5212 15098
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5184 14074 5212 14418
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5460 14006 5488 14418
rect 5448 14000 5500 14006
rect 5448 13942 5500 13948
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 5092 12918 5120 13330
rect 5080 12912 5132 12918
rect 5078 12880 5080 12889
rect 5132 12880 5134 12889
rect 5078 12815 5134 12824
rect 5184 9926 5212 13806
rect 5460 11898 5488 13942
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5552 10198 5580 16351
rect 5644 16114 5672 16662
rect 5736 16182 5764 16730
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5828 16250 5856 16526
rect 5956 16348 6252 16368
rect 6012 16346 6036 16348
rect 6092 16346 6116 16348
rect 6172 16346 6196 16348
rect 6034 16294 6036 16346
rect 6098 16294 6110 16346
rect 6172 16294 6174 16346
rect 6012 16292 6036 16294
rect 6092 16292 6116 16294
rect 6172 16292 6196 16294
rect 5956 16272 6252 16292
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 5724 16176 5776 16182
rect 5724 16118 5776 16124
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5956 15260 6252 15280
rect 6012 15258 6036 15260
rect 6092 15258 6116 15260
rect 6172 15258 6196 15260
rect 6034 15206 6036 15258
rect 6098 15206 6110 15258
rect 6172 15206 6174 15258
rect 6012 15204 6036 15206
rect 6092 15204 6116 15206
rect 6172 15204 6196 15206
rect 5956 15184 6252 15204
rect 5956 14172 6252 14192
rect 6012 14170 6036 14172
rect 6092 14170 6116 14172
rect 6172 14170 6196 14172
rect 6034 14118 6036 14170
rect 6098 14118 6110 14170
rect 6172 14118 6174 14170
rect 6012 14116 6036 14118
rect 6092 14116 6116 14118
rect 6172 14116 6196 14118
rect 5956 14096 6252 14116
rect 5956 13084 6252 13104
rect 6012 13082 6036 13084
rect 6092 13082 6116 13084
rect 6172 13082 6196 13084
rect 6034 13030 6036 13082
rect 6098 13030 6110 13082
rect 6172 13030 6174 13082
rect 6012 13028 6036 13030
rect 6092 13028 6116 13030
rect 6172 13028 6196 13030
rect 5956 13008 6252 13028
rect 5630 12336 5686 12345
rect 5630 12271 5686 12280
rect 5644 12170 5672 12271
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5956 11996 6252 12016
rect 6012 11994 6036 11996
rect 6092 11994 6116 11996
rect 6172 11994 6196 11996
rect 6034 11942 6036 11994
rect 6098 11942 6110 11994
rect 6172 11942 6174 11994
rect 6012 11940 6036 11942
rect 6092 11940 6116 11942
rect 6172 11940 6196 11942
rect 5956 11920 6252 11940
rect 5956 10908 6252 10928
rect 6012 10906 6036 10908
rect 6092 10906 6116 10908
rect 6172 10906 6196 10908
rect 6034 10854 6036 10906
rect 6098 10854 6110 10906
rect 6172 10854 6174 10906
rect 6012 10852 6036 10854
rect 6092 10852 6116 10854
rect 6172 10852 6196 10854
rect 5956 10832 6252 10852
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 6288 9994 6316 10406
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 5092 5914 5120 6190
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 5184 3738 5212 9862
rect 5956 9820 6252 9840
rect 6012 9818 6036 9820
rect 6092 9818 6116 9820
rect 6172 9818 6196 9820
rect 6034 9766 6036 9818
rect 6098 9766 6110 9818
rect 6172 9766 6174 9818
rect 6012 9764 6036 9766
rect 6092 9764 6116 9766
rect 6172 9764 6196 9766
rect 5956 9744 6252 9764
rect 6288 9722 6316 9930
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6564 9625 6592 19110
rect 6748 18902 6776 19858
rect 6920 19780 6972 19786
rect 6920 19722 6972 19728
rect 6932 19666 6960 19722
rect 6840 19638 6960 19666
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 6736 18896 6788 18902
rect 6736 18838 6788 18844
rect 6840 18426 6868 19638
rect 7208 19174 7236 19654
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 7116 18154 7144 19110
rect 7208 18970 7236 19110
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 7196 18624 7248 18630
rect 7196 18566 7248 18572
rect 7208 18290 7236 18566
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 7104 18148 7156 18154
rect 7104 18090 7156 18096
rect 7116 17882 7144 18090
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7116 16658 7144 17478
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 6840 16266 6868 16594
rect 6840 16238 6960 16266
rect 7116 16250 7144 16594
rect 6840 15162 6868 16238
rect 6932 16182 6960 16238
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6840 13530 6868 15098
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7024 13734 7052 13806
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 7024 13530 7052 13670
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 6840 12850 6868 13466
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6748 11082 6776 12650
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6932 11762 6960 12038
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6748 10742 6776 11018
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 6748 10266 6776 10678
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6550 9616 6606 9625
rect 6550 9551 6606 9560
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5368 8838 5396 9386
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5630 9344 5686 9353
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5368 7886 5396 8774
rect 5552 8498 5580 9318
rect 5630 9279 5686 9288
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5552 8022 5580 8434
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5368 7342 5396 7822
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5460 6322 5488 6598
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5552 6202 5580 7414
rect 5460 6186 5580 6202
rect 5448 6180 5580 6186
rect 5500 6174 5580 6180
rect 5448 6122 5500 6128
rect 5460 5914 5488 6122
rect 5644 6066 5672 9279
rect 5956 8732 6252 8752
rect 6012 8730 6036 8732
rect 6092 8730 6116 8732
rect 6172 8730 6196 8732
rect 6034 8678 6036 8730
rect 6098 8678 6110 8730
rect 6172 8678 6174 8730
rect 6012 8676 6036 8678
rect 6092 8676 6116 8678
rect 6172 8676 6196 8678
rect 5956 8656 6252 8676
rect 5724 8016 5776 8022
rect 5724 7958 5776 7964
rect 5736 7546 5764 7958
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 5956 7644 6252 7664
rect 6012 7642 6036 7644
rect 6092 7642 6116 7644
rect 6172 7642 6196 7644
rect 6034 7590 6036 7642
rect 6098 7590 6110 7642
rect 6172 7590 6174 7642
rect 6012 7588 6036 7590
rect 6092 7588 6116 7590
rect 6172 7588 6196 7590
rect 5956 7568 6252 7588
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 6380 7274 6408 7686
rect 6642 7440 6698 7449
rect 6642 7375 6698 7384
rect 6656 7342 6684 7375
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6368 7268 6420 7274
rect 6368 7210 6420 7216
rect 5814 7032 5870 7041
rect 5814 6967 5870 6976
rect 6182 7032 6238 7041
rect 6182 6967 6184 6976
rect 5828 6458 5856 6967
rect 6236 6967 6238 6976
rect 6184 6938 6236 6944
rect 6380 6798 6408 7210
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 5956 6556 6252 6576
rect 6012 6554 6036 6556
rect 6092 6554 6116 6556
rect 6172 6554 6196 6556
rect 6034 6502 6036 6554
rect 6098 6502 6110 6554
rect 6172 6502 6174 6554
rect 6012 6500 6036 6502
rect 6092 6500 6116 6502
rect 6172 6500 6196 6502
rect 5956 6480 6252 6500
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 6288 6225 6316 6734
rect 6274 6216 6330 6225
rect 6274 6151 6330 6160
rect 5552 6038 5672 6066
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4988 3664 5040 3670
rect 4988 3606 5040 3612
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4908 3194 4936 3334
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 5000 2990 5028 3606
rect 5184 3194 5212 3674
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5276 3058 5304 4014
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5172 2848 5224 2854
rect 4066 2816 4122 2825
rect 5172 2790 5224 2796
rect 4066 2751 4122 2760
rect 4080 2514 4108 2751
rect 5184 2650 5212 2790
rect 5460 2650 5488 3334
rect 5552 2922 5580 6038
rect 6288 5914 6316 6151
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 5956 5468 6252 5488
rect 6012 5466 6036 5468
rect 6092 5466 6116 5468
rect 6172 5466 6196 5468
rect 6034 5414 6036 5466
rect 6098 5414 6110 5466
rect 6172 5414 6174 5466
rect 6012 5412 6036 5414
rect 6092 5412 6116 5414
rect 6172 5412 6196 5414
rect 5956 5392 6252 5412
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5828 4486 5856 4966
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5644 2514 5672 3674
rect 5828 3534 5856 4422
rect 5956 4380 6252 4400
rect 6012 4378 6036 4380
rect 6092 4378 6116 4380
rect 6172 4378 6196 4380
rect 6034 4326 6036 4378
rect 6098 4326 6110 4378
rect 6172 4326 6174 4378
rect 6012 4324 6036 4326
rect 6092 4324 6116 4326
rect 6172 4324 6196 4326
rect 5956 4304 6252 4324
rect 6288 3602 6316 5850
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6656 4049 6684 5306
rect 6642 4040 6698 4049
rect 6642 3975 6698 3984
rect 6840 3738 6868 11494
rect 6932 11354 6960 11698
rect 7196 11552 7248 11558
rect 7194 11520 7196 11529
rect 7248 11520 7250 11529
rect 7194 11455 7250 11464
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6932 10810 6960 11154
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6932 10266 6960 10746
rect 7024 10538 7052 11086
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 7024 10266 7052 10474
rect 7300 10441 7328 21082
rect 7564 20800 7616 20806
rect 7564 20742 7616 20748
rect 7576 18970 7604 20742
rect 8312 20618 8340 23520
rect 10956 21244 11252 21264
rect 11012 21242 11036 21244
rect 11092 21242 11116 21244
rect 11172 21242 11196 21244
rect 11034 21190 11036 21242
rect 11098 21190 11110 21242
rect 11172 21190 11174 21242
rect 11012 21188 11036 21190
rect 11092 21188 11116 21190
rect 11172 21188 11196 21190
rect 10956 21168 11252 21188
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8220 20602 8340 20618
rect 8208 20596 8340 20602
rect 8260 20590 8340 20596
rect 8208 20538 8260 20544
rect 8404 20398 8432 20742
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 7746 19816 7802 19825
rect 7746 19751 7748 19760
rect 7800 19751 7802 19760
rect 7748 19722 7800 19728
rect 7852 19666 7880 20198
rect 8024 19984 8076 19990
rect 8024 19926 8076 19932
rect 7760 19638 7880 19666
rect 7760 19378 7788 19638
rect 8036 19514 8064 19926
rect 8404 19922 8432 20334
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 8024 19508 8076 19514
rect 8024 19450 8076 19456
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 7380 18896 7432 18902
rect 7380 18838 7432 18844
rect 7392 18290 7420 18838
rect 7576 18426 7604 18906
rect 7760 18766 7788 19314
rect 8114 19272 8170 19281
rect 8114 19207 8116 19216
rect 8168 19207 8170 19216
rect 8220 19224 8248 19790
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8760 19372 8812 19378
rect 8760 19314 8812 19320
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8300 19236 8352 19242
rect 8220 19196 8300 19224
rect 8116 19178 8168 19184
rect 8300 19178 8352 19184
rect 8312 18970 8340 19178
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8404 18850 8432 19246
rect 8772 18902 8800 19314
rect 8864 19310 8892 19654
rect 9692 19378 9720 20198
rect 10956 20156 11252 20176
rect 11012 20154 11036 20156
rect 11092 20154 11116 20156
rect 11172 20154 11196 20156
rect 11034 20102 11036 20154
rect 11098 20102 11110 20154
rect 11172 20102 11174 20154
rect 11012 20100 11036 20102
rect 11092 20100 11116 20102
rect 11172 20100 11196 20102
rect 10956 20080 11252 20100
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 10692 19916 10744 19922
rect 10744 19876 10824 19904
rect 10692 19858 10744 19864
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 10796 19174 10824 19876
rect 10980 19310 11008 19926
rect 11624 19922 11652 23520
rect 12072 22160 12124 22166
rect 12072 22102 12124 22108
rect 11612 19916 11664 19922
rect 11612 19858 11664 19864
rect 11428 19712 11480 19718
rect 11428 19654 11480 19660
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 10600 19168 10652 19174
rect 10600 19110 10652 19116
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 8220 18822 8432 18850
rect 8760 18896 8812 18902
rect 8760 18838 8812 18844
rect 7656 18760 7708 18766
rect 7654 18728 7656 18737
rect 7748 18760 7800 18766
rect 7708 18728 7710 18737
rect 7748 18702 7800 18708
rect 7654 18663 7710 18672
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7576 18193 7604 18362
rect 7562 18184 7618 18193
rect 7562 18119 7618 18128
rect 7668 17814 7696 18663
rect 7760 18358 7788 18702
rect 7748 18352 7800 18358
rect 7748 18294 7800 18300
rect 8220 17882 8248 18822
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 7656 17808 7708 17814
rect 7656 17750 7708 17756
rect 8022 17776 8078 17785
rect 8022 17711 8024 17720
rect 8076 17711 8078 17720
rect 8024 17682 8076 17688
rect 8036 16998 8064 17682
rect 8588 17678 8616 18702
rect 9324 18630 9352 19110
rect 10612 18766 10640 19110
rect 10956 19068 11252 19088
rect 11012 19066 11036 19068
rect 11092 19066 11116 19068
rect 11172 19066 11196 19068
rect 11034 19014 11036 19066
rect 11098 19014 11110 19066
rect 11172 19014 11174 19066
rect 11012 19012 11036 19014
rect 11092 19012 11116 19014
rect 11172 19012 11196 19014
rect 10956 18992 11252 19012
rect 11440 18902 11468 19654
rect 11794 19408 11850 19417
rect 11794 19343 11796 19352
rect 11848 19343 11850 19352
rect 11796 19314 11848 19320
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 11428 18896 11480 18902
rect 11428 18838 11480 18844
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9772 18624 9824 18630
rect 9772 18566 9824 18572
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 9784 18426 9812 18566
rect 9772 18420 9824 18426
rect 9772 18362 9824 18368
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9600 17678 9628 18226
rect 9968 18222 9996 18566
rect 10428 18290 10456 18566
rect 10416 18284 10468 18290
rect 10416 18226 10468 18232
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 8496 17338 8524 17614
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8588 17202 8616 17614
rect 9496 17264 9548 17270
rect 9496 17206 9548 17212
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 9508 17105 9536 17206
rect 9494 17096 9550 17105
rect 9494 17031 9550 17040
rect 8024 16992 8076 16998
rect 8022 16960 8024 16969
rect 8076 16960 8078 16969
rect 8022 16895 8078 16904
rect 9968 16794 9996 18158
rect 10324 18148 10376 18154
rect 10324 18090 10376 18096
rect 10336 17882 10364 18090
rect 10612 18086 10640 18702
rect 10888 18426 10916 18838
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 10704 17513 10732 17682
rect 10888 17678 10916 18362
rect 10956 17980 11252 18000
rect 11012 17978 11036 17980
rect 11092 17978 11116 17980
rect 11172 17978 11196 17980
rect 11034 17926 11036 17978
rect 11098 17926 11110 17978
rect 11172 17926 11174 17978
rect 11012 17924 11036 17926
rect 11092 17924 11116 17926
rect 11172 17924 11196 17926
rect 10956 17904 11252 17924
rect 10784 17672 10836 17678
rect 10782 17640 10784 17649
rect 10876 17672 10928 17678
rect 10836 17640 10838 17649
rect 10876 17614 10928 17620
rect 10782 17575 10838 17584
rect 10690 17504 10746 17513
rect 10690 17439 10746 17448
rect 10704 17270 10732 17439
rect 10692 17264 10744 17270
rect 10692 17206 10744 17212
rect 10796 17066 10824 17575
rect 10888 17338 10916 17614
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9864 16720 9916 16726
rect 9862 16688 9864 16697
rect 9916 16688 9918 16697
rect 9862 16623 9918 16632
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7668 15026 7696 15302
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7484 13938 7512 14350
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7484 13410 7512 13874
rect 7852 13870 7880 14418
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7562 13424 7618 13433
rect 7484 13382 7562 13410
rect 7562 13359 7618 13368
rect 7576 10792 7604 13359
rect 7852 13138 7880 13806
rect 7944 13258 7972 15098
rect 8220 14958 8248 16390
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8312 15162 8340 15506
rect 8864 15366 8892 15982
rect 9036 15972 9088 15978
rect 9036 15914 9088 15920
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8220 14414 8248 14894
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 8036 13938 8064 14214
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 8116 13728 8168 13734
rect 8116 13670 8168 13676
rect 7932 13252 7984 13258
rect 7932 13194 7984 13200
rect 7930 13152 7986 13161
rect 7852 13110 7930 13138
rect 7930 13087 7986 13096
rect 7944 12889 7972 13087
rect 8128 12889 8156 13670
rect 8220 13530 8248 14350
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8404 12986 8432 13330
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 7930 12880 7986 12889
rect 7930 12815 7986 12824
rect 8114 12880 8170 12889
rect 8114 12815 8170 12824
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 7392 10764 7604 10792
rect 7286 10432 7342 10441
rect 7286 10367 7342 10376
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7116 8634 7144 8978
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7208 7290 7236 9522
rect 7392 9518 7420 10764
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7472 10600 7524 10606
rect 7470 10568 7472 10577
rect 7524 10568 7526 10577
rect 7470 10503 7526 10512
rect 7472 10192 7524 10198
rect 7470 10160 7472 10169
rect 7524 10160 7526 10169
rect 7470 10095 7526 10104
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7286 7576 7342 7585
rect 7286 7511 7342 7520
rect 7300 7342 7328 7511
rect 7392 7410 7420 7686
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7116 7262 7236 7290
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6932 5370 6960 5646
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 7024 4826 7052 5510
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7116 4570 7144 7262
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7208 6866 7236 7142
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7300 6254 7328 6598
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7300 5234 7328 6190
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7392 4690 7420 6054
rect 7484 5896 7512 10095
rect 7576 9994 7604 10610
rect 7852 10470 7880 10950
rect 7944 10554 7972 12815
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8220 11830 8248 12582
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 8496 11762 8524 15302
rect 9048 15162 9076 15914
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9600 15178 9628 15506
rect 9600 15162 9720 15178
rect 9036 15156 9088 15162
rect 9600 15156 9732 15162
rect 9600 15150 9680 15156
rect 9036 15098 9088 15104
rect 9680 15098 9732 15104
rect 9048 14090 9076 15098
rect 10244 14657 10272 17002
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10336 16454 10364 16934
rect 10888 16590 10916 17274
rect 10956 16892 11252 16912
rect 11012 16890 11036 16892
rect 11092 16890 11116 16892
rect 11172 16890 11196 16892
rect 11034 16838 11036 16890
rect 11098 16838 11110 16890
rect 11172 16838 11174 16890
rect 11012 16836 11036 16838
rect 11092 16836 11116 16838
rect 11172 16836 11196 16838
rect 10956 16816 11252 16836
rect 11334 16824 11390 16833
rect 11334 16759 11390 16768
rect 11060 16720 11112 16726
rect 11348 16708 11376 16759
rect 11112 16680 11376 16708
rect 11060 16662 11112 16668
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10888 15706 10916 16526
rect 10980 16017 11008 16594
rect 11072 16250 11100 16662
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11336 16176 11388 16182
rect 11336 16118 11388 16124
rect 10966 16008 11022 16017
rect 10966 15943 10968 15952
rect 11020 15943 11022 15952
rect 10968 15914 11020 15920
rect 10956 15804 11252 15824
rect 11012 15802 11036 15804
rect 11092 15802 11116 15804
rect 11172 15802 11196 15804
rect 11034 15750 11036 15802
rect 11098 15750 11110 15802
rect 11172 15750 11174 15802
rect 11012 15748 11036 15750
rect 11092 15748 11116 15750
rect 11172 15748 11196 15750
rect 10956 15728 11252 15748
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 11348 15638 11376 16118
rect 11336 15632 11388 15638
rect 11336 15574 11388 15580
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11256 15162 11284 15438
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11348 14822 11376 15574
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 10956 14716 11252 14736
rect 11012 14714 11036 14716
rect 11092 14714 11116 14716
rect 11172 14714 11196 14716
rect 11034 14662 11036 14714
rect 11098 14662 11110 14714
rect 11172 14662 11174 14714
rect 11012 14660 11036 14662
rect 11092 14660 11116 14662
rect 11172 14660 11196 14662
rect 10230 14648 10286 14657
rect 10956 14640 11252 14660
rect 10230 14583 10286 14592
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 8956 14074 9076 14090
rect 8944 14068 9076 14074
rect 8996 14062 9076 14068
rect 8944 14010 8996 14016
rect 9036 14000 9088 14006
rect 9036 13942 9088 13948
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8588 13297 8616 13738
rect 9048 13530 9076 13942
rect 9232 13870 9260 14214
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9600 13818 9628 14010
rect 9678 13968 9734 13977
rect 9678 13903 9680 13912
rect 9732 13903 9734 13912
rect 9680 13874 9732 13880
rect 9772 13864 9824 13870
rect 9232 13530 9260 13806
rect 9600 13790 9720 13818
rect 9772 13806 9824 13812
rect 9954 13832 10010 13841
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 8574 13288 8630 13297
rect 9692 13258 9720 13790
rect 8574 13223 8630 13232
rect 9680 13252 9732 13258
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8312 10674 8340 11494
rect 8496 11354 8524 11698
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 7944 10526 8064 10554
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7930 10432 7986 10441
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7564 9988 7616 9994
rect 7564 9930 7616 9936
rect 7668 9722 7696 9998
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 7564 9376 7616 9382
rect 7562 9344 7564 9353
rect 7616 9344 7618 9353
rect 7562 9279 7618 9288
rect 7668 9178 7696 9658
rect 7760 9450 7788 10134
rect 7852 9722 7880 10406
rect 7930 10367 7986 10376
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7838 9480 7894 9489
rect 7748 9444 7800 9450
rect 7838 9415 7894 9424
rect 7748 9386 7800 9392
rect 7760 9178 7788 9386
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7668 6118 7696 6258
rect 7852 6254 7880 9415
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7484 5868 7604 5896
rect 7470 5808 7526 5817
rect 7470 5743 7472 5752
rect 7524 5743 7526 5752
rect 7472 5714 7524 5720
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7024 4542 7144 4570
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7024 4146 7052 4542
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 5724 2984 5776 2990
rect 5722 2952 5724 2961
rect 5776 2952 5778 2961
rect 5722 2887 5778 2896
rect 5828 2854 5856 3470
rect 5956 3292 6252 3312
rect 6012 3290 6036 3292
rect 6092 3290 6116 3292
rect 6172 3290 6196 3292
rect 6034 3238 6036 3290
rect 6098 3238 6110 3290
rect 6172 3238 6174 3290
rect 6012 3236 6036 3238
rect 6092 3236 6116 3238
rect 6172 3236 6196 3238
rect 5956 3216 6252 3236
rect 6564 3126 6592 3470
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6932 3058 6960 3334
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7116 2990 7144 4422
rect 7208 4282 7236 4558
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 6920 2916 6972 2922
rect 6920 2858 6972 2864
rect 5816 2848 5868 2854
rect 6828 2848 6880 2854
rect 5816 2790 5868 2796
rect 6826 2816 6828 2825
rect 6880 2816 6882 2825
rect 6826 2751 6882 2760
rect 6932 2650 6960 2858
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 3974 912 4030 921
rect 3974 847 4030 856
rect 4908 480 4936 2382
rect 7208 2378 7236 4218
rect 7392 4214 7420 4626
rect 7484 4282 7512 4762
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7576 3738 7604 5868
rect 7668 5710 7696 6054
rect 7748 5840 7800 5846
rect 7944 5828 7972 10367
rect 8036 9586 8064 10526
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8036 9382 8064 9522
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8128 9178 8156 9862
rect 8404 9602 8432 9862
rect 8312 9586 8432 9602
rect 8300 9580 8432 9586
rect 8352 9574 8432 9580
rect 8300 9522 8352 9528
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8036 8294 8064 8978
rect 8128 8634 8156 9114
rect 8404 8974 8432 9574
rect 8496 9110 8524 9862
rect 8588 9761 8616 13223
rect 9680 13194 9732 13200
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 8864 12345 8892 12922
rect 9680 12640 9732 12646
rect 9678 12608 9680 12617
rect 9732 12608 9734 12617
rect 9678 12543 9734 12552
rect 8850 12336 8906 12345
rect 8850 12271 8906 12280
rect 8864 10130 8892 12271
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9678 11520 9734 11529
rect 9600 11098 9628 11494
rect 9678 11455 9734 11464
rect 9692 11354 9720 11455
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9600 11082 9720 11098
rect 9600 11076 9732 11082
rect 9600 11070 9680 11076
rect 9600 10742 9628 11070
rect 9680 11018 9732 11024
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8574 9752 8630 9761
rect 8574 9687 8630 9696
rect 8574 9616 8630 9625
rect 8574 9551 8630 9560
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8588 9042 8616 9551
rect 8864 9178 8892 10066
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 9600 9042 9628 9862
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8404 8634 8432 8910
rect 9692 8906 9720 9318
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 7800 5800 7972 5828
rect 7748 5782 7800 5788
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7668 5098 7696 5646
rect 7760 5409 7788 5782
rect 7746 5400 7802 5409
rect 7746 5335 7748 5344
rect 7800 5335 7802 5344
rect 7748 5306 7800 5312
rect 7656 5092 7708 5098
rect 7656 5034 7708 5040
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7300 2514 7328 3334
rect 7576 3126 7604 3674
rect 8036 3602 8064 8230
rect 9324 7342 9352 8230
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 8772 6662 8800 7278
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8128 4826 8156 5102
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8128 4146 8156 4762
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 8772 3534 8800 6598
rect 9600 6322 9628 7210
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9600 5914 9628 6258
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9508 4622 9536 4966
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9402 3632 9458 3641
rect 9402 3567 9458 3576
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 7564 3120 7616 3126
rect 7564 3062 7616 3068
rect 8772 2990 8800 3470
rect 8760 2984 8812 2990
rect 9416 2961 9444 3567
rect 9508 2990 9536 4558
rect 9496 2984 9548 2990
rect 8760 2926 8812 2932
rect 9218 2952 9274 2961
rect 8772 2650 8800 2926
rect 9218 2887 9274 2896
rect 9402 2952 9458 2961
rect 9496 2926 9548 2932
rect 9402 2887 9458 2896
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7196 2372 7248 2378
rect 7196 2314 7248 2320
rect 5956 2204 6252 2224
rect 6012 2202 6036 2204
rect 6092 2202 6116 2204
rect 6172 2202 6196 2204
rect 6034 2150 6036 2202
rect 6098 2150 6110 2202
rect 6172 2150 6174 2202
rect 6012 2148 6036 2150
rect 6092 2148 6116 2150
rect 6172 2148 6196 2150
rect 5956 2128 6252 2148
rect 6366 1456 6422 1465
rect 6366 1391 6422 1400
rect 6380 480 6408 1391
rect 7760 480 7788 2518
rect 9232 480 9260 2887
rect 9692 2514 9720 6598
rect 9784 2553 9812 13806
rect 9954 13767 10010 13776
rect 9864 10464 9916 10470
rect 9862 10432 9864 10441
rect 9916 10432 9918 10441
rect 9862 10367 9918 10376
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9876 9382 9904 9454
rect 9968 9450 9996 13767
rect 10140 13320 10192 13326
rect 10138 13288 10140 13297
rect 10192 13288 10194 13297
rect 10138 13223 10194 13232
rect 10046 13152 10102 13161
rect 10046 13087 10102 13096
rect 10060 12782 10088 13087
rect 10152 12850 10180 13223
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10152 10810 10180 11086
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10048 10532 10100 10538
rect 10048 10474 10100 10480
rect 10060 9926 10088 10474
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9876 8945 9904 9318
rect 9862 8936 9918 8945
rect 9862 8871 9918 8880
rect 9876 3097 9904 8871
rect 10060 4185 10088 9862
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10152 7546 10180 8298
rect 10244 7698 10272 14583
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 11072 14362 11100 14418
rect 11348 14414 11376 14758
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 10888 14334 11100 14362
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11152 14340 11204 14346
rect 10506 13560 10562 13569
rect 10888 13530 10916 14334
rect 11152 14282 11204 14288
rect 11164 13870 11192 14282
rect 11348 13977 11376 14350
rect 11624 14074 11652 14418
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11334 13968 11390 13977
rect 11334 13903 11390 13912
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 10956 13628 11252 13648
rect 11012 13626 11036 13628
rect 11092 13626 11116 13628
rect 11172 13626 11196 13628
rect 11034 13574 11036 13626
rect 11098 13574 11110 13626
rect 11172 13574 11174 13626
rect 11012 13572 11036 13574
rect 11092 13572 11116 13574
rect 11172 13572 11196 13574
rect 10956 13552 11252 13572
rect 11348 13530 11376 13903
rect 11612 13796 11664 13802
rect 11612 13738 11664 13744
rect 10506 13495 10562 13504
rect 10876 13524 10928 13530
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10322 13152 10378 13161
rect 10322 13087 10378 13096
rect 10336 12889 10364 13087
rect 10428 12986 10456 13194
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10520 12889 10548 13495
rect 10876 13466 10928 13472
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11624 13326 11652 13738
rect 11716 13530 11744 14486
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 12084 13462 12112 22102
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13556 20398 13584 20742
rect 14936 20505 14964 23520
rect 15956 21788 16252 21808
rect 16012 21786 16036 21788
rect 16092 21786 16116 21788
rect 16172 21786 16196 21788
rect 16034 21734 16036 21786
rect 16098 21734 16110 21786
rect 16172 21734 16174 21786
rect 16012 21732 16036 21734
rect 16092 21732 16116 21734
rect 16172 21732 16196 21734
rect 15956 21712 16252 21732
rect 17040 20936 17092 20942
rect 17040 20878 17092 20884
rect 15956 20700 16252 20720
rect 16012 20698 16036 20700
rect 16092 20698 16116 20700
rect 16172 20698 16196 20700
rect 16034 20646 16036 20698
rect 16098 20646 16110 20698
rect 16172 20646 16174 20698
rect 16012 20644 16036 20646
rect 16092 20644 16116 20646
rect 16172 20644 16196 20646
rect 15956 20624 16252 20644
rect 14922 20496 14978 20505
rect 14922 20431 14978 20440
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 13544 20392 13596 20398
rect 13544 20334 13596 20340
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 12346 18864 12402 18873
rect 12346 18799 12402 18808
rect 12360 18698 12388 18799
rect 12348 18692 12400 18698
rect 12348 18634 12400 18640
rect 12348 18080 12400 18086
rect 12452 18068 12480 20334
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 15108 20256 15160 20262
rect 15160 20204 15240 20210
rect 15108 20198 15240 20204
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13096 19514 13124 19994
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 12400 18040 12480 18068
rect 12348 18022 12400 18028
rect 12360 16590 12388 18022
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12360 15162 12388 16526
rect 12544 16402 12572 16594
rect 12452 16374 12572 16402
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12452 15910 12480 16374
rect 12728 16153 12756 16390
rect 12714 16144 12770 16153
rect 12636 16102 12714 16130
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12452 15366 12480 15846
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12452 13938 12480 15302
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12162 13560 12218 13569
rect 12162 13495 12164 13504
rect 12216 13495 12218 13504
rect 12164 13466 12216 13472
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10322 12880 10378 12889
rect 10322 12815 10378 12824
rect 10506 12880 10562 12889
rect 10506 12815 10562 12824
rect 10796 12617 10824 13194
rect 11624 12986 11652 13262
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 12084 12918 12112 13398
rect 12176 12986 12204 13466
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12072 12912 12124 12918
rect 11334 12880 11390 12889
rect 11334 12815 11390 12824
rect 11992 12860 12072 12866
rect 11992 12854 12124 12860
rect 11992 12838 12112 12854
rect 11348 12617 11376 12815
rect 10782 12608 10838 12617
rect 11334 12608 11390 12617
rect 10782 12543 10838 12552
rect 10956 12540 11252 12560
rect 11334 12543 11390 12552
rect 11012 12538 11036 12540
rect 11092 12538 11116 12540
rect 11172 12538 11196 12540
rect 11034 12486 11036 12538
rect 11098 12486 11110 12538
rect 11172 12486 11174 12538
rect 11012 12484 11036 12486
rect 11092 12484 11116 12486
rect 11172 12484 11196 12486
rect 10956 12464 11252 12484
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10336 11218 10364 12038
rect 10428 11558 10456 12174
rect 10612 11898 10640 12242
rect 10784 12232 10836 12238
rect 10704 12192 10784 12220
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10428 10146 10456 11494
rect 10704 11014 10732 12192
rect 10784 12174 10836 12180
rect 10956 11452 11252 11472
rect 11012 11450 11036 11452
rect 11092 11450 11116 11452
rect 11172 11450 11196 11452
rect 11034 11398 11036 11450
rect 11098 11398 11110 11450
rect 11172 11398 11174 11450
rect 11012 11396 11036 11398
rect 11092 11396 11116 11398
rect 11172 11396 11196 11398
rect 10956 11376 11252 11396
rect 10968 11212 11020 11218
rect 11020 11172 11100 11200
rect 10968 11154 11020 11160
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10598 10704 10654 10713
rect 10704 10674 10732 10950
rect 11072 10810 11100 11172
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10598 10639 10654 10648
rect 10692 10668 10744 10674
rect 10612 10538 10640 10639
rect 10692 10610 10744 10616
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10956 10364 11252 10384
rect 11012 10362 11036 10364
rect 11092 10362 11116 10364
rect 11172 10362 11196 10364
rect 11034 10310 11036 10362
rect 11098 10310 11110 10362
rect 11172 10310 11174 10362
rect 11012 10308 11036 10310
rect 11092 10308 11116 10310
rect 11172 10308 11196 10310
rect 10956 10288 11252 10308
rect 11900 10266 11928 10610
rect 11992 10441 12020 12838
rect 12176 11257 12204 12922
rect 12544 12209 12572 13942
rect 12530 12200 12586 12209
rect 12530 12135 12586 12144
rect 12162 11248 12218 11257
rect 12162 11183 12218 11192
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 11978 10432 12034 10441
rect 11978 10367 12034 10376
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 10336 10118 10456 10146
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 10336 9489 10364 10118
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10322 9480 10378 9489
rect 10428 9450 10456 9998
rect 10704 9586 10732 10134
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10322 9415 10378 9424
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10428 8838 10456 9386
rect 10704 9382 10732 9522
rect 12452 9518 12480 11086
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10428 8430 10456 8774
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10520 8090 10548 8978
rect 10704 8634 10732 9318
rect 10956 9276 11252 9296
rect 11012 9274 11036 9276
rect 11092 9274 11116 9276
rect 11172 9274 11196 9276
rect 11034 9222 11036 9274
rect 11098 9222 11110 9274
rect 11172 9222 11174 9274
rect 11012 9220 11036 9222
rect 11092 9220 11116 9222
rect 11172 9220 11196 9222
rect 10956 9200 11252 9220
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10956 8188 11252 8208
rect 11012 8186 11036 8188
rect 11092 8186 11116 8188
rect 11172 8186 11196 8188
rect 11034 8134 11036 8186
rect 11098 8134 11110 8186
rect 11172 8134 11174 8186
rect 11012 8132 11036 8134
rect 11092 8132 11116 8134
rect 11172 8132 11196 8134
rect 10956 8112 11252 8132
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 10244 7670 10364 7698
rect 10140 7540 10192 7546
rect 10192 7500 10272 7528
rect 10140 7482 10192 7488
rect 10244 6798 10272 7500
rect 10336 6905 10364 7670
rect 11440 7342 11468 7822
rect 11532 7546 11560 7890
rect 12452 7546 12480 9454
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 10956 7100 11252 7120
rect 11012 7098 11036 7100
rect 11092 7098 11116 7100
rect 11172 7098 11196 7100
rect 11034 7046 11036 7098
rect 11098 7046 11110 7098
rect 11172 7046 11174 7098
rect 11012 7044 11036 7046
rect 11092 7044 11116 7046
rect 11172 7044 11196 7046
rect 10956 7024 11252 7044
rect 11532 6934 11560 7482
rect 12164 7200 12216 7206
rect 12162 7168 12164 7177
rect 12216 7168 12218 7177
rect 12162 7103 12218 7112
rect 11520 6928 11572 6934
rect 10322 6896 10378 6905
rect 11520 6870 11572 6876
rect 10322 6831 10378 6840
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10152 6458 10180 6734
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10244 6390 10272 6734
rect 11072 6662 11100 6802
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 6458 11100 6598
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10336 5914 10364 6054
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10704 4826 10732 5850
rect 10796 5370 10824 6122
rect 10956 6012 11252 6032
rect 11012 6010 11036 6012
rect 11092 6010 11116 6012
rect 11172 6010 11196 6012
rect 11034 5958 11036 6010
rect 11098 5958 11110 6010
rect 11172 5958 11174 6010
rect 11012 5956 11036 5958
rect 11092 5956 11116 5958
rect 11172 5956 11196 5958
rect 10956 5936 11252 5956
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10980 5681 11008 5714
rect 11532 5710 11560 6870
rect 11794 6760 11850 6769
rect 11794 6695 11850 6704
rect 11520 5704 11572 5710
rect 10966 5672 11022 5681
rect 11520 5646 11572 5652
rect 10966 5607 11022 5616
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10980 5302 11008 5607
rect 10968 5296 11020 5302
rect 10968 5238 11020 5244
rect 11532 5234 11560 5646
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 10956 4924 11252 4944
rect 11012 4922 11036 4924
rect 11092 4922 11116 4924
rect 11172 4922 11196 4924
rect 11034 4870 11036 4922
rect 11098 4870 11110 4922
rect 11172 4870 11174 4922
rect 11012 4868 11036 4870
rect 11092 4868 11116 4870
rect 11172 4868 11196 4870
rect 10956 4848 11252 4868
rect 11348 4826 11376 4966
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11532 4758 11560 5170
rect 11808 4826 11836 6695
rect 12072 5092 12124 5098
rect 12072 5034 12124 5040
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11900 4826 11928 4966
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11520 4752 11572 4758
rect 11520 4694 11572 4700
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11532 4282 11560 4558
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 11808 4214 11836 4762
rect 12084 4622 12112 5034
rect 12176 4729 12204 7103
rect 12346 6896 12402 6905
rect 12346 6831 12402 6840
rect 12360 5914 12388 6831
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12360 5370 12388 5850
rect 12452 5778 12480 7482
rect 12636 6610 12664 16102
rect 12714 16079 12770 16088
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 13004 15162 13032 15846
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12820 13802 12848 14350
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 13004 13326 13032 13874
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12728 11218 12756 12038
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12728 10810 12756 11154
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12820 6798 12848 7686
rect 13084 7472 13136 7478
rect 13084 7414 13136 7420
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 7002 12940 7142
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12544 6582 12664 6610
rect 12544 5846 12572 6582
rect 12820 6322 12848 6734
rect 12912 6458 12940 6938
rect 13096 6866 13124 7414
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13096 6458 13124 6802
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12714 6216 12770 6225
rect 12714 6151 12770 6160
rect 12728 5914 12756 6151
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12544 5370 12572 5782
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12162 4720 12218 4729
rect 12162 4655 12218 4664
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12084 4282 12112 4558
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 11796 4208 11848 4214
rect 10046 4176 10102 4185
rect 11796 4150 11848 4156
rect 10046 4111 10102 4120
rect 10956 3836 11252 3856
rect 11012 3834 11036 3836
rect 11092 3834 11116 3836
rect 11172 3834 11196 3836
rect 11034 3782 11036 3834
rect 11098 3782 11110 3834
rect 11172 3782 11174 3834
rect 11012 3780 11036 3782
rect 11092 3780 11116 3782
rect 11172 3780 11196 3782
rect 10956 3760 11252 3780
rect 12084 3738 12112 4218
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10796 3126 10824 3470
rect 11072 3194 11100 3538
rect 12544 3505 12572 5306
rect 12530 3496 12586 3505
rect 12530 3431 12586 3440
rect 13188 3194 13216 19654
rect 13464 18426 13492 20198
rect 15120 20182 15240 20198
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 15108 19848 15160 19854
rect 15212 19802 15240 20182
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 15160 19796 15240 19802
rect 15108 19790 15240 19796
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 13728 19780 13780 19786
rect 13728 19722 13780 19728
rect 13740 19514 13768 19722
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 13740 18970 13768 19450
rect 14016 19446 14044 19790
rect 15120 19774 15240 19790
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 14004 19440 14056 19446
rect 14004 19382 14056 19388
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 13636 18828 13688 18834
rect 13636 18770 13688 18776
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13556 17202 13584 18226
rect 13648 18154 13676 18770
rect 13832 18358 13860 18770
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13832 18170 13860 18294
rect 13636 18148 13688 18154
rect 13636 18090 13688 18096
rect 13740 18142 13860 18170
rect 13648 17610 13676 18090
rect 13740 17882 13768 18142
rect 13820 18080 13872 18086
rect 13924 18068 13952 19314
rect 15120 19310 15148 19654
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 15212 19258 15240 19774
rect 14740 19236 14792 19242
rect 14740 19178 14792 19184
rect 14280 19168 14332 19174
rect 14200 19116 14280 19122
rect 14200 19110 14332 19116
rect 14200 19094 14320 19110
rect 14200 18766 14228 19094
rect 14554 18864 14610 18873
rect 14554 18799 14610 18808
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14200 18426 14228 18702
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14568 18329 14596 18799
rect 14752 18329 14780 19178
rect 14554 18320 14610 18329
rect 14554 18255 14610 18264
rect 14738 18320 14794 18329
rect 14738 18255 14740 18264
rect 14792 18255 14794 18264
rect 14740 18226 14792 18232
rect 13872 18040 13952 18068
rect 13820 18022 13872 18028
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13636 17604 13688 17610
rect 13636 17546 13688 17552
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13832 16674 13860 18022
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 14016 17338 14044 17682
rect 14752 17678 14780 18226
rect 15120 17814 15148 19246
rect 15212 19230 15424 19258
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15108 17808 15160 17814
rect 15108 17750 15160 17756
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14830 17640 14886 17649
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 14108 17270 14136 17614
rect 14830 17575 14886 17584
rect 14096 17264 14148 17270
rect 14096 17206 14148 17212
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 13924 16998 13952 17138
rect 14844 17134 14872 17575
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13924 16794 13952 16934
rect 14844 16833 14872 17070
rect 14924 16992 14976 16998
rect 14924 16934 14976 16940
rect 14830 16824 14886 16833
rect 13912 16788 13964 16794
rect 14830 16759 14832 16768
rect 13912 16730 13964 16736
rect 14884 16759 14886 16768
rect 14832 16730 14884 16736
rect 14844 16699 14872 16730
rect 13832 16646 13952 16674
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13648 13530 13676 13738
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13634 13424 13690 13433
rect 13634 13359 13636 13368
rect 13688 13359 13690 13368
rect 13636 13330 13688 13336
rect 13648 12986 13676 13330
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13740 12442 13768 13262
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13634 11792 13690 11801
rect 13634 11727 13636 11736
rect 13688 11727 13690 11736
rect 13636 11698 13688 11704
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13280 9926 13308 10406
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13280 9518 13308 9862
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13556 9450 13584 10950
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 13556 9110 13584 9386
rect 13648 9178 13676 10134
rect 13832 10130 13860 10678
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13280 7002 13308 7346
rect 13450 7304 13506 7313
rect 13450 7239 13452 7248
rect 13504 7239 13506 7248
rect 13452 7210 13504 7216
rect 13360 7200 13412 7206
rect 13358 7168 13360 7177
rect 13412 7168 13414 7177
rect 13358 7103 13414 7112
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13280 5234 13308 5714
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13450 5128 13506 5137
rect 13648 5098 13676 5510
rect 13450 5063 13506 5072
rect 13636 5092 13688 5098
rect 13464 4826 13492 5063
rect 13636 5034 13688 5040
rect 13542 4992 13598 5001
rect 13542 4927 13598 4936
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13464 4282 13492 4762
rect 13556 4690 13584 4927
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13556 4214 13584 4626
rect 13648 4622 13676 5034
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13648 4282 13676 4558
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 10784 3120 10836 3126
rect 9862 3088 9918 3097
rect 10784 3062 10836 3068
rect 9862 3023 9918 3032
rect 13188 2990 13216 3130
rect 13176 2984 13228 2990
rect 13176 2926 13228 2932
rect 12072 2916 12124 2922
rect 12072 2858 12124 2864
rect 10956 2748 11252 2768
rect 11012 2746 11036 2748
rect 11092 2746 11116 2748
rect 11172 2746 11196 2748
rect 11034 2694 11036 2746
rect 11098 2694 11110 2746
rect 11172 2694 11174 2746
rect 11012 2692 11036 2694
rect 11092 2692 11116 2694
rect 11172 2692 11196 2694
rect 10956 2672 11252 2692
rect 9770 2544 9826 2553
rect 9680 2508 9732 2514
rect 9770 2479 9826 2488
rect 11058 2544 11114 2553
rect 11058 2479 11060 2488
rect 9680 2450 9732 2456
rect 11112 2479 11114 2488
rect 11060 2450 11112 2456
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 9968 1465 9996 2382
rect 9954 1456 10010 1465
rect 9954 1391 10010 1400
rect 10612 480 10640 2382
rect 12084 480 12112 2858
rect 13740 2650 13768 9862
rect 13832 9722 13860 10066
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13924 8673 13952 16646
rect 14936 16017 14964 16934
rect 15304 16794 15332 18022
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 14922 16008 14978 16017
rect 14922 15943 14978 15952
rect 14936 15473 14964 15943
rect 15396 15570 15424 19230
rect 15856 18970 15884 19790
rect 15956 19612 16252 19632
rect 16012 19610 16036 19612
rect 16092 19610 16116 19612
rect 16172 19610 16196 19612
rect 16034 19558 16036 19610
rect 16098 19558 16110 19610
rect 16172 19558 16174 19610
rect 16012 19556 16036 19558
rect 16092 19556 16116 19558
rect 16172 19556 16196 19558
rect 15956 19536 16252 19556
rect 16316 19174 16344 19790
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 16408 18902 16436 19858
rect 16684 19825 16712 20334
rect 17052 20058 17080 20878
rect 18340 20466 18368 23520
rect 20956 21244 21252 21264
rect 21012 21242 21036 21244
rect 21092 21242 21116 21244
rect 21172 21242 21196 21244
rect 21034 21190 21036 21242
rect 21098 21190 21110 21242
rect 21172 21190 21174 21242
rect 21012 21188 21036 21190
rect 21092 21188 21116 21190
rect 21172 21188 21196 21190
rect 20956 21168 21252 21188
rect 21652 20602 21680 23520
rect 24858 23080 24914 23089
rect 24858 23015 24914 23024
rect 24872 22166 24900 23015
rect 21824 22160 21876 22166
rect 21824 22102 21876 22108
rect 24860 22160 24912 22166
rect 24860 22102 24912 22108
rect 21640 20596 21692 20602
rect 21640 20538 21692 20544
rect 20628 20528 20680 20534
rect 20626 20496 20628 20505
rect 20680 20496 20682 20505
rect 18328 20460 18380 20466
rect 20626 20431 20682 20440
rect 18328 20402 18380 20408
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 19260 20058 19288 20334
rect 20720 20324 20772 20330
rect 20720 20266 20772 20272
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 17316 19984 17368 19990
rect 17316 19926 17368 19932
rect 16670 19816 16726 19825
rect 16670 19751 16726 19760
rect 17132 19440 17184 19446
rect 17132 19382 17184 19388
rect 16396 18896 16448 18902
rect 16396 18838 16448 18844
rect 17040 18828 17092 18834
rect 17040 18770 17092 18776
rect 16580 18692 16632 18698
rect 16580 18634 16632 18640
rect 15956 18524 16252 18544
rect 16012 18522 16036 18524
rect 16092 18522 16116 18524
rect 16172 18522 16196 18524
rect 16034 18470 16036 18522
rect 16098 18470 16110 18522
rect 16172 18470 16174 18522
rect 16012 18468 16036 18470
rect 16092 18468 16116 18470
rect 16172 18468 16196 18470
rect 15956 18448 16252 18468
rect 16592 18426 16620 18634
rect 17052 18465 17080 18770
rect 17144 18766 17172 19382
rect 17328 19174 17356 19926
rect 17696 19514 17724 19994
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17684 19508 17736 19514
rect 17684 19450 17736 19456
rect 17880 19446 17908 19790
rect 17868 19440 17920 19446
rect 17868 19382 17920 19388
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17328 18873 17356 19110
rect 19260 18902 19288 19994
rect 20732 19310 20760 20266
rect 20956 20156 21252 20176
rect 21012 20154 21036 20156
rect 21092 20154 21116 20156
rect 21172 20154 21196 20156
rect 21034 20102 21036 20154
rect 21098 20102 21110 20154
rect 21172 20102 21174 20154
rect 21012 20100 21036 20102
rect 21092 20100 21116 20102
rect 21172 20100 21196 20102
rect 20956 20080 21252 20100
rect 21548 19984 21600 19990
rect 21548 19926 21600 19932
rect 21638 19952 21694 19961
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 19248 18896 19300 18902
rect 17314 18864 17370 18873
rect 19248 18838 19300 18844
rect 17314 18799 17370 18808
rect 17868 18828 17920 18834
rect 17868 18770 17920 18776
rect 18420 18828 18472 18834
rect 18420 18770 18472 18776
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17038 18456 17094 18465
rect 16580 18420 16632 18426
rect 17144 18426 17172 18702
rect 17880 18426 17908 18770
rect 17038 18391 17040 18400
rect 16580 18362 16632 18368
rect 17092 18391 17094 18400
rect 17132 18420 17184 18426
rect 17040 18362 17092 18368
rect 17132 18362 17184 18368
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 17144 18329 17172 18362
rect 17130 18320 17186 18329
rect 17130 18255 17186 18264
rect 17144 17882 17172 18255
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 17880 17814 17908 18362
rect 18432 18086 18460 18770
rect 19338 18728 19394 18737
rect 19338 18663 19394 18672
rect 19352 18426 19380 18663
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 18420 18080 18472 18086
rect 18420 18022 18472 18028
rect 16304 17808 16356 17814
rect 17868 17808 17920 17814
rect 16304 17750 16356 17756
rect 17774 17776 17830 17785
rect 15752 17536 15804 17542
rect 15750 17504 15752 17513
rect 15804 17504 15806 17513
rect 15750 17439 15806 17448
rect 15956 17436 16252 17456
rect 16012 17434 16036 17436
rect 16092 17434 16116 17436
rect 16172 17434 16196 17436
rect 16034 17382 16036 17434
rect 16098 17382 16110 17434
rect 16172 17382 16174 17434
rect 16012 17380 16036 17382
rect 16092 17380 16116 17382
rect 16172 17380 16196 17382
rect 15956 17360 16252 17380
rect 15750 17232 15806 17241
rect 15750 17167 15806 17176
rect 15844 17196 15896 17202
rect 15658 17096 15714 17105
rect 15658 17031 15714 17040
rect 15672 16726 15700 17031
rect 15764 16794 15792 17167
rect 15844 17138 15896 17144
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15660 16720 15712 16726
rect 15660 16662 15712 16668
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 14922 15464 14978 15473
rect 14922 15399 14978 15408
rect 15304 14482 15332 15506
rect 15396 15162 15424 15506
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14292 13870 14320 14214
rect 15304 14006 15332 14418
rect 15396 14074 15424 14486
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15016 14000 15068 14006
rect 14922 13968 14978 13977
rect 15016 13942 15068 13948
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 14922 13903 14924 13912
rect 14976 13903 14978 13912
rect 14924 13874 14976 13880
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14660 13530 14688 13738
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 14016 12889 14044 13330
rect 14280 12912 14332 12918
rect 14002 12880 14058 12889
rect 14280 12854 14332 12860
rect 14002 12815 14058 12824
rect 14016 12782 14044 12815
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14292 11694 14320 12854
rect 14936 12850 14964 13874
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14648 12640 14700 12646
rect 14646 12608 14648 12617
rect 14740 12640 14792 12646
rect 14700 12608 14702 12617
rect 14740 12582 14792 12588
rect 14646 12543 14702 12552
rect 14752 12170 14780 12582
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14936 12102 14964 12786
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14924 11824 14976 11830
rect 14924 11766 14976 11772
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14464 11008 14516 11014
rect 14464 10950 14516 10956
rect 14200 10810 14228 10950
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14476 10606 14504 10950
rect 14936 10810 14964 11766
rect 15028 11762 15056 13942
rect 15396 13462 15424 14010
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15212 13161 15240 13262
rect 15198 13152 15254 13161
rect 15198 13087 15254 13096
rect 15212 12646 15240 13087
rect 15488 13002 15516 16186
rect 15672 16182 15700 16662
rect 15764 16250 15792 16730
rect 15856 16590 15884 17138
rect 16316 16794 16344 17750
rect 16488 17740 16540 17746
rect 17868 17750 17920 17756
rect 17774 17711 17830 17720
rect 16488 17682 16540 17688
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16408 17134 16436 17478
rect 16500 17202 16528 17682
rect 17788 17338 17816 17711
rect 18234 17640 18290 17649
rect 18234 17575 18236 17584
rect 18288 17575 18290 17584
rect 18236 17546 18288 17552
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 17788 17134 17816 17274
rect 18248 17202 18276 17546
rect 18432 17270 18460 18022
rect 19720 17678 19748 18566
rect 20720 18352 20772 18358
rect 20720 18294 20772 18300
rect 20168 18216 20220 18222
rect 20168 18158 20220 18164
rect 19800 18080 19852 18086
rect 19800 18022 19852 18028
rect 19812 17882 19840 18022
rect 19800 17876 19852 17882
rect 19800 17818 19852 17824
rect 19708 17672 19760 17678
rect 19708 17614 19760 17620
rect 19248 17536 19300 17542
rect 19248 17478 19300 17484
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 18510 17232 18566 17241
rect 18236 17196 18288 17202
rect 18510 17167 18566 17176
rect 18880 17196 18932 17202
rect 18236 17138 18288 17144
rect 18524 17134 18552 17167
rect 18880 17138 18932 17144
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15856 16250 15884 16526
rect 15956 16348 16252 16368
rect 16012 16346 16036 16348
rect 16092 16346 16116 16348
rect 16172 16346 16196 16348
rect 16034 16294 16036 16346
rect 16098 16294 16110 16346
rect 16172 16294 16174 16346
rect 16012 16292 16036 16294
rect 16092 16292 16116 16294
rect 16172 16292 16196 16294
rect 15956 16272 16252 16292
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15660 16176 15712 16182
rect 15660 16118 15712 16124
rect 15672 15450 15700 16118
rect 16316 15706 16344 16730
rect 16304 15700 16356 15706
rect 16304 15642 16356 15648
rect 15672 15422 15792 15450
rect 15396 12974 15516 13002
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15106 12336 15162 12345
rect 15396 12322 15424 12974
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15488 12481 15516 12582
rect 15474 12472 15530 12481
rect 15474 12407 15530 12416
rect 15396 12294 15608 12322
rect 15106 12271 15162 12280
rect 15120 11898 15148 12271
rect 15474 12200 15530 12209
rect 15474 12135 15530 12144
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 14936 10674 14964 10746
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14740 10532 14792 10538
rect 14740 10474 14792 10480
rect 14752 10266 14780 10474
rect 15212 10282 15240 11494
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15304 10810 15332 11086
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15304 10606 15332 10746
rect 15396 10674 15424 12038
rect 15488 11257 15516 12135
rect 15474 11248 15530 11257
rect 15474 11183 15530 11192
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15382 10568 15438 10577
rect 15580 10554 15608 12294
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15672 12209 15700 12242
rect 15658 12200 15714 12209
rect 15658 12135 15714 12144
rect 15672 11218 15700 12135
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15672 10713 15700 11154
rect 15658 10704 15714 10713
rect 15658 10639 15714 10648
rect 15382 10503 15438 10512
rect 15488 10526 15608 10554
rect 15396 10305 15424 10503
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 15120 10254 15240 10282
rect 15382 10296 15438 10305
rect 15120 10198 15148 10254
rect 15382 10231 15438 10240
rect 15108 10192 15160 10198
rect 15108 10134 15160 10140
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 14016 9382 14044 9998
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 13910 8664 13966 8673
rect 14476 8634 14504 9318
rect 14646 8936 14702 8945
rect 14646 8871 14702 8880
rect 14660 8838 14688 8871
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 13910 8599 13966 8608
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14660 8430 14688 8774
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14370 7576 14426 7585
rect 14370 7511 14426 7520
rect 14384 7274 14412 7511
rect 14660 7410 14688 7686
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14372 7268 14424 7274
rect 14372 7210 14424 7216
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14568 7002 14596 7142
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14660 5370 14688 7346
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 14924 7200 14976 7206
rect 14922 7168 14924 7177
rect 14976 7168 14978 7177
rect 14922 7103 14978 7112
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 15198 5264 15254 5273
rect 15198 5199 15254 5208
rect 15212 5166 15240 5199
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15396 4758 15424 7210
rect 15488 5681 15516 10526
rect 15658 10432 15714 10441
rect 15658 10367 15714 10376
rect 15672 10169 15700 10367
rect 15658 10160 15714 10169
rect 15658 10095 15660 10104
rect 15712 10095 15714 10104
rect 15660 10066 15712 10072
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15580 9382 15608 9998
rect 15672 9722 15700 10066
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15580 8537 15608 9318
rect 15658 8936 15714 8945
rect 15658 8871 15714 8880
rect 15566 8528 15622 8537
rect 15566 8463 15622 8472
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15580 7206 15608 7890
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15474 5672 15530 5681
rect 15474 5607 15530 5616
rect 15580 5137 15608 7142
rect 15672 5778 15700 8871
rect 15764 7342 15792 15422
rect 15956 15260 16252 15280
rect 16012 15258 16036 15260
rect 16092 15258 16116 15260
rect 16172 15258 16196 15260
rect 16034 15206 16036 15258
rect 16098 15206 16110 15258
rect 16172 15206 16174 15258
rect 16012 15204 16036 15206
rect 16092 15204 16116 15206
rect 16172 15204 16196 15206
rect 15956 15184 16252 15204
rect 16316 15162 16344 15642
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 16684 14550 16712 15302
rect 16672 14544 16724 14550
rect 16672 14486 16724 14492
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 15956 14172 16252 14192
rect 16012 14170 16036 14172
rect 16092 14170 16116 14172
rect 16172 14170 16196 14172
rect 16034 14118 16036 14170
rect 16098 14118 16110 14170
rect 16172 14118 16174 14170
rect 16012 14116 16036 14118
rect 16092 14116 16116 14118
rect 16172 14116 16196 14118
rect 15956 14096 16252 14116
rect 16684 13977 16712 14214
rect 16776 14074 16804 17070
rect 18604 17060 18656 17066
rect 18604 17002 18656 17008
rect 17960 16992 18012 16998
rect 17880 16940 17960 16946
rect 17880 16934 18012 16940
rect 17880 16918 18000 16934
rect 17880 16250 17908 16918
rect 17972 16794 18000 16918
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 18616 16697 18644 17002
rect 18602 16688 18658 16697
rect 18602 16623 18658 16632
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 17972 15162 18000 15506
rect 18432 15473 18460 15506
rect 18512 15496 18564 15502
rect 18418 15464 18474 15473
rect 18052 15428 18104 15434
rect 18512 15438 18564 15444
rect 18418 15399 18474 15408
rect 18052 15370 18104 15376
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17972 14657 18000 15098
rect 18064 15094 18092 15370
rect 18432 15162 18460 15399
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18052 15088 18104 15094
rect 18052 15030 18104 15036
rect 17958 14648 18014 14657
rect 18524 14618 18552 15438
rect 17958 14583 18014 14592
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17788 14074 17816 14418
rect 18512 14408 18564 14414
rect 18616 14396 18644 16623
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18708 16250 18736 16526
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18708 15706 18736 16186
rect 18800 16182 18828 16526
rect 18788 16176 18840 16182
rect 18788 16118 18840 16124
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18892 15434 18920 17138
rect 19260 16794 19288 17478
rect 19720 17202 19748 17614
rect 19812 17338 19840 17818
rect 20076 17808 20128 17814
rect 20180 17785 20208 18158
rect 20732 17898 20760 18294
rect 20640 17870 20760 17898
rect 20640 17814 20668 17870
rect 20628 17808 20680 17814
rect 20076 17750 20128 17756
rect 20166 17776 20222 17785
rect 20088 17338 20116 17750
rect 20628 17750 20680 17756
rect 20166 17711 20222 17720
rect 19800 17332 19852 17338
rect 19800 17274 19852 17280
rect 20076 17332 20128 17338
rect 20076 17274 20128 17280
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19260 16640 19288 16730
rect 19720 16658 19748 17138
rect 20824 16810 20852 19450
rect 21560 19174 21588 19926
rect 21638 19887 21640 19896
rect 21692 19887 21694 19896
rect 21640 19858 21692 19864
rect 21652 19514 21680 19858
rect 21640 19508 21692 19514
rect 21640 19450 21692 19456
rect 21548 19168 21600 19174
rect 21548 19110 21600 19116
rect 20956 19068 21252 19088
rect 21012 19066 21036 19068
rect 21092 19066 21116 19068
rect 21172 19066 21196 19068
rect 21034 19014 21036 19066
rect 21098 19014 21110 19066
rect 21172 19014 21174 19066
rect 21012 19012 21036 19014
rect 21092 19012 21116 19014
rect 21172 19012 21196 19014
rect 20956 18992 21252 19012
rect 21178 18864 21234 18873
rect 21178 18799 21234 18808
rect 21192 18426 21220 18799
rect 21364 18760 21416 18766
rect 21364 18702 21416 18708
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 21192 18154 21220 18362
rect 21284 18290 21312 18566
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21376 18222 21404 18702
rect 21560 18426 21588 19110
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 21364 18216 21416 18222
rect 21364 18158 21416 18164
rect 21180 18148 21232 18154
rect 21180 18090 21232 18096
rect 20956 17980 21252 18000
rect 21012 17978 21036 17980
rect 21092 17978 21116 17980
rect 21172 17978 21196 17980
rect 21034 17926 21036 17978
rect 21098 17926 21110 17978
rect 21172 17926 21174 17978
rect 21012 17924 21036 17926
rect 21092 17924 21116 17926
rect 21172 17924 21196 17926
rect 20956 17904 21252 17924
rect 21376 17882 21404 18158
rect 21836 18154 21864 22102
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 23676 20398 23704 20742
rect 23664 20392 23716 20398
rect 23664 20334 23716 20340
rect 23676 19961 23704 20334
rect 24676 20324 24728 20330
rect 24676 20266 24728 20272
rect 23662 19952 23718 19961
rect 23662 19887 23718 19896
rect 22928 19712 22980 19718
rect 22928 19654 22980 19660
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 22940 19378 22968 19654
rect 23480 19508 23532 19514
rect 23480 19450 23532 19456
rect 22928 19372 22980 19378
rect 22928 19314 22980 19320
rect 22468 19304 22520 19310
rect 22468 19246 22520 19252
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 21824 18148 21876 18154
rect 21824 18090 21876 18096
rect 21364 17876 21416 17882
rect 21364 17818 21416 17824
rect 20956 16892 21252 16912
rect 21012 16890 21036 16892
rect 21092 16890 21116 16892
rect 21172 16890 21196 16892
rect 21034 16838 21036 16890
rect 21098 16838 21110 16890
rect 21172 16838 21174 16890
rect 21012 16836 21036 16838
rect 21092 16836 21116 16838
rect 21172 16836 21196 16838
rect 20956 16816 21252 16836
rect 20732 16782 20852 16810
rect 19229 16612 19288 16640
rect 19708 16652 19760 16658
rect 19229 16538 19257 16612
rect 19708 16594 19760 16600
rect 20732 16590 20760 16782
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 20720 16584 20772 16590
rect 19229 16510 19288 16538
rect 20720 16526 20772 16532
rect 19156 16448 19208 16454
rect 19260 16436 19288 16510
rect 19260 16408 19380 16436
rect 19156 16390 19208 16396
rect 19168 16114 19196 16390
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 18880 15428 18932 15434
rect 18880 15370 18932 15376
rect 18972 14952 19024 14958
rect 18694 14920 18750 14929
rect 18972 14894 19024 14900
rect 18694 14855 18750 14864
rect 18708 14482 18736 14855
rect 18880 14816 18932 14822
rect 18880 14758 18932 14764
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18892 14414 18920 14758
rect 18984 14550 19012 14894
rect 18972 14544 19024 14550
rect 18972 14486 19024 14492
rect 18564 14368 18644 14396
rect 18880 14408 18932 14414
rect 18512 14350 18564 14356
rect 18880 14350 18932 14356
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 16670 13968 16726 13977
rect 16670 13903 16726 13912
rect 16854 13968 16910 13977
rect 16854 13903 16910 13912
rect 18236 13932 18288 13938
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 15844 13456 15896 13462
rect 15844 13398 15896 13404
rect 15856 12986 15884 13398
rect 16316 13297 16344 13466
rect 16868 13433 16896 13903
rect 18236 13874 18288 13880
rect 17868 13796 17920 13802
rect 17868 13738 17920 13744
rect 16854 13424 16910 13433
rect 16854 13359 16910 13368
rect 16302 13288 16358 13297
rect 16302 13223 16358 13232
rect 15956 13084 16252 13104
rect 16012 13082 16036 13084
rect 16092 13082 16116 13084
rect 16172 13082 16196 13084
rect 16034 13030 16036 13082
rect 16098 13030 16110 13082
rect 16172 13030 16174 13082
rect 16012 13028 16036 13030
rect 16092 13028 16116 13030
rect 16172 13028 16196 13030
rect 15956 13008 16252 13028
rect 15844 12980 15896 12986
rect 15896 12940 15976 12968
rect 15844 12922 15896 12928
rect 15948 12238 15976 12940
rect 16316 12918 16344 13223
rect 17880 12986 17908 13738
rect 18248 13462 18276 13874
rect 17960 13456 18012 13462
rect 17960 13398 18012 13404
rect 18236 13456 18288 13462
rect 18236 13398 18288 13404
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16764 12708 16816 12714
rect 16764 12650 16816 12656
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 15856 11082 15884 12174
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 15956 11996 16252 12016
rect 16012 11994 16036 11996
rect 16092 11994 16116 11996
rect 16172 11994 16196 11996
rect 16034 11942 16036 11994
rect 16098 11942 16110 11994
rect 16172 11942 16174 11994
rect 16012 11940 16036 11942
rect 16092 11940 16116 11942
rect 16172 11940 16196 11942
rect 15956 11920 16252 11940
rect 16316 11762 16344 12038
rect 16684 11898 16712 12174
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16132 11354 16160 11698
rect 16776 11354 16804 12650
rect 17972 12594 18000 13398
rect 18524 13190 18552 14350
rect 18892 14074 18920 14350
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18694 13968 18750 13977
rect 18694 13903 18750 13912
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 17880 12566 18000 12594
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18142 12608 18198 12617
rect 17880 12306 17908 12566
rect 17960 12368 18012 12374
rect 17960 12310 18012 12316
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 17224 11280 17276 11286
rect 16394 11248 16450 11257
rect 17224 11222 17276 11228
rect 16394 11183 16450 11192
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15856 10305 15884 11018
rect 15956 10908 16252 10928
rect 16012 10906 16036 10908
rect 16092 10906 16116 10908
rect 16172 10906 16196 10908
rect 16034 10854 16036 10906
rect 16098 10854 16110 10906
rect 16172 10854 16174 10906
rect 16012 10852 16036 10854
rect 16092 10852 16116 10854
rect 16172 10852 16196 10854
rect 15956 10832 16252 10852
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 15842 10296 15898 10305
rect 16316 10266 16344 10610
rect 16408 10538 16436 11183
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16486 10840 16542 10849
rect 16486 10775 16542 10784
rect 16396 10532 16448 10538
rect 16396 10474 16448 10480
rect 15842 10231 15898 10240
rect 16304 10260 16356 10266
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15856 6361 15884 10231
rect 16304 10202 16356 10208
rect 16316 10062 16344 10202
rect 16500 10130 16528 10775
rect 16868 10266 16896 11018
rect 17236 10266 17264 11222
rect 17420 11150 17448 11766
rect 17880 11354 17908 12242
rect 17972 11830 18000 12310
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17420 10810 17448 11086
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17868 10804 17920 10810
rect 17972 10792 18000 11154
rect 17920 10764 18000 10792
rect 17868 10746 17920 10752
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 15956 9820 16252 9840
rect 16012 9818 16036 9820
rect 16092 9818 16116 9820
rect 16172 9818 16196 9820
rect 16034 9766 16036 9818
rect 16098 9766 16110 9818
rect 16172 9766 16174 9818
rect 16012 9764 16036 9766
rect 16092 9764 16116 9766
rect 16172 9764 16196 9766
rect 15956 9744 16252 9764
rect 16316 9722 16344 9998
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16764 8968 16816 8974
rect 16762 8936 16764 8945
rect 16816 8936 16818 8945
rect 16762 8871 16818 8880
rect 15956 8732 16252 8752
rect 16012 8730 16036 8732
rect 16092 8730 16116 8732
rect 16172 8730 16196 8732
rect 16034 8678 16036 8730
rect 16098 8678 16110 8730
rect 16172 8678 16174 8730
rect 16012 8676 16036 8678
rect 16092 8676 16116 8678
rect 16172 8676 16196 8678
rect 15956 8656 16252 8676
rect 16776 8566 16804 8871
rect 16868 8634 16896 8978
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 15956 7644 16252 7664
rect 16012 7642 16036 7644
rect 16092 7642 16116 7644
rect 16172 7642 16196 7644
rect 16034 7590 16036 7642
rect 16098 7590 16110 7642
rect 16172 7590 16174 7642
rect 16012 7588 16036 7590
rect 16092 7588 16116 7590
rect 16172 7588 16196 7590
rect 15956 7568 16252 7588
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16132 6798 16160 7142
rect 16120 6792 16172 6798
rect 16118 6760 16120 6769
rect 16172 6760 16174 6769
rect 16118 6695 16174 6704
rect 15956 6556 16252 6576
rect 16012 6554 16036 6556
rect 16092 6554 16116 6556
rect 16172 6554 16196 6556
rect 16034 6502 16036 6554
rect 16098 6502 16110 6554
rect 16172 6502 16174 6554
rect 16012 6500 16036 6502
rect 16092 6500 16116 6502
rect 16172 6500 16196 6502
rect 15956 6480 16252 6500
rect 15842 6352 15898 6361
rect 16316 6322 16344 7686
rect 16408 7478 16436 7822
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 16592 7342 16620 7822
rect 16670 7440 16726 7449
rect 16868 7410 16896 8570
rect 16670 7375 16726 7384
rect 16856 7404 16908 7410
rect 16580 7336 16632 7342
rect 16500 7296 16580 7324
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 15842 6287 15898 6296
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 15752 6180 15804 6186
rect 15752 6122 15804 6128
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15566 5128 15622 5137
rect 15672 5098 15700 5714
rect 15764 5370 15792 6122
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15566 5063 15622 5072
rect 15660 5092 15712 5098
rect 15660 5034 15712 5040
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 15672 3670 15700 5034
rect 15856 4162 15884 6054
rect 16304 5840 16356 5846
rect 16304 5782 16356 5788
rect 15956 5468 16252 5488
rect 16012 5466 16036 5468
rect 16092 5466 16116 5468
rect 16172 5466 16196 5468
rect 16034 5414 16036 5466
rect 16098 5414 16110 5466
rect 16172 5414 16174 5466
rect 16012 5412 16036 5414
rect 16092 5412 16116 5414
rect 16172 5412 16196 5414
rect 15956 5392 16252 5412
rect 16316 5370 16344 5782
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16212 5092 16264 5098
rect 16212 5034 16264 5040
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16132 4826 16160 4966
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16224 4690 16252 5034
rect 16408 4842 16436 6598
rect 16500 5846 16528 7296
rect 16580 7278 16632 7284
rect 16684 7274 16712 7375
rect 16856 7346 16908 7352
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16868 6866 16896 7346
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17512 6458 17540 6734
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17604 6390 17632 6734
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 17592 6384 17644 6390
rect 17592 6326 17644 6332
rect 17236 5914 17264 6326
rect 17972 6118 18000 6149
rect 17960 6112 18012 6118
rect 17958 6080 17960 6089
rect 18012 6080 18014 6089
rect 17958 6015 18014 6024
rect 17972 5914 18000 6015
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 16488 5840 16540 5846
rect 16488 5782 16540 5788
rect 16486 5536 16542 5545
rect 16486 5471 16542 5480
rect 16500 5166 16528 5471
rect 16670 5400 16726 5409
rect 16670 5335 16726 5344
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16684 5030 16712 5335
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16316 4814 16436 4842
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 15956 4380 16252 4400
rect 16012 4378 16036 4380
rect 16092 4378 16116 4380
rect 16172 4378 16196 4380
rect 16034 4326 16036 4378
rect 16098 4326 16110 4378
rect 16172 4326 16174 4378
rect 16012 4324 16036 4326
rect 16092 4324 16116 4326
rect 16172 4324 16196 4326
rect 15956 4304 16252 4324
rect 15856 4146 15976 4162
rect 15856 4140 15988 4146
rect 15856 4134 15936 4140
rect 15936 4082 15988 4088
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15660 3664 15712 3670
rect 15660 3606 15712 3612
rect 15856 3194 15884 3878
rect 15948 3738 15976 4082
rect 16316 4010 16344 4814
rect 17236 4758 17264 5850
rect 17224 4752 17276 4758
rect 17224 4694 17276 4700
rect 16670 4448 16726 4457
rect 16670 4383 16726 4392
rect 16394 4176 16450 4185
rect 16394 4111 16450 4120
rect 16488 4140 16540 4146
rect 16304 4004 16356 4010
rect 16304 3946 16356 3952
rect 15936 3732 15988 3738
rect 15936 3674 15988 3680
rect 15956 3292 16252 3312
rect 16012 3290 16036 3292
rect 16092 3290 16116 3292
rect 16172 3290 16196 3292
rect 16034 3238 16036 3290
rect 16098 3238 16110 3290
rect 16172 3238 16174 3290
rect 16012 3236 16036 3238
rect 16092 3236 16116 3238
rect 16172 3236 16196 3238
rect 15956 3216 16252 3236
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 14924 2916 14976 2922
rect 14924 2858 14976 2864
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 13452 2440 13504 2446
rect 13452 2382 13504 2388
rect 13464 480 13492 2382
rect 14936 480 14964 2858
rect 16408 2650 16436 4111
rect 16488 4082 16540 4088
rect 16500 3670 16528 4082
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 16684 3194 16712 4383
rect 17236 4282 17264 4694
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17604 3670 17632 4422
rect 17592 3664 17644 3670
rect 17592 3606 17644 3612
rect 17604 3194 17632 3606
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17788 3194 17816 3538
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 16684 2990 16712 3130
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 17776 2984 17828 2990
rect 17776 2926 17828 2932
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 15956 2204 16252 2224
rect 16012 2202 16036 2204
rect 16092 2202 16116 2204
rect 16172 2202 16196 2204
rect 16034 2150 16036 2202
rect 16098 2150 16110 2202
rect 16172 2150 16174 2202
rect 16012 2148 16036 2150
rect 16092 2148 16116 2150
rect 16172 2148 16196 2150
rect 15956 2128 16252 2148
rect 16316 480 16344 2382
rect 17788 480 17816 2926
rect 18064 2530 18092 12582
rect 18142 12543 18198 12552
rect 18156 11626 18184 12543
rect 18144 11620 18196 11626
rect 18144 11562 18196 11568
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18432 11286 18460 11494
rect 18420 11280 18472 11286
rect 18420 11222 18472 11228
rect 18420 11076 18472 11082
rect 18420 11018 18472 11024
rect 18432 10266 18460 11018
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18236 10192 18288 10198
rect 18236 10134 18288 10140
rect 18248 9382 18276 10134
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18156 7342 18184 8774
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18156 6798 18184 7278
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18156 6322 18184 6734
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 18248 2582 18276 9318
rect 18524 7449 18552 13126
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18616 12442 18644 12786
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 18708 11336 18736 13903
rect 18892 13530 18920 14010
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 19076 12832 19104 15846
rect 19168 15706 19196 16050
rect 19352 16046 19380 16408
rect 20732 16182 20760 16526
rect 21008 16250 21036 16594
rect 21824 16448 21876 16454
rect 21824 16390 21876 16396
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 20720 16176 20772 16182
rect 20720 16118 20772 16124
rect 21732 16176 21784 16182
rect 21732 16118 21784 16124
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 20956 15804 21252 15824
rect 21012 15802 21036 15804
rect 21092 15802 21116 15804
rect 21172 15802 21196 15804
rect 21034 15750 21036 15802
rect 21098 15750 21110 15802
rect 21172 15750 21174 15802
rect 21012 15748 21036 15750
rect 21092 15748 21116 15750
rect 21172 15748 21196 15750
rect 20956 15728 21252 15748
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 21744 15570 21772 16118
rect 21836 16114 21864 16390
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 21836 15638 21864 16050
rect 21824 15632 21876 15638
rect 21824 15574 21876 15580
rect 21732 15564 21784 15570
rect 21732 15506 21784 15512
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19260 15144 19288 15370
rect 21744 15162 21772 15506
rect 21836 15162 21864 15574
rect 19340 15156 19392 15162
rect 19260 15116 19340 15144
rect 19340 15098 19392 15104
rect 21732 15156 21784 15162
rect 21732 15098 21784 15104
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 19892 14884 19944 14890
rect 19892 14826 19944 14832
rect 19904 14657 19932 14826
rect 20956 14716 21252 14736
rect 21012 14714 21036 14716
rect 21092 14714 21116 14716
rect 21172 14714 21196 14716
rect 21034 14662 21036 14714
rect 21098 14662 21110 14714
rect 21172 14662 21174 14714
rect 21012 14660 21036 14662
rect 21092 14660 21116 14662
rect 21172 14660 21196 14662
rect 19890 14648 19946 14657
rect 20956 14640 21252 14660
rect 19890 14583 19892 14592
rect 19944 14583 19946 14592
rect 19892 14554 19944 14560
rect 20444 14544 20496 14550
rect 20444 14486 20496 14492
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 18984 12804 19104 12832
rect 19168 12832 19196 13194
rect 20456 12850 20484 14486
rect 21744 14482 21772 15098
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 20548 13870 20576 14418
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20732 13977 20760 14010
rect 20718 13968 20774 13977
rect 20718 13903 20774 13912
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20444 12844 20496 12850
rect 19168 12804 19257 12832
rect 18880 11552 18932 11558
rect 18880 11494 18932 11500
rect 18616 11308 18736 11336
rect 18616 10130 18644 11308
rect 18696 11212 18748 11218
rect 18696 11154 18748 11160
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18708 9654 18736 11154
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18800 10538 18828 11086
rect 18892 10810 18920 11494
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18800 10266 18828 10474
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18696 9648 18748 9654
rect 18696 9590 18748 9596
rect 18800 9382 18828 10066
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18510 7440 18566 7449
rect 18510 7375 18566 7384
rect 18418 7304 18474 7313
rect 18418 7239 18474 7248
rect 18432 6254 18460 7239
rect 18696 6724 18748 6730
rect 18696 6666 18748 6672
rect 18708 6610 18736 6666
rect 18616 6582 18736 6610
rect 18510 6488 18566 6497
rect 18510 6423 18566 6432
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18524 6118 18552 6423
rect 18616 6322 18644 6582
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18512 6112 18564 6118
rect 18512 6054 18564 6060
rect 18616 5914 18644 6258
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18616 3058 18644 3334
rect 18800 3233 18828 9318
rect 18984 7290 19012 12804
rect 19229 12753 19257 12804
rect 20444 12786 20496 12792
rect 19229 12744 19302 12753
rect 19229 12702 19246 12744
rect 19246 12679 19302 12688
rect 19156 12640 19208 12646
rect 19154 12608 19156 12617
rect 19208 12608 19210 12617
rect 19154 12543 19210 12552
rect 20456 12442 20484 12786
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 20548 12345 20576 13806
rect 20956 13628 21252 13648
rect 21012 13626 21036 13628
rect 21092 13626 21116 13628
rect 21172 13626 21196 13628
rect 21034 13574 21036 13626
rect 21098 13574 21110 13626
rect 21172 13574 21174 13626
rect 21012 13572 21036 13574
rect 21092 13572 21116 13574
rect 21172 13572 21196 13574
rect 20956 13552 21252 13572
rect 20718 13016 20774 13025
rect 20718 12951 20774 12960
rect 20732 12730 20760 12951
rect 20640 12702 20760 12730
rect 21730 12744 21786 12753
rect 20812 12708 20864 12714
rect 20534 12336 20590 12345
rect 20640 12322 20668 12702
rect 21730 12679 21732 12688
rect 20812 12650 20864 12656
rect 21784 12679 21786 12688
rect 21732 12650 21784 12656
rect 20718 12608 20774 12617
rect 20718 12543 20774 12552
rect 20732 12442 20760 12543
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20640 12294 20760 12322
rect 20534 12271 20590 12280
rect 19156 11756 19208 11762
rect 19156 11698 19208 11704
rect 19064 11620 19116 11626
rect 19064 11562 19116 11568
rect 19076 10713 19104 11562
rect 19168 11150 19196 11698
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 19062 10704 19118 10713
rect 19444 10674 19472 11018
rect 19522 10976 19578 10985
rect 19522 10911 19578 10920
rect 19062 10639 19118 10648
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19156 10464 19208 10470
rect 19156 10406 19208 10412
rect 19062 10296 19118 10305
rect 19062 10231 19064 10240
rect 19116 10231 19118 10240
rect 19064 10202 19116 10208
rect 19168 10033 19196 10406
rect 19444 10062 19472 10610
rect 19536 10538 19564 10911
rect 19524 10532 19576 10538
rect 19524 10474 19576 10480
rect 19432 10056 19484 10062
rect 19154 10024 19210 10033
rect 19432 9998 19484 10004
rect 19154 9959 19210 9968
rect 19154 9616 19210 9625
rect 19444 9586 19472 9998
rect 19154 9551 19210 9560
rect 19432 9580 19484 9586
rect 19168 9382 19196 9551
rect 19432 9522 19484 9528
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19338 9480 19394 9489
rect 19156 9376 19208 9382
rect 19156 9318 19208 9324
rect 19168 9178 19196 9318
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 19260 8838 19288 9454
rect 19338 9415 19394 9424
rect 19352 9110 19380 9415
rect 19340 9104 19392 9110
rect 19340 9046 19392 9052
rect 19248 8832 19300 8838
rect 19246 8800 19248 8809
rect 19300 8800 19302 8809
rect 19246 8735 19302 8744
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19260 8378 19288 8502
rect 19260 8350 19380 8378
rect 19062 7984 19118 7993
rect 19062 7919 19118 7928
rect 18892 7262 19012 7290
rect 18786 3224 18842 3233
rect 18786 3159 18842 3168
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18616 2650 18644 2994
rect 18892 2990 18920 7262
rect 18972 7200 19024 7206
rect 19076 7177 19104 7919
rect 19352 7342 19380 8350
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 18972 7142 19024 7148
rect 19062 7168 19118 7177
rect 18984 7002 19012 7142
rect 19062 7103 19118 7112
rect 18972 6996 19024 7002
rect 18972 6938 19024 6944
rect 19076 6866 19104 7103
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 19076 6458 19104 6802
rect 19352 6458 19380 6938
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19260 5370 19288 5850
rect 19536 5817 19564 10474
rect 20548 10130 20576 12271
rect 20536 10124 20588 10130
rect 20536 10066 20588 10072
rect 20352 9920 20404 9926
rect 20352 9862 20404 9868
rect 19616 9444 19668 9450
rect 19616 9386 19668 9392
rect 19628 9178 19656 9386
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 20364 9042 20392 9862
rect 20548 9722 20576 10066
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20444 9104 20496 9110
rect 20444 9046 20496 9052
rect 20352 9036 20404 9042
rect 20352 8978 20404 8984
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20180 8430 20208 8774
rect 20364 8634 20392 8978
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20180 7750 20208 8366
rect 20168 7744 20220 7750
rect 20168 7686 20220 7692
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 19904 7002 19932 7278
rect 19892 6996 19944 7002
rect 19892 6938 19944 6944
rect 19522 5808 19578 5817
rect 19522 5743 19578 5752
rect 19708 5704 19760 5710
rect 19708 5646 19760 5652
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19248 5364 19300 5370
rect 19248 5306 19300 5312
rect 19352 4826 19380 5510
rect 19444 5030 19472 5578
rect 19720 5370 19748 5646
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 20180 5030 20208 7686
rect 20456 6458 20484 9046
rect 20640 7342 20668 9454
rect 20732 8809 20760 12294
rect 20824 11762 20852 12650
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 20956 12540 21252 12560
rect 21012 12538 21036 12540
rect 21092 12538 21116 12540
rect 21172 12538 21196 12540
rect 21034 12486 21036 12538
rect 21098 12486 21110 12538
rect 21172 12486 21174 12538
rect 21012 12484 21036 12486
rect 21092 12484 21116 12486
rect 21172 12484 21196 12486
rect 20956 12464 21252 12484
rect 21560 12238 21588 12582
rect 21730 12472 21786 12481
rect 21730 12407 21786 12416
rect 21640 12300 21692 12306
rect 21640 12242 21692 12248
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21376 11898 21404 12174
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 21272 11688 21324 11694
rect 21270 11656 21272 11665
rect 21324 11656 21326 11665
rect 21270 11591 21326 11600
rect 20956 11452 21252 11472
rect 21012 11450 21036 11452
rect 21092 11450 21116 11452
rect 21172 11450 21196 11452
rect 21034 11398 21036 11450
rect 21098 11398 21110 11450
rect 21172 11398 21174 11450
rect 21012 11396 21036 11398
rect 21092 11396 21116 11398
rect 21172 11396 21196 11398
rect 20956 11376 21252 11396
rect 21376 11354 21404 11834
rect 21560 11830 21588 12174
rect 21548 11824 21600 11830
rect 21548 11766 21600 11772
rect 21652 11626 21680 12242
rect 21744 11914 21772 12407
rect 21744 11886 21864 11914
rect 21640 11620 21692 11626
rect 21640 11562 21692 11568
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21468 11082 21496 11494
rect 21652 11354 21680 11562
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 21744 11121 21772 11154
rect 21730 11112 21786 11121
rect 21456 11076 21508 11082
rect 21730 11047 21786 11056
rect 21456 11018 21508 11024
rect 21468 10849 21496 11018
rect 21454 10840 21510 10849
rect 21744 10810 21772 11047
rect 21454 10775 21510 10784
rect 21732 10804 21784 10810
rect 21732 10746 21784 10752
rect 20956 10364 21252 10384
rect 21012 10362 21036 10364
rect 21092 10362 21116 10364
rect 21172 10362 21196 10364
rect 21034 10310 21036 10362
rect 21098 10310 21110 10362
rect 21172 10310 21174 10362
rect 21012 10308 21036 10310
rect 21092 10308 21116 10310
rect 21172 10308 21196 10310
rect 20956 10288 21252 10308
rect 21362 10296 21418 10305
rect 21362 10231 21418 10240
rect 21376 10062 21404 10231
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 21364 10056 21416 10062
rect 21364 9998 21416 10004
rect 20824 9382 20852 9998
rect 21468 9382 21496 10066
rect 21546 10024 21602 10033
rect 21546 9959 21602 9968
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 20956 9276 21252 9296
rect 21012 9274 21036 9276
rect 21092 9274 21116 9276
rect 21172 9274 21196 9276
rect 21034 9222 21036 9274
rect 21098 9222 21110 9274
rect 21172 9222 21174 9274
rect 21012 9220 21036 9222
rect 21092 9220 21116 9222
rect 21172 9220 21196 9222
rect 20956 9200 21252 9220
rect 21284 8838 21312 9318
rect 21272 8832 21324 8838
rect 20718 8800 20774 8809
rect 21272 8774 21324 8780
rect 21362 8800 21418 8809
rect 20718 8735 20774 8744
rect 21362 8735 21418 8744
rect 20812 8356 20864 8362
rect 20812 8298 20864 8304
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 20456 6254 20484 6394
rect 20444 6248 20496 6254
rect 20444 6190 20496 6196
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 20548 5914 20576 6054
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20534 5808 20590 5817
rect 20534 5743 20590 5752
rect 20350 5264 20406 5273
rect 20350 5199 20352 5208
rect 20404 5199 20406 5208
rect 20352 5170 20404 5176
rect 20548 5098 20576 5743
rect 20536 5092 20588 5098
rect 20536 5034 20588 5040
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 20168 5024 20220 5030
rect 20168 4966 20220 4972
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19248 4480 19300 4486
rect 19248 4422 19300 4428
rect 19260 4185 19288 4422
rect 19246 4176 19302 4185
rect 19246 4111 19302 4120
rect 19352 3738 19380 4762
rect 19444 4078 19472 4966
rect 19708 4616 19760 4622
rect 19892 4616 19944 4622
rect 19708 4558 19760 4564
rect 19890 4584 19892 4593
rect 19944 4584 19946 4593
rect 19720 4146 19748 4558
rect 19890 4519 19946 4528
rect 19904 4282 19932 4519
rect 19892 4276 19944 4282
rect 19892 4218 19944 4224
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19982 3224 20038 3233
rect 19982 3159 20038 3168
rect 18880 2984 18932 2990
rect 18880 2926 18932 2932
rect 19156 2916 19208 2922
rect 19156 2858 19208 2864
rect 19168 2825 19196 2858
rect 19154 2816 19210 2825
rect 19154 2751 19210 2760
rect 19996 2650 20024 3159
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 17880 2514 18092 2530
rect 18236 2576 18288 2582
rect 18236 2518 18288 2524
rect 17868 2508 18092 2514
rect 17920 2502 18092 2508
rect 17868 2450 17920 2456
rect 20088 2446 20116 2994
rect 20180 2990 20208 4966
rect 20548 4826 20576 5034
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 20732 4457 20760 7686
rect 20824 7546 20852 8298
rect 20956 8188 21252 8208
rect 21012 8186 21036 8188
rect 21092 8186 21116 8188
rect 21172 8186 21196 8188
rect 21034 8134 21036 8186
rect 21098 8134 21110 8186
rect 21172 8134 21174 8186
rect 21012 8132 21036 8134
rect 21092 8132 21116 8134
rect 21172 8132 21196 8134
rect 20956 8112 21252 8132
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20956 7100 21252 7120
rect 21012 7098 21036 7100
rect 21092 7098 21116 7100
rect 21172 7098 21196 7100
rect 21034 7046 21036 7098
rect 21098 7046 21110 7098
rect 21172 7046 21174 7098
rect 21012 7044 21036 7046
rect 21092 7044 21116 7046
rect 21172 7044 21196 7046
rect 20956 7024 21252 7044
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 21100 6322 21128 6598
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 21100 6202 21128 6258
rect 21100 6174 21312 6202
rect 20812 6112 20864 6118
rect 20812 6054 20864 6060
rect 20824 5914 20852 6054
rect 20956 6012 21252 6032
rect 21012 6010 21036 6012
rect 21092 6010 21116 6012
rect 21172 6010 21196 6012
rect 21034 5958 21036 6010
rect 21098 5958 21110 6010
rect 21172 5958 21174 6010
rect 21012 5956 21036 5958
rect 21092 5956 21116 5958
rect 21172 5956 21196 5958
rect 20956 5936 21252 5956
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 21284 5234 21312 6174
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 20956 4924 21252 4944
rect 21012 4922 21036 4924
rect 21092 4922 21116 4924
rect 21172 4922 21196 4924
rect 21034 4870 21036 4922
rect 21098 4870 21110 4922
rect 21172 4870 21174 4922
rect 21012 4868 21036 4870
rect 21092 4868 21116 4870
rect 21172 4868 21196 4870
rect 20956 4848 21252 4868
rect 20718 4448 20774 4457
rect 20718 4383 20774 4392
rect 21284 4282 21312 5170
rect 21376 4486 21404 8735
rect 21468 8634 21496 9318
rect 21456 8628 21508 8634
rect 21456 8570 21508 8576
rect 21560 8242 21588 9959
rect 21836 9625 21864 11886
rect 21822 9616 21878 9625
rect 21468 8214 21588 8242
rect 21744 9574 21822 9602
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21468 4298 21496 8214
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21560 6934 21588 8026
rect 21744 7970 21772 9574
rect 21822 9551 21878 9560
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21836 8634 21864 8978
rect 21928 8838 21956 19110
rect 22480 18902 22508 19246
rect 22652 19168 22704 19174
rect 22652 19110 22704 19116
rect 22664 18970 22692 19110
rect 22652 18964 22704 18970
rect 22652 18906 22704 18912
rect 22468 18896 22520 18902
rect 22468 18838 22520 18844
rect 23020 18828 23072 18834
rect 23020 18770 23072 18776
rect 23032 18358 23060 18770
rect 23492 18766 23520 19450
rect 23768 19378 23796 19654
rect 24688 19446 24716 20266
rect 24676 19440 24728 19446
rect 24676 19382 24728 19388
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 23768 18970 23796 19314
rect 24122 19272 24178 19281
rect 24122 19207 24178 19216
rect 23756 18964 23808 18970
rect 23756 18906 23808 18912
rect 23112 18760 23164 18766
rect 23112 18702 23164 18708
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23020 18352 23072 18358
rect 23020 18294 23072 18300
rect 23032 17882 23060 18294
rect 23124 17882 23152 18702
rect 23492 18426 23520 18702
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 23572 18216 23624 18222
rect 23570 18184 23572 18193
rect 23624 18184 23626 18193
rect 23570 18119 23626 18128
rect 23940 18148 23992 18154
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 23020 17876 23072 17882
rect 23020 17818 23072 17824
rect 23112 17876 23164 17882
rect 23112 17818 23164 17824
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 23124 17338 23152 17614
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 23492 17241 23520 18022
rect 23478 17232 23534 17241
rect 23478 17167 23534 17176
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23110 16144 23166 16153
rect 23110 16079 23166 16088
rect 23124 16046 23152 16079
rect 23112 16040 23164 16046
rect 23112 15982 23164 15988
rect 23112 15360 23164 15366
rect 23112 15302 23164 15308
rect 23124 14550 23152 15302
rect 23492 14929 23520 17070
rect 23478 14920 23534 14929
rect 23478 14855 23534 14864
rect 23112 14544 23164 14550
rect 23112 14486 23164 14492
rect 22560 14476 22612 14482
rect 22560 14418 22612 14424
rect 22572 13977 22600 14418
rect 23124 14074 23152 14486
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 22558 13968 22614 13977
rect 22558 13903 22614 13912
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22112 13190 22140 13670
rect 22572 13530 22600 13903
rect 23480 13728 23532 13734
rect 23480 13670 23532 13676
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 22112 12889 22140 13126
rect 22098 12880 22154 12889
rect 22098 12815 22154 12824
rect 23492 12481 23520 13670
rect 23478 12472 23534 12481
rect 23478 12407 23534 12416
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22006 11792 22062 11801
rect 22006 11727 22062 11736
rect 22284 11756 22336 11762
rect 22020 11558 22048 11727
rect 22284 11698 22336 11704
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22112 10810 22140 11290
rect 22296 11150 22324 11698
rect 22480 11354 22508 12174
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22284 11144 22336 11150
rect 22284 11086 22336 11092
rect 22468 11144 22520 11150
rect 22468 11086 22520 11092
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22480 10470 22508 11086
rect 22468 10464 22520 10470
rect 23480 10464 23532 10470
rect 22468 10406 22520 10412
rect 23400 10412 23480 10418
rect 23400 10406 23532 10412
rect 22480 10266 22508 10406
rect 23400 10390 23520 10406
rect 22468 10260 22520 10266
rect 22468 10202 22520 10208
rect 23296 9988 23348 9994
rect 23296 9930 23348 9936
rect 22558 9616 22614 9625
rect 22192 9580 22244 9586
rect 22558 9551 22560 9560
rect 22192 9522 22244 9528
rect 22612 9551 22614 9560
rect 22560 9522 22612 9528
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21916 8560 21968 8566
rect 21914 8528 21916 8537
rect 21968 8528 21970 8537
rect 21914 8463 21970 8472
rect 22020 8090 22048 9318
rect 22204 9178 22232 9522
rect 22572 9450 22600 9522
rect 23308 9518 23336 9930
rect 23400 9586 23428 10390
rect 23492 10266 23520 10390
rect 23480 10260 23532 10266
rect 23480 10202 23532 10208
rect 23584 10033 23612 18119
rect 23940 18090 23992 18096
rect 23756 17740 23808 17746
rect 23756 17682 23808 17688
rect 23768 17066 23796 17682
rect 23756 17060 23808 17066
rect 23756 17002 23808 17008
rect 23768 16658 23796 17002
rect 23848 16992 23900 16998
rect 23848 16934 23900 16940
rect 23860 16697 23888 16934
rect 23846 16688 23902 16697
rect 23756 16652 23808 16658
rect 23846 16623 23902 16632
rect 23756 16594 23808 16600
rect 23952 16250 23980 18090
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 24044 17921 24072 18022
rect 24030 17912 24086 17921
rect 24030 17847 24086 17856
rect 24032 17740 24084 17746
rect 24032 17682 24084 17688
rect 24044 16998 24072 17682
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 24044 16794 24072 16934
rect 24032 16788 24084 16794
rect 24032 16730 24084 16736
rect 23940 16244 23992 16250
rect 23940 16186 23992 16192
rect 23940 15904 23992 15910
rect 23940 15846 23992 15852
rect 23754 15464 23810 15473
rect 23754 15399 23810 15408
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23676 13462 23704 13670
rect 23664 13456 23716 13462
rect 23664 13398 23716 13404
rect 23676 12986 23704 13398
rect 23664 12980 23716 12986
rect 23664 12922 23716 12928
rect 23570 10024 23626 10033
rect 23570 9959 23626 9968
rect 23584 9586 23612 9959
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23572 9580 23624 9586
rect 23572 9522 23624 9528
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 23296 9512 23348 9518
rect 23296 9454 23348 9460
rect 22560 9444 22612 9450
rect 22560 9386 22612 9392
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 21640 7948 21692 7954
rect 21744 7942 21864 7970
rect 21640 7890 21692 7896
rect 21652 7002 21680 7890
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21744 7546 21772 7822
rect 21732 7540 21784 7546
rect 21732 7482 21784 7488
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 21548 6928 21600 6934
rect 21548 6870 21600 6876
rect 21652 6730 21680 6938
rect 21640 6724 21692 6730
rect 21640 6666 21692 6672
rect 21640 4480 21692 4486
rect 21640 4422 21692 4428
rect 21272 4276 21324 4282
rect 21272 4218 21324 4224
rect 21376 4270 21496 4298
rect 21376 4146 21404 4270
rect 21456 4208 21508 4214
rect 21456 4150 21508 4156
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 20640 4049 20668 4082
rect 20626 4040 20682 4049
rect 20352 4004 20404 4010
rect 20626 3975 20682 3984
rect 20352 3946 20404 3952
rect 20364 3670 20392 3946
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20456 3738 20484 3878
rect 20956 3836 21252 3856
rect 21012 3834 21036 3836
rect 21092 3834 21116 3836
rect 21172 3834 21196 3836
rect 21034 3782 21036 3834
rect 21098 3782 21110 3834
rect 21172 3782 21174 3834
rect 21012 3780 21036 3782
rect 21092 3780 21116 3782
rect 21172 3780 21196 3782
rect 20956 3760 21252 3780
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 20352 3664 20404 3670
rect 20352 3606 20404 3612
rect 20812 3664 20864 3670
rect 20812 3606 20864 3612
rect 20720 3528 20772 3534
rect 20548 3476 20720 3482
rect 20548 3470 20772 3476
rect 20548 3454 20760 3470
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 20180 2650 20208 2926
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 19168 480 19196 2382
rect 20548 2378 20576 3454
rect 20626 2816 20682 2825
rect 20626 2751 20682 2760
rect 20536 2372 20588 2378
rect 20536 2314 20588 2320
rect 20640 480 20668 2751
rect 20824 2650 20852 3606
rect 21468 3534 21496 4150
rect 21652 4146 21680 4422
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 21836 3738 21864 7942
rect 22006 5672 22062 5681
rect 22006 5607 22062 5616
rect 22020 5137 22048 5607
rect 22006 5128 22062 5137
rect 22006 5063 22062 5072
rect 22008 4004 22060 4010
rect 22008 3946 22060 3952
rect 22020 3913 22048 3946
rect 22006 3904 22062 3913
rect 22006 3839 22062 3848
rect 21824 3732 21876 3738
rect 21824 3674 21876 3680
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21376 3194 21404 3470
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 21468 3126 21496 3470
rect 21456 3120 21508 3126
rect 21284 3068 21456 3074
rect 21284 3062 21508 3068
rect 21284 3046 21496 3062
rect 20956 2748 21252 2768
rect 21012 2746 21036 2748
rect 21092 2746 21116 2748
rect 21172 2746 21196 2748
rect 21034 2694 21036 2746
rect 21098 2694 21110 2746
rect 21172 2694 21174 2746
rect 21012 2692 21036 2694
rect 21092 2692 21116 2694
rect 21172 2692 21196 2694
rect 20956 2672 21252 2692
rect 21284 2650 21312 3046
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 22296 2514 22324 8774
rect 22572 6798 22600 9386
rect 22664 9178 22692 9454
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 23296 9036 23348 9042
rect 23296 8978 23348 8984
rect 23204 8832 23256 8838
rect 23204 8774 23256 8780
rect 23216 7002 23244 8774
rect 23308 8566 23336 8978
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23296 8560 23348 8566
rect 23296 8502 23348 8508
rect 23388 8560 23440 8566
rect 23388 8502 23440 8508
rect 23204 6996 23256 7002
rect 23204 6938 23256 6944
rect 22928 6860 22980 6866
rect 22928 6802 22980 6808
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22572 6458 22600 6734
rect 22940 6458 22968 6802
rect 23216 6458 23244 6938
rect 23308 6934 23336 8502
rect 23296 6928 23348 6934
rect 23296 6870 23348 6876
rect 23400 6866 23428 8502
rect 23676 8090 23704 8910
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 23768 6866 23796 15399
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23860 13938 23888 14214
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 23860 13190 23888 13874
rect 23848 13184 23900 13190
rect 23848 13126 23900 13132
rect 23860 12170 23888 13126
rect 23952 12238 23980 15846
rect 24032 13864 24084 13870
rect 24032 13806 24084 13812
rect 24044 13530 24072 13806
rect 24032 13524 24084 13530
rect 24032 13466 24084 13472
rect 23940 12232 23992 12238
rect 23940 12174 23992 12180
rect 23848 12164 23900 12170
rect 23848 12106 23900 12112
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23860 10606 23888 11630
rect 23848 10600 23900 10606
rect 23848 10542 23900 10548
rect 24136 10198 24164 19207
rect 24688 18766 24716 19382
rect 24860 19304 24912 19310
rect 24858 19272 24860 19281
rect 24912 19272 24914 19281
rect 24858 19207 24914 19216
rect 24768 18828 24820 18834
rect 24768 18770 24820 18776
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 24214 18456 24270 18465
rect 24214 18391 24270 18400
rect 24228 15178 24256 18391
rect 24688 18290 24716 18702
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24688 17882 24716 18226
rect 24780 18222 24808 18770
rect 24768 18216 24820 18222
rect 24768 18158 24820 18164
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 24676 17876 24728 17882
rect 24676 17818 24728 17824
rect 24872 17762 24900 18022
rect 24688 17734 24900 17762
rect 24306 17640 24362 17649
rect 24306 17575 24362 17584
rect 24320 16658 24348 17575
rect 24688 17542 24716 17734
rect 24676 17536 24728 17542
rect 24676 17478 24728 17484
rect 24688 17202 24716 17478
rect 24676 17196 24728 17202
rect 24676 17138 24728 17144
rect 24308 16652 24360 16658
rect 24308 16594 24360 16600
rect 24320 15366 24348 16594
rect 24688 16590 24716 17138
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 24676 16584 24728 16590
rect 24676 16526 24728 16532
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24400 16040 24452 16046
rect 24400 15982 24452 15988
rect 24308 15360 24360 15366
rect 24308 15302 24360 15308
rect 24228 15150 24348 15178
rect 24320 12594 24348 15150
rect 24412 14657 24440 15982
rect 24504 15706 24532 16526
rect 24872 16250 24900 16526
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 24872 15706 24900 16186
rect 24492 15700 24544 15706
rect 24492 15642 24544 15648
rect 24860 15700 24912 15706
rect 24860 15642 24912 15648
rect 24504 15473 24532 15642
rect 24490 15464 24546 15473
rect 24490 15399 24546 15408
rect 24768 15360 24820 15366
rect 24768 15302 24820 15308
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24398 14648 24454 14657
rect 24398 14583 24454 14592
rect 24320 12566 24440 12594
rect 24308 12368 24360 12374
rect 24308 12310 24360 12316
rect 24216 12096 24268 12102
rect 24216 12038 24268 12044
rect 24228 11694 24256 12038
rect 24216 11688 24268 11694
rect 24216 11630 24268 11636
rect 24228 10305 24256 11630
rect 24214 10296 24270 10305
rect 24214 10231 24270 10240
rect 24124 10192 24176 10198
rect 24124 10134 24176 10140
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 23940 9648 23992 9654
rect 23940 9590 23992 9596
rect 23848 9444 23900 9450
rect 23848 9386 23900 9392
rect 23388 6860 23440 6866
rect 23388 6802 23440 6808
rect 23756 6860 23808 6866
rect 23756 6802 23808 6808
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22928 6452 22980 6458
rect 22928 6394 22980 6400
rect 23204 6452 23256 6458
rect 23204 6394 23256 6400
rect 22468 5772 22520 5778
rect 22468 5714 22520 5720
rect 22376 5704 22428 5710
rect 22376 5646 22428 5652
rect 22388 5030 22416 5646
rect 22480 5302 22508 5714
rect 23768 5681 23796 6802
rect 23860 6225 23888 9386
rect 23952 7970 23980 9590
rect 24044 9364 24072 9862
rect 24136 9722 24164 10134
rect 24216 10056 24268 10062
rect 24216 9998 24268 10004
rect 24124 9716 24176 9722
rect 24124 9658 24176 9664
rect 24228 9586 24256 9998
rect 24320 9654 24348 12310
rect 24412 9926 24440 12566
rect 24504 12458 24532 14758
rect 24780 13433 24808 15302
rect 24860 14544 24912 14550
rect 24860 14486 24912 14492
rect 24766 13424 24822 13433
rect 24766 13359 24822 13368
rect 24676 13184 24728 13190
rect 24676 13126 24728 13132
rect 24495 12430 24532 12458
rect 24495 12374 24523 12430
rect 24492 12368 24544 12374
rect 24492 12310 24544 12316
rect 24584 12368 24636 12374
rect 24584 12310 24636 12316
rect 24688 12322 24716 13126
rect 24780 12442 24808 13359
rect 24872 12646 24900 14486
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 24964 12442 24992 23520
rect 25134 21312 25190 21321
rect 25134 21247 25190 21256
rect 25044 20256 25096 20262
rect 25044 20198 25096 20204
rect 25056 19378 25084 20198
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 25148 18986 25176 21247
rect 25226 20088 25282 20097
rect 25226 20023 25282 20032
rect 25056 18958 25176 18986
rect 25056 14929 25084 18958
rect 25136 18828 25188 18834
rect 25136 18770 25188 18776
rect 25148 18737 25176 18770
rect 25134 18728 25190 18737
rect 25134 18663 25190 18672
rect 25148 18358 25176 18663
rect 25136 18352 25188 18358
rect 25134 18320 25136 18329
rect 25188 18320 25190 18329
rect 25134 18255 25190 18264
rect 25240 15994 25268 20023
rect 25318 19408 25374 19417
rect 25318 19343 25374 19352
rect 25332 18465 25360 19343
rect 25318 18456 25374 18465
rect 25318 18391 25374 18400
rect 25318 17640 25374 17649
rect 25318 17575 25374 17584
rect 25148 15966 25268 15994
rect 25332 15994 25360 17575
rect 25424 16232 25452 23559
rect 28262 23520 28318 24000
rect 25594 22400 25650 22409
rect 25594 22335 25650 22344
rect 25608 19802 25636 22335
rect 25956 21788 26252 21808
rect 26012 21786 26036 21788
rect 26092 21786 26116 21788
rect 26172 21786 26196 21788
rect 26034 21734 26036 21786
rect 26098 21734 26110 21786
rect 26172 21734 26174 21786
rect 26012 21732 26036 21734
rect 26092 21732 26116 21734
rect 26172 21732 26196 21734
rect 25956 21712 26252 21732
rect 25870 21584 25926 21593
rect 25870 21519 25926 21528
rect 25778 20496 25834 20505
rect 25778 20431 25834 20440
rect 25608 19774 25728 19802
rect 25596 19712 25648 19718
rect 25596 19654 25648 19660
rect 25608 19310 25636 19654
rect 25596 19304 25648 19310
rect 25596 19246 25648 19252
rect 25424 16204 25636 16232
rect 25502 16144 25558 16153
rect 25502 16079 25558 16088
rect 25332 15966 25452 15994
rect 25042 14920 25098 14929
rect 25042 14855 25098 14864
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 25056 14618 25084 14758
rect 25044 14612 25096 14618
rect 25044 14554 25096 14560
rect 25056 13530 25084 14554
rect 25044 13524 25096 13530
rect 25044 13466 25096 13472
rect 25042 13016 25098 13025
rect 25042 12951 25098 12960
rect 25056 12782 25084 12951
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 25044 12640 25096 12646
rect 25148 12617 25176 15966
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 25240 15026 25268 15846
rect 25228 15020 25280 15026
rect 25228 14962 25280 14968
rect 25240 14074 25268 14962
rect 25424 14550 25452 15966
rect 25412 14544 25464 14550
rect 25412 14486 25464 14492
rect 25228 14068 25280 14074
rect 25228 14010 25280 14016
rect 25228 13388 25280 13394
rect 25228 13330 25280 13336
rect 25240 12986 25268 13330
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25228 12980 25280 12986
rect 25228 12922 25280 12928
rect 25332 12918 25360 13262
rect 25516 13190 25544 16079
rect 25504 13184 25556 13190
rect 25504 13126 25556 13132
rect 25320 12912 25372 12918
rect 25320 12854 25372 12860
rect 25320 12708 25372 12714
rect 25320 12650 25372 12656
rect 25044 12582 25096 12588
rect 25134 12608 25190 12617
rect 24768 12436 24820 12442
rect 24768 12378 24820 12384
rect 24952 12436 25004 12442
rect 24952 12378 25004 12384
rect 24492 12232 24544 12238
rect 24492 12174 24544 12180
rect 24400 9920 24452 9926
rect 24400 9862 24452 9868
rect 24504 9654 24532 12174
rect 24596 9654 24624 12310
rect 24688 12294 24992 12322
rect 24768 12164 24820 12170
rect 24768 12106 24820 12112
rect 24780 11694 24808 12106
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24872 11694 24900 12038
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24780 11354 24808 11630
rect 24768 11348 24820 11354
rect 24768 11290 24820 11296
rect 24964 10985 24992 12294
rect 25056 12209 25084 12582
rect 25134 12543 25190 12552
rect 25228 12300 25280 12306
rect 25228 12242 25280 12248
rect 25240 12209 25268 12242
rect 25042 12200 25098 12209
rect 25042 12135 25098 12144
rect 25226 12200 25282 12209
rect 25226 12135 25282 12144
rect 25042 12064 25098 12073
rect 25042 11999 25098 12008
rect 24950 10976 25006 10985
rect 24950 10911 25006 10920
rect 24860 10192 24912 10198
rect 24860 10134 24912 10140
rect 24308 9648 24360 9654
rect 24308 9590 24360 9596
rect 24492 9648 24544 9654
rect 24492 9590 24544 9596
rect 24584 9648 24636 9654
rect 24584 9590 24636 9596
rect 24216 9580 24268 9586
rect 24216 9522 24268 9528
rect 24124 9376 24176 9382
rect 24044 9336 24124 9364
rect 24124 9318 24176 9324
rect 24136 9081 24164 9318
rect 24122 9072 24178 9081
rect 24122 9007 24178 9016
rect 24228 8974 24256 9522
rect 24216 8968 24268 8974
rect 24216 8910 24268 8916
rect 24228 8838 24256 8910
rect 24216 8832 24268 8838
rect 24216 8774 24268 8780
rect 24228 8498 24256 8774
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 24124 8084 24176 8090
rect 24124 8026 24176 8032
rect 23952 7942 24072 7970
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23952 7206 23980 7822
rect 23940 7200 23992 7206
rect 23940 7142 23992 7148
rect 23846 6216 23902 6225
rect 23846 6151 23902 6160
rect 23860 5710 23888 6151
rect 23848 5704 23900 5710
rect 23754 5672 23810 5681
rect 23848 5646 23900 5652
rect 23754 5607 23810 5616
rect 23848 5568 23900 5574
rect 23952 5545 23980 7142
rect 23848 5510 23900 5516
rect 23938 5536 23994 5545
rect 22468 5296 22520 5302
rect 22468 5238 22520 5244
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 23572 5024 23624 5030
rect 23572 4966 23624 4972
rect 23584 4690 23612 4966
rect 23860 4690 23888 5510
rect 23938 5471 23994 5480
rect 23952 5137 23980 5471
rect 23938 5128 23994 5137
rect 23938 5063 23994 5072
rect 23572 4684 23624 4690
rect 23572 4626 23624 4632
rect 23848 4684 23900 4690
rect 23848 4626 23900 4632
rect 23584 4282 23612 4626
rect 23572 4276 23624 4282
rect 23572 4218 23624 4224
rect 23860 4078 23888 4626
rect 23848 4072 23900 4078
rect 23846 4040 23848 4049
rect 23900 4040 23902 4049
rect 23846 3975 23902 3984
rect 23846 2952 23902 2961
rect 23846 2887 23902 2896
rect 23860 2854 23888 2887
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 24044 2514 24072 7942
rect 24136 7002 24164 8026
rect 24228 8022 24256 8434
rect 24492 8356 24544 8362
rect 24492 8298 24544 8304
rect 24400 8288 24452 8294
rect 24400 8230 24452 8236
rect 24216 8016 24268 8022
rect 24216 7958 24268 7964
rect 24412 7546 24440 8230
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 24216 7472 24268 7478
rect 24214 7440 24216 7449
rect 24268 7440 24270 7449
rect 24214 7375 24270 7384
rect 24228 7342 24256 7375
rect 24216 7336 24268 7342
rect 24216 7278 24268 7284
rect 24124 6996 24176 7002
rect 24124 6938 24176 6944
rect 24136 6497 24164 6938
rect 24400 6860 24452 6866
rect 24400 6802 24452 6808
rect 24122 6488 24178 6497
rect 24412 6458 24440 6802
rect 24504 6730 24532 8298
rect 24768 8084 24820 8090
rect 24872 8072 24900 10134
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 24820 8044 24900 8072
rect 24768 8026 24820 8032
rect 24964 7002 24992 9590
rect 25056 9110 25084 11999
rect 25240 11898 25268 12135
rect 25228 11892 25280 11898
rect 25228 11834 25280 11840
rect 25226 11520 25282 11529
rect 25226 11455 25282 11464
rect 25044 9104 25096 9110
rect 25044 9046 25096 9052
rect 25240 7993 25268 11455
rect 25332 11218 25360 12650
rect 25412 12368 25464 12374
rect 25412 12310 25464 12316
rect 25320 11212 25372 11218
rect 25320 11154 25372 11160
rect 25332 10810 25360 11154
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 25226 7984 25282 7993
rect 25226 7919 25282 7928
rect 25044 7744 25096 7750
rect 25044 7686 25096 7692
rect 25056 7410 25084 7686
rect 25044 7404 25096 7410
rect 25044 7346 25096 7352
rect 24768 6996 24820 7002
rect 24768 6938 24820 6944
rect 24952 6996 25004 7002
rect 24952 6938 25004 6944
rect 24492 6724 24544 6730
rect 24492 6666 24544 6672
rect 24122 6423 24178 6432
rect 24400 6452 24452 6458
rect 24400 6394 24452 6400
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24688 2582 24716 6394
rect 24780 6118 24808 6938
rect 25056 6798 25084 7346
rect 25044 6792 25096 6798
rect 25044 6734 25096 6740
rect 25056 6458 25084 6734
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 24780 5409 24808 6054
rect 24766 5400 24822 5409
rect 24766 5335 24822 5344
rect 24952 5024 25004 5030
rect 24952 4966 25004 4972
rect 24964 4593 24992 4966
rect 24950 4584 25006 4593
rect 24950 4519 24952 4528
rect 25004 4519 25006 4528
rect 24952 4490 25004 4496
rect 24858 3768 24914 3777
rect 24858 3703 24914 3712
rect 24676 2576 24728 2582
rect 24676 2518 24728 2524
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 24032 2508 24084 2514
rect 24032 2450 24084 2456
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 24216 2440 24268 2446
rect 24216 2382 24268 2388
rect 22006 1456 22062 1465
rect 22006 1391 22062 1400
rect 22020 480 22048 1391
rect 23492 480 23520 2382
rect 24228 1465 24256 2382
rect 24214 1456 24270 1465
rect 24214 1391 24270 1400
rect 24872 480 24900 3703
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 25332 3097 25360 3538
rect 25424 3194 25452 12310
rect 25608 12306 25636 16204
rect 25596 12300 25648 12306
rect 25596 12242 25648 12248
rect 25502 11384 25558 11393
rect 25608 11370 25636 12242
rect 25558 11342 25636 11370
rect 25700 11354 25728 19774
rect 25792 15609 25820 20431
rect 25884 19242 25912 21519
rect 25956 20700 26252 20720
rect 26012 20698 26036 20700
rect 26092 20698 26116 20700
rect 26172 20698 26196 20700
rect 26034 20646 26036 20698
rect 26098 20646 26110 20698
rect 26172 20646 26174 20698
rect 26012 20644 26036 20646
rect 26092 20644 26116 20646
rect 26172 20644 26196 20646
rect 25956 20624 26252 20644
rect 26330 20360 26386 20369
rect 26330 20295 26386 20304
rect 26344 20262 26372 20295
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 26884 20256 26936 20262
rect 26884 20198 26936 20204
rect 26792 19916 26844 19922
rect 26792 19858 26844 19864
rect 25956 19612 26252 19632
rect 26012 19610 26036 19612
rect 26092 19610 26116 19612
rect 26172 19610 26196 19612
rect 26034 19558 26036 19610
rect 26098 19558 26110 19610
rect 26172 19558 26174 19610
rect 26012 19556 26036 19558
rect 26092 19556 26116 19558
rect 26172 19556 26196 19558
rect 25956 19536 26252 19556
rect 26148 19372 26200 19378
rect 26148 19314 26200 19320
rect 26160 19258 26188 19314
rect 25872 19236 25924 19242
rect 26160 19230 26372 19258
rect 25872 19178 25924 19184
rect 25956 18524 26252 18544
rect 26012 18522 26036 18524
rect 26092 18522 26116 18524
rect 26172 18522 26196 18524
rect 26034 18470 26036 18522
rect 26098 18470 26110 18522
rect 26172 18470 26174 18522
rect 26012 18468 26036 18470
rect 26092 18468 26116 18470
rect 26172 18468 26196 18470
rect 25956 18448 26252 18468
rect 26344 18426 26372 19230
rect 26804 19174 26832 19858
rect 26792 19168 26844 19174
rect 26792 19110 26844 19116
rect 26332 18420 26384 18426
rect 26332 18362 26384 18368
rect 26148 18216 26200 18222
rect 26148 18158 26200 18164
rect 26160 17898 26188 18158
rect 26514 17912 26570 17921
rect 26160 17882 26280 17898
rect 26160 17876 26292 17882
rect 26160 17870 26240 17876
rect 26514 17847 26570 17856
rect 26240 17818 26292 17824
rect 26252 17626 26280 17818
rect 26422 17776 26478 17785
rect 26422 17711 26478 17720
rect 26252 17598 26372 17626
rect 25956 17436 26252 17456
rect 26012 17434 26036 17436
rect 26092 17434 26116 17436
rect 26172 17434 26196 17436
rect 26034 17382 26036 17434
rect 26098 17382 26110 17434
rect 26172 17382 26174 17434
rect 26012 17380 26036 17382
rect 26092 17380 26116 17382
rect 26172 17380 26196 17382
rect 25956 17360 26252 17380
rect 25872 16992 25924 16998
rect 25872 16934 25924 16940
rect 25778 15600 25834 15609
rect 25778 15535 25834 15544
rect 25778 15464 25834 15473
rect 25778 15399 25834 15408
rect 25792 13841 25820 15399
rect 25778 13832 25834 13841
rect 25778 13767 25834 13776
rect 25778 13696 25834 13705
rect 25778 13631 25834 13640
rect 25792 12782 25820 13631
rect 25780 12776 25832 12782
rect 25780 12718 25832 12724
rect 25778 12608 25834 12617
rect 25778 12543 25834 12552
rect 25792 11801 25820 12543
rect 25778 11792 25834 11801
rect 25778 11727 25834 11736
rect 25780 11620 25832 11626
rect 25780 11562 25832 11568
rect 25688 11348 25740 11354
rect 25502 11319 25558 11328
rect 25516 11286 25544 11319
rect 25688 11290 25740 11296
rect 25504 11280 25556 11286
rect 25504 11222 25556 11228
rect 25596 11280 25648 11286
rect 25596 11222 25648 11228
rect 25504 11076 25556 11082
rect 25504 11018 25556 11024
rect 25516 6905 25544 11018
rect 25608 7546 25636 11222
rect 25688 9512 25740 9518
rect 25688 9454 25740 9460
rect 25700 8838 25728 9454
rect 25688 8832 25740 8838
rect 25688 8774 25740 8780
rect 25700 7750 25728 8774
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25608 7274 25636 7482
rect 25700 7410 25728 7686
rect 25688 7404 25740 7410
rect 25688 7346 25740 7352
rect 25596 7268 25648 7274
rect 25596 7210 25648 7216
rect 25502 6896 25558 6905
rect 25502 6831 25558 6840
rect 25504 5568 25556 5574
rect 25700 5556 25728 7346
rect 25792 6225 25820 11562
rect 25884 11121 25912 16934
rect 25956 16348 26252 16368
rect 26012 16346 26036 16348
rect 26092 16346 26116 16348
rect 26172 16346 26196 16348
rect 26034 16294 26036 16346
rect 26098 16294 26110 16346
rect 26172 16294 26174 16346
rect 26012 16292 26036 16294
rect 26092 16292 26116 16294
rect 26172 16292 26196 16294
rect 25956 16272 26252 16292
rect 26344 16164 26372 17598
rect 26436 17134 26464 17711
rect 26424 17128 26476 17134
rect 26424 17070 26476 17076
rect 25976 16136 26372 16164
rect 25976 16046 26004 16136
rect 25964 16040 26016 16046
rect 25964 15982 26016 15988
rect 25976 15706 26004 15982
rect 25964 15700 26016 15706
rect 25964 15642 26016 15648
rect 26160 15450 26188 16136
rect 26528 15570 26556 17847
rect 26516 15564 26568 15570
rect 26516 15506 26568 15512
rect 26160 15422 26372 15450
rect 25956 15260 26252 15280
rect 26012 15258 26036 15260
rect 26092 15258 26116 15260
rect 26172 15258 26196 15260
rect 26034 15206 26036 15258
rect 26098 15206 26110 15258
rect 26172 15206 26174 15258
rect 26012 15204 26036 15206
rect 26092 15204 26116 15206
rect 26172 15204 26196 15206
rect 25956 15184 26252 15204
rect 26148 14884 26200 14890
rect 26148 14826 26200 14832
rect 26160 14634 26188 14826
rect 26344 14770 26372 15422
rect 26528 15162 26556 15506
rect 26516 15156 26568 15162
rect 26516 15098 26568 15104
rect 26344 14742 26464 14770
rect 26160 14606 26372 14634
rect 25956 14172 26252 14192
rect 26012 14170 26036 14172
rect 26092 14170 26116 14172
rect 26172 14170 26196 14172
rect 26034 14118 26036 14170
rect 26098 14118 26110 14170
rect 26172 14118 26174 14170
rect 26012 14116 26036 14118
rect 26092 14116 26116 14118
rect 26172 14116 26196 14118
rect 25956 14096 26252 14116
rect 26146 13968 26202 13977
rect 26146 13903 26202 13912
rect 26160 13870 26188 13903
rect 26148 13864 26200 13870
rect 26200 13812 26280 13818
rect 26148 13806 26280 13812
rect 26160 13790 26280 13806
rect 26056 13728 26108 13734
rect 26056 13670 26108 13676
rect 26068 13326 26096 13670
rect 26252 13530 26280 13790
rect 26240 13524 26292 13530
rect 26240 13466 26292 13472
rect 26056 13320 26108 13326
rect 26056 13262 26108 13268
rect 25956 13084 26252 13104
rect 26012 13082 26036 13084
rect 26092 13082 26116 13084
rect 26172 13082 26196 13084
rect 26034 13030 26036 13082
rect 26098 13030 26110 13082
rect 26172 13030 26174 13082
rect 26012 13028 26036 13030
rect 26092 13028 26116 13030
rect 26172 13028 26196 13030
rect 25956 13008 26252 13028
rect 26056 12844 26108 12850
rect 26056 12786 26108 12792
rect 26068 12170 26096 12786
rect 26056 12164 26108 12170
rect 26056 12106 26108 12112
rect 25956 11996 26252 12016
rect 26012 11994 26036 11996
rect 26092 11994 26116 11996
rect 26172 11994 26196 11996
rect 26034 11942 26036 11994
rect 26098 11942 26110 11994
rect 26172 11942 26174 11994
rect 26012 11940 26036 11942
rect 26092 11940 26116 11942
rect 26172 11940 26196 11942
rect 25956 11920 26252 11940
rect 26344 11898 26372 14606
rect 26436 13530 26464 14742
rect 26424 13524 26476 13530
rect 26424 13466 26476 13472
rect 26516 13320 26568 13326
rect 26516 13262 26568 13268
rect 26528 12442 26556 13262
rect 26516 12436 26568 12442
rect 26516 12378 26568 12384
rect 26700 12436 26752 12442
rect 26700 12378 26752 12384
rect 26424 12368 26476 12374
rect 26424 12310 26476 12316
rect 26332 11892 26384 11898
rect 26332 11834 26384 11840
rect 26436 11830 26464 12310
rect 26516 12300 26568 12306
rect 26516 12242 26568 12248
rect 26424 11824 26476 11830
rect 26424 11766 26476 11772
rect 26528 11558 26556 12242
rect 26712 11762 26740 12378
rect 26700 11756 26752 11762
rect 26700 11698 26752 11704
rect 26698 11656 26754 11665
rect 26698 11591 26754 11600
rect 26516 11552 26568 11558
rect 26516 11494 26568 11500
rect 26528 11218 26556 11494
rect 26712 11354 26740 11591
rect 26700 11348 26752 11354
rect 26700 11290 26752 11296
rect 26516 11212 26568 11218
rect 26516 11154 26568 11160
rect 25870 11112 25926 11121
rect 25870 11047 25926 11056
rect 25956 10908 26252 10928
rect 26012 10906 26036 10908
rect 26092 10906 26116 10908
rect 26172 10906 26196 10908
rect 26034 10854 26036 10906
rect 26098 10854 26110 10906
rect 26172 10854 26174 10906
rect 26012 10852 26036 10854
rect 26092 10852 26116 10854
rect 26172 10852 26196 10854
rect 25956 10832 26252 10852
rect 26528 10810 26556 11154
rect 26516 10804 26568 10810
rect 26516 10746 26568 10752
rect 26528 10169 26556 10746
rect 26608 10464 26660 10470
rect 26606 10432 26608 10441
rect 26660 10432 26662 10441
rect 26606 10367 26662 10376
rect 26514 10160 26570 10169
rect 26424 10124 26476 10130
rect 26514 10095 26570 10104
rect 26424 10066 26476 10072
rect 26436 10033 26464 10066
rect 26422 10024 26478 10033
rect 26478 9982 26556 10010
rect 26422 9959 26478 9968
rect 25956 9820 26252 9840
rect 26012 9818 26036 9820
rect 26092 9818 26116 9820
rect 26172 9818 26196 9820
rect 26034 9766 26036 9818
rect 26098 9766 26110 9818
rect 26172 9766 26174 9818
rect 26012 9764 26036 9766
rect 26092 9764 26116 9766
rect 26172 9764 26196 9766
rect 25956 9744 26252 9764
rect 26528 9722 26556 9982
rect 26700 9920 26752 9926
rect 26698 9888 26700 9897
rect 26752 9888 26754 9897
rect 26698 9823 26754 9832
rect 26516 9716 26568 9722
rect 26516 9658 26568 9664
rect 26698 9344 26754 9353
rect 26698 9279 26754 9288
rect 26712 9178 26740 9279
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26424 9036 26476 9042
rect 26424 8978 26476 8984
rect 25956 8732 26252 8752
rect 26012 8730 26036 8732
rect 26092 8730 26116 8732
rect 26172 8730 26196 8732
rect 26034 8678 26036 8730
rect 26098 8678 26110 8730
rect 26172 8678 26174 8730
rect 26012 8676 26036 8678
rect 26092 8676 26116 8678
rect 26172 8676 26196 8678
rect 25956 8656 26252 8676
rect 26436 8362 26464 8978
rect 26698 8664 26754 8673
rect 26698 8599 26754 8608
rect 26424 8356 26476 8362
rect 26424 8298 26476 8304
rect 25872 7948 25924 7954
rect 25872 7890 25924 7896
rect 25884 7528 25912 7890
rect 25956 7644 26252 7664
rect 26012 7642 26036 7644
rect 26092 7642 26116 7644
rect 26172 7642 26196 7644
rect 26034 7590 26036 7642
rect 26098 7590 26110 7642
rect 26172 7590 26174 7642
rect 26012 7588 26036 7590
rect 26092 7588 26116 7590
rect 26172 7588 26196 7590
rect 25956 7568 26252 7588
rect 25884 7500 26004 7528
rect 25976 7342 26004 7500
rect 26330 7440 26386 7449
rect 26330 7375 26386 7384
rect 25964 7336 26016 7342
rect 25962 7304 25964 7313
rect 26016 7304 26018 7313
rect 25962 7239 26018 7248
rect 25956 6556 26252 6576
rect 26012 6554 26036 6556
rect 26092 6554 26116 6556
rect 26172 6554 26196 6556
rect 26034 6502 26036 6554
rect 26098 6502 26110 6554
rect 26172 6502 26174 6554
rect 26012 6500 26036 6502
rect 26092 6500 26116 6502
rect 26172 6500 26196 6502
rect 25956 6480 26252 6500
rect 26238 6352 26294 6361
rect 26238 6287 26240 6296
rect 26292 6287 26294 6296
rect 26240 6258 26292 6264
rect 25778 6216 25834 6225
rect 25778 6151 25834 6160
rect 25556 5528 25728 5556
rect 25504 5510 25556 5516
rect 25516 5166 25544 5510
rect 25956 5468 26252 5488
rect 26012 5466 26036 5468
rect 26092 5466 26116 5468
rect 26172 5466 26196 5468
rect 26034 5414 26036 5466
rect 26098 5414 26110 5466
rect 26172 5414 26174 5466
rect 26012 5412 26036 5414
rect 26092 5412 26116 5414
rect 26172 5412 26196 5414
rect 25956 5392 26252 5412
rect 25504 5160 25556 5166
rect 25504 5102 25556 5108
rect 25956 4380 26252 4400
rect 26012 4378 26036 4380
rect 26092 4378 26116 4380
rect 26172 4378 26196 4380
rect 26034 4326 26036 4378
rect 26098 4326 26110 4378
rect 26172 4326 26174 4378
rect 26012 4324 26036 4326
rect 26092 4324 26116 4326
rect 26172 4324 26196 4326
rect 25956 4304 26252 4324
rect 26344 4078 26372 7375
rect 26436 5273 26464 8298
rect 26712 8090 26740 8599
rect 26700 8084 26752 8090
rect 26700 8026 26752 8032
rect 26804 7750 26832 19110
rect 26792 7744 26844 7750
rect 26792 7686 26844 7692
rect 26698 7440 26754 7449
rect 26698 7375 26754 7384
rect 26712 6730 26740 7375
rect 26792 7268 26844 7274
rect 26792 7210 26844 7216
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 26804 6662 26832 7210
rect 26792 6656 26844 6662
rect 26792 6598 26844 6604
rect 26804 6458 26832 6598
rect 26792 6452 26844 6458
rect 26792 6394 26844 6400
rect 26608 6112 26660 6118
rect 26608 6054 26660 6060
rect 26514 5808 26570 5817
rect 26514 5743 26516 5752
rect 26568 5743 26570 5752
rect 26516 5714 26568 5720
rect 26528 5370 26556 5714
rect 26620 5681 26648 6054
rect 26606 5672 26662 5681
rect 26606 5607 26662 5616
rect 26700 5568 26752 5574
rect 26700 5510 26752 5516
rect 26516 5364 26568 5370
rect 26516 5306 26568 5312
rect 26422 5264 26478 5273
rect 26422 5199 26478 5208
rect 26712 5137 26740 5510
rect 26804 5302 26832 6394
rect 26792 5296 26844 5302
rect 26792 5238 26844 5244
rect 26514 5128 26570 5137
rect 26514 5063 26570 5072
rect 26698 5128 26754 5137
rect 26698 5063 26754 5072
rect 26528 4690 26556 5063
rect 26516 4684 26568 4690
rect 26516 4626 26568 4632
rect 26700 4480 26752 4486
rect 26700 4422 26752 4428
rect 26712 4185 26740 4422
rect 26698 4176 26754 4185
rect 26698 4111 26754 4120
rect 26332 4072 26384 4078
rect 26332 4014 26384 4020
rect 26608 4072 26660 4078
rect 26896 4049 26924 20198
rect 28276 20058 28304 23520
rect 28264 20052 28316 20058
rect 28264 19994 28316 20000
rect 26974 18864 27030 18873
rect 26974 18799 27030 18808
rect 26988 13569 27016 18799
rect 27344 17060 27396 17066
rect 27344 17002 27396 17008
rect 27252 15360 27304 15366
rect 27252 15302 27304 15308
rect 26974 13560 27030 13569
rect 26974 13495 27030 13504
rect 26988 12442 27016 13495
rect 26976 12436 27028 12442
rect 26976 12378 27028 12384
rect 27068 12232 27120 12238
rect 27068 12174 27120 12180
rect 27080 11354 27108 12174
rect 27160 12096 27212 12102
rect 27160 12038 27212 12044
rect 27172 11762 27200 12038
rect 27160 11756 27212 11762
rect 27160 11698 27212 11704
rect 27172 11354 27200 11698
rect 27264 11626 27292 15302
rect 27356 12345 27384 17002
rect 27434 15872 27490 15881
rect 27434 15807 27490 15816
rect 27342 12336 27398 12345
rect 27342 12271 27398 12280
rect 27252 11620 27304 11626
rect 27252 11562 27304 11568
rect 27068 11348 27120 11354
rect 27068 11290 27120 11296
rect 27160 11348 27212 11354
rect 27160 11290 27212 11296
rect 27356 11286 27384 12271
rect 27344 11280 27396 11286
rect 27344 11222 27396 11228
rect 27448 10198 27476 15807
rect 27618 12200 27674 12209
rect 27618 12135 27674 12144
rect 27528 12096 27580 12102
rect 27528 12038 27580 12044
rect 27540 11694 27568 12038
rect 27528 11688 27580 11694
rect 27528 11630 27580 11636
rect 27632 11354 27660 12135
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 27526 10704 27582 10713
rect 27526 10639 27582 10648
rect 27540 10606 27568 10639
rect 27528 10600 27580 10606
rect 27528 10542 27580 10548
rect 27712 10464 27764 10470
rect 27712 10406 27764 10412
rect 27436 10192 27488 10198
rect 27436 10134 27488 10140
rect 26976 9648 27028 9654
rect 26974 9616 26976 9625
rect 27028 9616 27030 9625
rect 26974 9551 27030 9560
rect 27528 9444 27580 9450
rect 27528 9386 27580 9392
rect 27068 7744 27120 7750
rect 27068 7686 27120 7692
rect 26976 6860 27028 6866
rect 26976 6802 27028 6808
rect 26988 6458 27016 6802
rect 26976 6452 27028 6458
rect 26976 6394 27028 6400
rect 26608 4014 26660 4020
rect 26882 4040 26938 4049
rect 26620 3913 26648 4014
rect 26882 3975 26938 3984
rect 26700 3936 26752 3942
rect 26606 3904 26662 3913
rect 26700 3878 26752 3884
rect 26606 3839 26662 3848
rect 25502 3496 25558 3505
rect 26712 3482 26740 3878
rect 27080 3777 27108 7686
rect 27540 7546 27568 9386
rect 27724 8129 27752 10406
rect 27710 8120 27766 8129
rect 27710 8055 27766 8064
rect 27528 7540 27580 7546
rect 27528 7482 27580 7488
rect 27436 5704 27488 5710
rect 27436 5646 27488 5652
rect 27160 4684 27212 4690
rect 27160 4626 27212 4632
rect 27172 4282 27200 4626
rect 27160 4276 27212 4282
rect 27160 4218 27212 4224
rect 27066 3768 27122 3777
rect 27066 3703 27122 3712
rect 27344 3596 27396 3602
rect 27344 3538 27396 3544
rect 26712 3454 26832 3482
rect 25502 3431 25504 3440
rect 25556 3431 25558 3440
rect 25504 3402 25556 3408
rect 26700 3392 26752 3398
rect 26700 3334 26752 3340
rect 25956 3292 26252 3312
rect 26012 3290 26036 3292
rect 26092 3290 26116 3292
rect 26172 3290 26196 3292
rect 26034 3238 26036 3290
rect 26098 3238 26110 3290
rect 26172 3238 26174 3290
rect 26012 3236 26036 3238
rect 26092 3236 26116 3238
rect 26172 3236 26196 3238
rect 25956 3216 26252 3236
rect 25412 3188 25464 3194
rect 25412 3130 25464 3136
rect 26332 3120 26384 3126
rect 25318 3088 25374 3097
rect 26332 3062 26384 3068
rect 26422 3088 26478 3097
rect 25318 3023 25320 3032
rect 25372 3023 25374 3032
rect 25320 2994 25372 3000
rect 25872 2304 25924 2310
rect 25872 2246 25924 2252
rect 25884 1465 25912 2246
rect 25956 2204 26252 2224
rect 26012 2202 26036 2204
rect 26092 2202 26116 2204
rect 26172 2202 26196 2204
rect 26034 2150 26036 2202
rect 26098 2150 26110 2202
rect 26172 2150 26174 2202
rect 26012 2148 26036 2150
rect 26092 2148 26116 2150
rect 26172 2148 26196 2150
rect 25956 2128 26252 2148
rect 25870 1456 25926 1465
rect 25870 1391 25926 1400
rect 26344 480 26372 3062
rect 26422 3023 26478 3032
rect 26436 2990 26464 3023
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 26608 2848 26660 2854
rect 26608 2790 26660 2796
rect 26620 921 26648 2790
rect 26712 2145 26740 3334
rect 26698 2136 26754 2145
rect 26698 2071 26754 2080
rect 26606 912 26662 921
rect 26606 847 26662 856
rect 1398 368 1454 377
rect 1398 303 1454 312
rect 2042 0 2098 480
rect 3514 0 3570 480
rect 4894 0 4950 480
rect 6366 0 6422 480
rect 7746 0 7802 480
rect 9218 0 9274 480
rect 10598 0 10654 480
rect 12070 0 12126 480
rect 13450 0 13506 480
rect 14922 0 14978 480
rect 16302 0 16358 480
rect 17774 0 17830 480
rect 19154 0 19210 480
rect 20626 0 20682 480
rect 22006 0 22062 480
rect 23478 0 23534 480
rect 24858 0 24914 480
rect 26330 0 26386 480
rect 26804 377 26832 3454
rect 27356 3194 27384 3538
rect 27344 3188 27396 3194
rect 27344 3130 27396 3136
rect 27448 2990 27476 5646
rect 27526 4448 27582 4457
rect 27526 4383 27582 4392
rect 27540 3942 27568 4383
rect 27618 4040 27674 4049
rect 27618 3975 27674 3984
rect 27528 3936 27580 3942
rect 27528 3878 27580 3884
rect 27436 2984 27488 2990
rect 27436 2926 27488 2932
rect 27632 2666 27660 3975
rect 27712 2848 27764 2854
rect 27710 2816 27712 2825
rect 27764 2816 27766 2825
rect 27710 2751 27766 2760
rect 27632 2638 27752 2666
rect 27724 480 27752 2638
rect 29184 2304 29236 2310
rect 29184 2246 29236 2252
rect 29196 480 29224 2246
rect 26790 368 26846 377
rect 26790 303 26846 312
rect 27710 0 27766 480
rect 29182 0 29238 480
<< via2 >>
rect 3330 23568 3386 23624
rect 2778 22344 2834 22400
rect 2042 18672 2098 18728
rect 754 15272 810 15328
rect 1858 12588 1860 12608
rect 1860 12588 1912 12608
rect 1912 12588 1914 12608
rect 1858 12552 1914 12588
rect 1582 11056 1638 11112
rect 1582 10412 1584 10432
rect 1584 10412 1636 10432
rect 1636 10412 1638 10432
rect 1582 10376 1638 10412
rect 1582 9324 1584 9344
rect 1584 9324 1636 9344
rect 1636 9324 1638 9344
rect 1582 9288 1638 9324
rect 1490 8608 1546 8664
rect 1582 8064 1638 8120
rect 1398 7384 1454 7440
rect 1582 6840 1638 6896
rect 662 3576 718 3632
rect 1582 5616 1638 5672
rect 1582 5072 1638 5128
rect 1490 4392 1546 4448
rect 1582 3848 1638 3904
rect 2318 17856 2374 17912
rect 2318 16904 2374 16960
rect 2686 16904 2742 16960
rect 2318 12008 2374 12064
rect 2134 11736 2190 11792
rect 2042 9036 2098 9072
rect 2042 9016 2044 9036
rect 2044 9016 2096 9036
rect 2096 9016 2098 9036
rect 1950 7384 2006 7440
rect 25410 23568 25466 23624
rect 4158 23024 4214 23080
rect 4066 21800 4122 21856
rect 3974 21256 4030 21312
rect 3790 20576 3846 20632
rect 3330 20032 3386 20088
rect 2962 18808 3018 18864
rect 2870 16632 2926 16688
rect 3054 18028 3056 18048
rect 3056 18028 3108 18048
rect 3108 18028 3110 18048
rect 3054 17992 3110 18028
rect 3606 18264 3662 18320
rect 3606 17584 3662 17640
rect 3330 13504 3386 13560
rect 3606 13368 3662 13424
rect 3054 12552 3110 12608
rect 2778 11464 2834 11520
rect 2778 11192 2834 11248
rect 2686 9832 2742 9888
rect 3146 12280 3202 12336
rect 3606 12688 3662 12744
rect 3514 11600 3570 11656
rect 2962 11056 3018 11112
rect 3698 10512 3754 10568
rect 2962 9444 3018 9480
rect 2962 9424 2964 9444
rect 2964 9424 3016 9444
rect 3016 9424 3018 9444
rect 3146 9596 3148 9616
rect 3148 9596 3200 9616
rect 3200 9596 3202 9616
rect 3146 9560 3202 9596
rect 3054 8880 3110 8936
rect 2410 8492 2466 8528
rect 2410 8472 2412 8492
rect 2412 8472 2464 8492
rect 2464 8472 2466 8492
rect 2042 6704 2098 6760
rect 1858 6296 1914 6352
rect 2226 5480 2282 5536
rect 2042 4684 2098 4720
rect 2042 4664 2044 4684
rect 2044 4664 2096 4684
rect 2096 4664 2098 4684
rect 2134 4120 2190 4176
rect 2042 4004 2098 4040
rect 2042 3984 2044 4004
rect 2044 3984 2096 4004
rect 2096 3984 2098 4004
rect 1582 1400 1638 1456
rect 4066 20032 4122 20088
rect 5956 21786 6012 21788
rect 6036 21786 6092 21788
rect 6116 21786 6172 21788
rect 6196 21786 6252 21788
rect 5956 21734 5982 21786
rect 5982 21734 6012 21786
rect 6036 21734 6046 21786
rect 6046 21734 6092 21786
rect 6116 21734 6162 21786
rect 6162 21734 6172 21786
rect 6196 21734 6226 21786
rect 6226 21734 6252 21786
rect 5956 21732 6012 21734
rect 6036 21732 6092 21734
rect 6116 21732 6172 21734
rect 6196 21732 6252 21734
rect 5956 20698 6012 20700
rect 6036 20698 6092 20700
rect 6116 20698 6172 20700
rect 6196 20698 6252 20700
rect 5956 20646 5982 20698
rect 5982 20646 6012 20698
rect 6036 20646 6046 20698
rect 6046 20646 6092 20698
rect 6116 20646 6162 20698
rect 6162 20646 6172 20698
rect 6196 20646 6226 20698
rect 6226 20646 6252 20698
rect 5956 20644 6012 20646
rect 6036 20644 6092 20646
rect 6116 20644 6172 20646
rect 6196 20644 6252 20646
rect 4986 20304 5042 20360
rect 4434 18844 4436 18864
rect 4436 18844 4488 18864
rect 4488 18844 4490 18864
rect 4434 18808 4490 18844
rect 4526 18708 4528 18728
rect 4528 18708 4580 18728
rect 4580 18708 4582 18728
rect 4526 18672 4582 18708
rect 4526 17584 4582 17640
rect 4434 17040 4490 17096
rect 4066 16768 4122 16824
rect 4250 15972 4306 16008
rect 4250 15952 4252 15972
rect 4252 15952 4304 15972
rect 4304 15952 4306 15972
rect 3882 15816 3938 15872
rect 3790 6976 3846 7032
rect 6642 20052 6698 20088
rect 6642 20032 6644 20052
rect 6644 20032 6696 20052
rect 6696 20032 6698 20052
rect 5956 19610 6012 19612
rect 6036 19610 6092 19612
rect 6116 19610 6172 19612
rect 6196 19610 6252 19612
rect 5956 19558 5982 19610
rect 5982 19558 6012 19610
rect 6036 19558 6046 19610
rect 6046 19558 6092 19610
rect 6116 19558 6162 19610
rect 6162 19558 6172 19610
rect 6196 19558 6226 19610
rect 6226 19558 6252 19610
rect 5956 19556 6012 19558
rect 6036 19556 6092 19558
rect 6116 19556 6172 19558
rect 6196 19556 6252 19558
rect 5956 18522 6012 18524
rect 6036 18522 6092 18524
rect 6116 18522 6172 18524
rect 6196 18522 6252 18524
rect 5956 18470 5982 18522
rect 5982 18470 6012 18522
rect 6036 18470 6046 18522
rect 6046 18470 6092 18522
rect 6116 18470 6162 18522
rect 6162 18470 6172 18522
rect 6196 18470 6226 18522
rect 6226 18470 6252 18522
rect 5956 18468 6012 18470
rect 6036 18468 6092 18470
rect 6116 18468 6172 18470
rect 6196 18468 6252 18470
rect 5630 17992 5686 18048
rect 4066 14068 4122 14104
rect 4066 14048 4068 14068
rect 4068 14048 4120 14068
rect 4120 14048 4122 14068
rect 3974 12144 4030 12200
rect 4250 12552 4306 12608
rect 4158 11872 4214 11928
rect 4710 13404 4712 13424
rect 4712 13404 4764 13424
rect 4764 13404 4766 13424
rect 4710 13368 4766 13404
rect 4710 12824 4766 12880
rect 4434 12008 4490 12064
rect 2502 3440 2558 3496
rect 4526 6704 4582 6760
rect 2778 3304 2834 3360
rect 2870 2624 2926 2680
rect 4710 5480 4766 5536
rect 4342 5208 4398 5264
rect 4710 5072 4766 5128
rect 2778 2080 2834 2136
rect 5956 17434 6012 17436
rect 6036 17434 6092 17436
rect 6116 17434 6172 17436
rect 6196 17434 6252 17436
rect 5956 17382 5982 17434
rect 5982 17382 6012 17434
rect 6036 17382 6046 17434
rect 6046 17382 6092 17434
rect 6116 17382 6162 17434
rect 6162 17382 6172 17434
rect 6196 17382 6226 17434
rect 6226 17382 6252 17434
rect 5956 17380 6012 17382
rect 6036 17380 6092 17382
rect 6116 17380 6172 17382
rect 6196 17380 6252 17382
rect 5722 16788 5778 16824
rect 5722 16768 5724 16788
rect 5724 16768 5776 16788
rect 5776 16768 5778 16788
rect 5538 16360 5594 16416
rect 5078 12860 5080 12880
rect 5080 12860 5132 12880
rect 5132 12860 5134 12880
rect 5078 12824 5134 12860
rect 5956 16346 6012 16348
rect 6036 16346 6092 16348
rect 6116 16346 6172 16348
rect 6196 16346 6252 16348
rect 5956 16294 5982 16346
rect 5982 16294 6012 16346
rect 6036 16294 6046 16346
rect 6046 16294 6092 16346
rect 6116 16294 6162 16346
rect 6162 16294 6172 16346
rect 6196 16294 6226 16346
rect 6226 16294 6252 16346
rect 5956 16292 6012 16294
rect 6036 16292 6092 16294
rect 6116 16292 6172 16294
rect 6196 16292 6252 16294
rect 5956 15258 6012 15260
rect 6036 15258 6092 15260
rect 6116 15258 6172 15260
rect 6196 15258 6252 15260
rect 5956 15206 5982 15258
rect 5982 15206 6012 15258
rect 6036 15206 6046 15258
rect 6046 15206 6092 15258
rect 6116 15206 6162 15258
rect 6162 15206 6172 15258
rect 6196 15206 6226 15258
rect 6226 15206 6252 15258
rect 5956 15204 6012 15206
rect 6036 15204 6092 15206
rect 6116 15204 6172 15206
rect 6196 15204 6252 15206
rect 5956 14170 6012 14172
rect 6036 14170 6092 14172
rect 6116 14170 6172 14172
rect 6196 14170 6252 14172
rect 5956 14118 5982 14170
rect 5982 14118 6012 14170
rect 6036 14118 6046 14170
rect 6046 14118 6092 14170
rect 6116 14118 6162 14170
rect 6162 14118 6172 14170
rect 6196 14118 6226 14170
rect 6226 14118 6252 14170
rect 5956 14116 6012 14118
rect 6036 14116 6092 14118
rect 6116 14116 6172 14118
rect 6196 14116 6252 14118
rect 5956 13082 6012 13084
rect 6036 13082 6092 13084
rect 6116 13082 6172 13084
rect 6196 13082 6252 13084
rect 5956 13030 5982 13082
rect 5982 13030 6012 13082
rect 6036 13030 6046 13082
rect 6046 13030 6092 13082
rect 6116 13030 6162 13082
rect 6162 13030 6172 13082
rect 6196 13030 6226 13082
rect 6226 13030 6252 13082
rect 5956 13028 6012 13030
rect 6036 13028 6092 13030
rect 6116 13028 6172 13030
rect 6196 13028 6252 13030
rect 5630 12280 5686 12336
rect 5956 11994 6012 11996
rect 6036 11994 6092 11996
rect 6116 11994 6172 11996
rect 6196 11994 6252 11996
rect 5956 11942 5982 11994
rect 5982 11942 6012 11994
rect 6036 11942 6046 11994
rect 6046 11942 6092 11994
rect 6116 11942 6162 11994
rect 6162 11942 6172 11994
rect 6196 11942 6226 11994
rect 6226 11942 6252 11994
rect 5956 11940 6012 11942
rect 6036 11940 6092 11942
rect 6116 11940 6172 11942
rect 6196 11940 6252 11942
rect 5956 10906 6012 10908
rect 6036 10906 6092 10908
rect 6116 10906 6172 10908
rect 6196 10906 6252 10908
rect 5956 10854 5982 10906
rect 5982 10854 6012 10906
rect 6036 10854 6046 10906
rect 6046 10854 6092 10906
rect 6116 10854 6162 10906
rect 6162 10854 6172 10906
rect 6196 10854 6226 10906
rect 6226 10854 6252 10906
rect 5956 10852 6012 10854
rect 6036 10852 6092 10854
rect 6116 10852 6172 10854
rect 6196 10852 6252 10854
rect 5956 9818 6012 9820
rect 6036 9818 6092 9820
rect 6116 9818 6172 9820
rect 6196 9818 6252 9820
rect 5956 9766 5982 9818
rect 5982 9766 6012 9818
rect 6036 9766 6046 9818
rect 6046 9766 6092 9818
rect 6116 9766 6162 9818
rect 6162 9766 6172 9818
rect 6196 9766 6226 9818
rect 6226 9766 6252 9818
rect 5956 9764 6012 9766
rect 6036 9764 6092 9766
rect 6116 9764 6172 9766
rect 6196 9764 6252 9766
rect 6550 9560 6606 9616
rect 5630 9288 5686 9344
rect 5956 8730 6012 8732
rect 6036 8730 6092 8732
rect 6116 8730 6172 8732
rect 6196 8730 6252 8732
rect 5956 8678 5982 8730
rect 5982 8678 6012 8730
rect 6036 8678 6046 8730
rect 6046 8678 6092 8730
rect 6116 8678 6162 8730
rect 6162 8678 6172 8730
rect 6196 8678 6226 8730
rect 6226 8678 6252 8730
rect 5956 8676 6012 8678
rect 6036 8676 6092 8678
rect 6116 8676 6172 8678
rect 6196 8676 6252 8678
rect 5956 7642 6012 7644
rect 6036 7642 6092 7644
rect 6116 7642 6172 7644
rect 6196 7642 6252 7644
rect 5956 7590 5982 7642
rect 5982 7590 6012 7642
rect 6036 7590 6046 7642
rect 6046 7590 6092 7642
rect 6116 7590 6162 7642
rect 6162 7590 6172 7642
rect 6196 7590 6226 7642
rect 6226 7590 6252 7642
rect 5956 7588 6012 7590
rect 6036 7588 6092 7590
rect 6116 7588 6172 7590
rect 6196 7588 6252 7590
rect 6642 7384 6698 7440
rect 5814 6976 5870 7032
rect 6182 6996 6238 7032
rect 6182 6976 6184 6996
rect 6184 6976 6236 6996
rect 6236 6976 6238 6996
rect 5956 6554 6012 6556
rect 6036 6554 6092 6556
rect 6116 6554 6172 6556
rect 6196 6554 6252 6556
rect 5956 6502 5982 6554
rect 5982 6502 6012 6554
rect 6036 6502 6046 6554
rect 6046 6502 6092 6554
rect 6116 6502 6162 6554
rect 6162 6502 6172 6554
rect 6196 6502 6226 6554
rect 6226 6502 6252 6554
rect 5956 6500 6012 6502
rect 6036 6500 6092 6502
rect 6116 6500 6172 6502
rect 6196 6500 6252 6502
rect 6274 6160 6330 6216
rect 4066 2760 4122 2816
rect 5956 5466 6012 5468
rect 6036 5466 6092 5468
rect 6116 5466 6172 5468
rect 6196 5466 6252 5468
rect 5956 5414 5982 5466
rect 5982 5414 6012 5466
rect 6036 5414 6046 5466
rect 6046 5414 6092 5466
rect 6116 5414 6162 5466
rect 6162 5414 6172 5466
rect 6196 5414 6226 5466
rect 6226 5414 6252 5466
rect 5956 5412 6012 5414
rect 6036 5412 6092 5414
rect 6116 5412 6172 5414
rect 6196 5412 6252 5414
rect 5956 4378 6012 4380
rect 6036 4378 6092 4380
rect 6116 4378 6172 4380
rect 6196 4378 6252 4380
rect 5956 4326 5982 4378
rect 5982 4326 6012 4378
rect 6036 4326 6046 4378
rect 6046 4326 6092 4378
rect 6116 4326 6162 4378
rect 6162 4326 6172 4378
rect 6196 4326 6226 4378
rect 6226 4326 6252 4378
rect 5956 4324 6012 4326
rect 6036 4324 6092 4326
rect 6116 4324 6172 4326
rect 6196 4324 6252 4326
rect 6642 3984 6698 4040
rect 7194 11500 7196 11520
rect 7196 11500 7248 11520
rect 7248 11500 7250 11520
rect 7194 11464 7250 11500
rect 10956 21242 11012 21244
rect 11036 21242 11092 21244
rect 11116 21242 11172 21244
rect 11196 21242 11252 21244
rect 10956 21190 10982 21242
rect 10982 21190 11012 21242
rect 11036 21190 11046 21242
rect 11046 21190 11092 21242
rect 11116 21190 11162 21242
rect 11162 21190 11172 21242
rect 11196 21190 11226 21242
rect 11226 21190 11252 21242
rect 10956 21188 11012 21190
rect 11036 21188 11092 21190
rect 11116 21188 11172 21190
rect 11196 21188 11252 21190
rect 7746 19780 7802 19816
rect 7746 19760 7748 19780
rect 7748 19760 7800 19780
rect 7800 19760 7802 19780
rect 8114 19236 8170 19272
rect 8114 19216 8116 19236
rect 8116 19216 8168 19236
rect 8168 19216 8170 19236
rect 10956 20154 11012 20156
rect 11036 20154 11092 20156
rect 11116 20154 11172 20156
rect 11196 20154 11252 20156
rect 10956 20102 10982 20154
rect 10982 20102 11012 20154
rect 11036 20102 11046 20154
rect 11046 20102 11092 20154
rect 11116 20102 11162 20154
rect 11162 20102 11172 20154
rect 11196 20102 11226 20154
rect 11226 20102 11252 20154
rect 10956 20100 11012 20102
rect 11036 20100 11092 20102
rect 11116 20100 11172 20102
rect 11196 20100 11252 20102
rect 7654 18708 7656 18728
rect 7656 18708 7708 18728
rect 7708 18708 7710 18728
rect 7654 18672 7710 18708
rect 7562 18128 7618 18184
rect 8022 17740 8078 17776
rect 8022 17720 8024 17740
rect 8024 17720 8076 17740
rect 8076 17720 8078 17740
rect 10956 19066 11012 19068
rect 11036 19066 11092 19068
rect 11116 19066 11172 19068
rect 11196 19066 11252 19068
rect 10956 19014 10982 19066
rect 10982 19014 11012 19066
rect 11036 19014 11046 19066
rect 11046 19014 11092 19066
rect 11116 19014 11162 19066
rect 11162 19014 11172 19066
rect 11196 19014 11226 19066
rect 11226 19014 11252 19066
rect 10956 19012 11012 19014
rect 11036 19012 11092 19014
rect 11116 19012 11172 19014
rect 11196 19012 11252 19014
rect 11794 19372 11850 19408
rect 11794 19352 11796 19372
rect 11796 19352 11848 19372
rect 11848 19352 11850 19372
rect 9494 17040 9550 17096
rect 8022 16940 8024 16960
rect 8024 16940 8076 16960
rect 8076 16940 8078 16960
rect 8022 16904 8078 16940
rect 10956 17978 11012 17980
rect 11036 17978 11092 17980
rect 11116 17978 11172 17980
rect 11196 17978 11252 17980
rect 10956 17926 10982 17978
rect 10982 17926 11012 17978
rect 11036 17926 11046 17978
rect 11046 17926 11092 17978
rect 11116 17926 11162 17978
rect 11162 17926 11172 17978
rect 11196 17926 11226 17978
rect 11226 17926 11252 17978
rect 10956 17924 11012 17926
rect 11036 17924 11092 17926
rect 11116 17924 11172 17926
rect 11196 17924 11252 17926
rect 10782 17620 10784 17640
rect 10784 17620 10836 17640
rect 10836 17620 10838 17640
rect 10782 17584 10838 17620
rect 10690 17448 10746 17504
rect 9862 16668 9864 16688
rect 9864 16668 9916 16688
rect 9916 16668 9918 16688
rect 9862 16632 9918 16668
rect 7562 13368 7618 13424
rect 7930 13096 7986 13152
rect 7930 12824 7986 12880
rect 8114 12824 8170 12880
rect 7286 10376 7342 10432
rect 7470 10548 7472 10568
rect 7472 10548 7524 10568
rect 7524 10548 7526 10568
rect 7470 10512 7526 10548
rect 7470 10140 7472 10160
rect 7472 10140 7524 10160
rect 7524 10140 7526 10160
rect 7470 10104 7526 10140
rect 7286 7520 7342 7576
rect 10956 16890 11012 16892
rect 11036 16890 11092 16892
rect 11116 16890 11172 16892
rect 11196 16890 11252 16892
rect 10956 16838 10982 16890
rect 10982 16838 11012 16890
rect 11036 16838 11046 16890
rect 11046 16838 11092 16890
rect 11116 16838 11162 16890
rect 11162 16838 11172 16890
rect 11196 16838 11226 16890
rect 11226 16838 11252 16890
rect 10956 16836 11012 16838
rect 11036 16836 11092 16838
rect 11116 16836 11172 16838
rect 11196 16836 11252 16838
rect 11334 16768 11390 16824
rect 10966 15972 11022 16008
rect 10966 15952 10968 15972
rect 10968 15952 11020 15972
rect 11020 15952 11022 15972
rect 10956 15802 11012 15804
rect 11036 15802 11092 15804
rect 11116 15802 11172 15804
rect 11196 15802 11252 15804
rect 10956 15750 10982 15802
rect 10982 15750 11012 15802
rect 11036 15750 11046 15802
rect 11046 15750 11092 15802
rect 11116 15750 11162 15802
rect 11162 15750 11172 15802
rect 11196 15750 11226 15802
rect 11226 15750 11252 15802
rect 10956 15748 11012 15750
rect 11036 15748 11092 15750
rect 11116 15748 11172 15750
rect 11196 15748 11252 15750
rect 10956 14714 11012 14716
rect 11036 14714 11092 14716
rect 11116 14714 11172 14716
rect 11196 14714 11252 14716
rect 10956 14662 10982 14714
rect 10982 14662 11012 14714
rect 11036 14662 11046 14714
rect 11046 14662 11092 14714
rect 11116 14662 11162 14714
rect 11162 14662 11172 14714
rect 11196 14662 11226 14714
rect 11226 14662 11252 14714
rect 10956 14660 11012 14662
rect 11036 14660 11092 14662
rect 11116 14660 11172 14662
rect 11196 14660 11252 14662
rect 10230 14592 10286 14648
rect 9678 13932 9734 13968
rect 9678 13912 9680 13932
rect 9680 13912 9732 13932
rect 9732 13912 9734 13932
rect 8574 13232 8630 13288
rect 7562 9324 7564 9344
rect 7564 9324 7616 9344
rect 7616 9324 7618 9344
rect 7562 9288 7618 9324
rect 7930 10376 7986 10432
rect 7838 9424 7894 9480
rect 7470 5772 7526 5808
rect 7470 5752 7472 5772
rect 7472 5752 7524 5772
rect 7524 5752 7526 5772
rect 5722 2932 5724 2952
rect 5724 2932 5776 2952
rect 5776 2932 5778 2952
rect 5722 2896 5778 2932
rect 5956 3290 6012 3292
rect 6036 3290 6092 3292
rect 6116 3290 6172 3292
rect 6196 3290 6252 3292
rect 5956 3238 5982 3290
rect 5982 3238 6012 3290
rect 6036 3238 6046 3290
rect 6046 3238 6092 3290
rect 6116 3238 6162 3290
rect 6162 3238 6172 3290
rect 6196 3238 6226 3290
rect 6226 3238 6252 3290
rect 5956 3236 6012 3238
rect 6036 3236 6092 3238
rect 6116 3236 6172 3238
rect 6196 3236 6252 3238
rect 6826 2796 6828 2816
rect 6828 2796 6880 2816
rect 6880 2796 6882 2816
rect 6826 2760 6882 2796
rect 3974 856 4030 912
rect 9678 12588 9680 12608
rect 9680 12588 9732 12608
rect 9732 12588 9734 12608
rect 9678 12552 9734 12588
rect 8850 12280 8906 12336
rect 9678 11464 9734 11520
rect 8574 9696 8630 9752
rect 8574 9560 8630 9616
rect 7746 5364 7802 5400
rect 7746 5344 7748 5364
rect 7748 5344 7800 5364
rect 7800 5344 7802 5364
rect 9402 3576 9458 3632
rect 9218 2896 9274 2952
rect 9402 2896 9458 2952
rect 5956 2202 6012 2204
rect 6036 2202 6092 2204
rect 6116 2202 6172 2204
rect 6196 2202 6252 2204
rect 5956 2150 5982 2202
rect 5982 2150 6012 2202
rect 6036 2150 6046 2202
rect 6046 2150 6092 2202
rect 6116 2150 6162 2202
rect 6162 2150 6172 2202
rect 6196 2150 6226 2202
rect 6226 2150 6252 2202
rect 5956 2148 6012 2150
rect 6036 2148 6092 2150
rect 6116 2148 6172 2150
rect 6196 2148 6252 2150
rect 6366 1400 6422 1456
rect 9954 13776 10010 13832
rect 9862 10412 9864 10432
rect 9864 10412 9916 10432
rect 9916 10412 9918 10432
rect 9862 10376 9918 10412
rect 10138 13268 10140 13288
rect 10140 13268 10192 13288
rect 10192 13268 10194 13288
rect 10138 13232 10194 13268
rect 10046 13096 10102 13152
rect 9862 8880 9918 8936
rect 10506 13504 10562 13560
rect 11334 13912 11390 13968
rect 10956 13626 11012 13628
rect 11036 13626 11092 13628
rect 11116 13626 11172 13628
rect 11196 13626 11252 13628
rect 10956 13574 10982 13626
rect 10982 13574 11012 13626
rect 11036 13574 11046 13626
rect 11046 13574 11092 13626
rect 11116 13574 11162 13626
rect 11162 13574 11172 13626
rect 11196 13574 11226 13626
rect 11226 13574 11252 13626
rect 10956 13572 11012 13574
rect 11036 13572 11092 13574
rect 11116 13572 11172 13574
rect 11196 13572 11252 13574
rect 10322 13096 10378 13152
rect 15956 21786 16012 21788
rect 16036 21786 16092 21788
rect 16116 21786 16172 21788
rect 16196 21786 16252 21788
rect 15956 21734 15982 21786
rect 15982 21734 16012 21786
rect 16036 21734 16046 21786
rect 16046 21734 16092 21786
rect 16116 21734 16162 21786
rect 16162 21734 16172 21786
rect 16196 21734 16226 21786
rect 16226 21734 16252 21786
rect 15956 21732 16012 21734
rect 16036 21732 16092 21734
rect 16116 21732 16172 21734
rect 16196 21732 16252 21734
rect 15956 20698 16012 20700
rect 16036 20698 16092 20700
rect 16116 20698 16172 20700
rect 16196 20698 16252 20700
rect 15956 20646 15982 20698
rect 15982 20646 16012 20698
rect 16036 20646 16046 20698
rect 16046 20646 16092 20698
rect 16116 20646 16162 20698
rect 16162 20646 16172 20698
rect 16196 20646 16226 20698
rect 16226 20646 16252 20698
rect 15956 20644 16012 20646
rect 16036 20644 16092 20646
rect 16116 20644 16172 20646
rect 16196 20644 16252 20646
rect 14922 20440 14978 20496
rect 12346 18808 12402 18864
rect 12162 13524 12218 13560
rect 12162 13504 12164 13524
rect 12164 13504 12216 13524
rect 12216 13504 12218 13524
rect 10322 12824 10378 12880
rect 10506 12824 10562 12880
rect 11334 12824 11390 12880
rect 10782 12552 10838 12608
rect 11334 12552 11390 12608
rect 10956 12538 11012 12540
rect 11036 12538 11092 12540
rect 11116 12538 11172 12540
rect 11196 12538 11252 12540
rect 10956 12486 10982 12538
rect 10982 12486 11012 12538
rect 11036 12486 11046 12538
rect 11046 12486 11092 12538
rect 11116 12486 11162 12538
rect 11162 12486 11172 12538
rect 11196 12486 11226 12538
rect 11226 12486 11252 12538
rect 10956 12484 11012 12486
rect 11036 12484 11092 12486
rect 11116 12484 11172 12486
rect 11196 12484 11252 12486
rect 10956 11450 11012 11452
rect 11036 11450 11092 11452
rect 11116 11450 11172 11452
rect 11196 11450 11252 11452
rect 10956 11398 10982 11450
rect 10982 11398 11012 11450
rect 11036 11398 11046 11450
rect 11046 11398 11092 11450
rect 11116 11398 11162 11450
rect 11162 11398 11172 11450
rect 11196 11398 11226 11450
rect 11226 11398 11252 11450
rect 10956 11396 11012 11398
rect 11036 11396 11092 11398
rect 11116 11396 11172 11398
rect 11196 11396 11252 11398
rect 10598 10648 10654 10704
rect 10956 10362 11012 10364
rect 11036 10362 11092 10364
rect 11116 10362 11172 10364
rect 11196 10362 11252 10364
rect 10956 10310 10982 10362
rect 10982 10310 11012 10362
rect 11036 10310 11046 10362
rect 11046 10310 11092 10362
rect 11116 10310 11162 10362
rect 11162 10310 11172 10362
rect 11196 10310 11226 10362
rect 11226 10310 11252 10362
rect 10956 10308 11012 10310
rect 11036 10308 11092 10310
rect 11116 10308 11172 10310
rect 11196 10308 11252 10310
rect 12530 12144 12586 12200
rect 12162 11192 12218 11248
rect 11978 10376 12034 10432
rect 10322 9424 10378 9480
rect 10956 9274 11012 9276
rect 11036 9274 11092 9276
rect 11116 9274 11172 9276
rect 11196 9274 11252 9276
rect 10956 9222 10982 9274
rect 10982 9222 11012 9274
rect 11036 9222 11046 9274
rect 11046 9222 11092 9274
rect 11116 9222 11162 9274
rect 11162 9222 11172 9274
rect 11196 9222 11226 9274
rect 11226 9222 11252 9274
rect 10956 9220 11012 9222
rect 11036 9220 11092 9222
rect 11116 9220 11172 9222
rect 11196 9220 11252 9222
rect 10956 8186 11012 8188
rect 11036 8186 11092 8188
rect 11116 8186 11172 8188
rect 11196 8186 11252 8188
rect 10956 8134 10982 8186
rect 10982 8134 11012 8186
rect 11036 8134 11046 8186
rect 11046 8134 11092 8186
rect 11116 8134 11162 8186
rect 11162 8134 11172 8186
rect 11196 8134 11226 8186
rect 11226 8134 11252 8186
rect 10956 8132 11012 8134
rect 11036 8132 11092 8134
rect 11116 8132 11172 8134
rect 11196 8132 11252 8134
rect 10956 7098 11012 7100
rect 11036 7098 11092 7100
rect 11116 7098 11172 7100
rect 11196 7098 11252 7100
rect 10956 7046 10982 7098
rect 10982 7046 11012 7098
rect 11036 7046 11046 7098
rect 11046 7046 11092 7098
rect 11116 7046 11162 7098
rect 11162 7046 11172 7098
rect 11196 7046 11226 7098
rect 11226 7046 11252 7098
rect 10956 7044 11012 7046
rect 11036 7044 11092 7046
rect 11116 7044 11172 7046
rect 11196 7044 11252 7046
rect 12162 7148 12164 7168
rect 12164 7148 12216 7168
rect 12216 7148 12218 7168
rect 12162 7112 12218 7148
rect 10322 6840 10378 6896
rect 10956 6010 11012 6012
rect 11036 6010 11092 6012
rect 11116 6010 11172 6012
rect 11196 6010 11252 6012
rect 10956 5958 10982 6010
rect 10982 5958 11012 6010
rect 11036 5958 11046 6010
rect 11046 5958 11092 6010
rect 11116 5958 11162 6010
rect 11162 5958 11172 6010
rect 11196 5958 11226 6010
rect 11226 5958 11252 6010
rect 10956 5956 11012 5958
rect 11036 5956 11092 5958
rect 11116 5956 11172 5958
rect 11196 5956 11252 5958
rect 11794 6704 11850 6760
rect 10966 5616 11022 5672
rect 10956 4922 11012 4924
rect 11036 4922 11092 4924
rect 11116 4922 11172 4924
rect 11196 4922 11252 4924
rect 10956 4870 10982 4922
rect 10982 4870 11012 4922
rect 11036 4870 11046 4922
rect 11046 4870 11092 4922
rect 11116 4870 11162 4922
rect 11162 4870 11172 4922
rect 11196 4870 11226 4922
rect 11226 4870 11252 4922
rect 10956 4868 11012 4870
rect 11036 4868 11092 4870
rect 11116 4868 11172 4870
rect 11196 4868 11252 4870
rect 12346 6840 12402 6896
rect 12714 16088 12770 16144
rect 12714 6160 12770 6216
rect 12162 4664 12218 4720
rect 10046 4120 10102 4176
rect 10956 3834 11012 3836
rect 11036 3834 11092 3836
rect 11116 3834 11172 3836
rect 11196 3834 11252 3836
rect 10956 3782 10982 3834
rect 10982 3782 11012 3834
rect 11036 3782 11046 3834
rect 11046 3782 11092 3834
rect 11116 3782 11162 3834
rect 11162 3782 11172 3834
rect 11196 3782 11226 3834
rect 11226 3782 11252 3834
rect 10956 3780 11012 3782
rect 11036 3780 11092 3782
rect 11116 3780 11172 3782
rect 11196 3780 11252 3782
rect 12530 3440 12586 3496
rect 14554 18808 14610 18864
rect 14554 18264 14610 18320
rect 14738 18284 14794 18320
rect 14738 18264 14740 18284
rect 14740 18264 14792 18284
rect 14792 18264 14794 18284
rect 14830 17584 14886 17640
rect 14830 16788 14886 16824
rect 14830 16768 14832 16788
rect 14832 16768 14884 16788
rect 14884 16768 14886 16788
rect 13634 13388 13690 13424
rect 13634 13368 13636 13388
rect 13636 13368 13688 13388
rect 13688 13368 13690 13388
rect 13634 11756 13690 11792
rect 13634 11736 13636 11756
rect 13636 11736 13688 11756
rect 13688 11736 13690 11756
rect 13450 7268 13506 7304
rect 13450 7248 13452 7268
rect 13452 7248 13504 7268
rect 13504 7248 13506 7268
rect 13358 7148 13360 7168
rect 13360 7148 13412 7168
rect 13412 7148 13414 7168
rect 13358 7112 13414 7148
rect 13450 5072 13506 5128
rect 13542 4936 13598 4992
rect 9862 3032 9918 3088
rect 10956 2746 11012 2748
rect 11036 2746 11092 2748
rect 11116 2746 11172 2748
rect 11196 2746 11252 2748
rect 10956 2694 10982 2746
rect 10982 2694 11012 2746
rect 11036 2694 11046 2746
rect 11046 2694 11092 2746
rect 11116 2694 11162 2746
rect 11162 2694 11172 2746
rect 11196 2694 11226 2746
rect 11226 2694 11252 2746
rect 10956 2692 11012 2694
rect 11036 2692 11092 2694
rect 11116 2692 11172 2694
rect 11196 2692 11252 2694
rect 9770 2488 9826 2544
rect 11058 2508 11114 2544
rect 11058 2488 11060 2508
rect 11060 2488 11112 2508
rect 11112 2488 11114 2508
rect 9954 1400 10010 1456
rect 14922 15952 14978 16008
rect 15956 19610 16012 19612
rect 16036 19610 16092 19612
rect 16116 19610 16172 19612
rect 16196 19610 16252 19612
rect 15956 19558 15982 19610
rect 15982 19558 16012 19610
rect 16036 19558 16046 19610
rect 16046 19558 16092 19610
rect 16116 19558 16162 19610
rect 16162 19558 16172 19610
rect 16196 19558 16226 19610
rect 16226 19558 16252 19610
rect 15956 19556 16012 19558
rect 16036 19556 16092 19558
rect 16116 19556 16172 19558
rect 16196 19556 16252 19558
rect 20956 21242 21012 21244
rect 21036 21242 21092 21244
rect 21116 21242 21172 21244
rect 21196 21242 21252 21244
rect 20956 21190 20982 21242
rect 20982 21190 21012 21242
rect 21036 21190 21046 21242
rect 21046 21190 21092 21242
rect 21116 21190 21162 21242
rect 21162 21190 21172 21242
rect 21196 21190 21226 21242
rect 21226 21190 21252 21242
rect 20956 21188 21012 21190
rect 21036 21188 21092 21190
rect 21116 21188 21172 21190
rect 21196 21188 21252 21190
rect 24858 23024 24914 23080
rect 20626 20476 20628 20496
rect 20628 20476 20680 20496
rect 20680 20476 20682 20496
rect 20626 20440 20682 20476
rect 16670 19760 16726 19816
rect 15956 18522 16012 18524
rect 16036 18522 16092 18524
rect 16116 18522 16172 18524
rect 16196 18522 16252 18524
rect 15956 18470 15982 18522
rect 15982 18470 16012 18522
rect 16036 18470 16046 18522
rect 16046 18470 16092 18522
rect 16116 18470 16162 18522
rect 16162 18470 16172 18522
rect 16196 18470 16226 18522
rect 16226 18470 16252 18522
rect 15956 18468 16012 18470
rect 16036 18468 16092 18470
rect 16116 18468 16172 18470
rect 16196 18468 16252 18470
rect 20956 20154 21012 20156
rect 21036 20154 21092 20156
rect 21116 20154 21172 20156
rect 21196 20154 21252 20156
rect 20956 20102 20982 20154
rect 20982 20102 21012 20154
rect 21036 20102 21046 20154
rect 21046 20102 21092 20154
rect 21116 20102 21162 20154
rect 21162 20102 21172 20154
rect 21196 20102 21226 20154
rect 21226 20102 21252 20154
rect 20956 20100 21012 20102
rect 21036 20100 21092 20102
rect 21116 20100 21172 20102
rect 21196 20100 21252 20102
rect 17314 18808 17370 18864
rect 17038 18420 17094 18456
rect 17038 18400 17040 18420
rect 17040 18400 17092 18420
rect 17092 18400 17094 18420
rect 17130 18264 17186 18320
rect 19338 18672 19394 18728
rect 15750 17484 15752 17504
rect 15752 17484 15804 17504
rect 15804 17484 15806 17504
rect 15750 17448 15806 17484
rect 15956 17434 16012 17436
rect 16036 17434 16092 17436
rect 16116 17434 16172 17436
rect 16196 17434 16252 17436
rect 15956 17382 15982 17434
rect 15982 17382 16012 17434
rect 16036 17382 16046 17434
rect 16046 17382 16092 17434
rect 16116 17382 16162 17434
rect 16162 17382 16172 17434
rect 16196 17382 16226 17434
rect 16226 17382 16252 17434
rect 15956 17380 16012 17382
rect 16036 17380 16092 17382
rect 16116 17380 16172 17382
rect 16196 17380 16252 17382
rect 15750 17176 15806 17232
rect 15658 17040 15714 17096
rect 14922 15408 14978 15464
rect 14922 13932 14978 13968
rect 14922 13912 14924 13932
rect 14924 13912 14976 13932
rect 14976 13912 14978 13932
rect 14002 12824 14058 12880
rect 14646 12588 14648 12608
rect 14648 12588 14700 12608
rect 14700 12588 14702 12608
rect 14646 12552 14702 12588
rect 15198 13096 15254 13152
rect 17774 17720 17830 17776
rect 18234 17604 18290 17640
rect 18234 17584 18236 17604
rect 18236 17584 18288 17604
rect 18288 17584 18290 17604
rect 18510 17176 18566 17232
rect 15956 16346 16012 16348
rect 16036 16346 16092 16348
rect 16116 16346 16172 16348
rect 16196 16346 16252 16348
rect 15956 16294 15982 16346
rect 15982 16294 16012 16346
rect 16036 16294 16046 16346
rect 16046 16294 16092 16346
rect 16116 16294 16162 16346
rect 16162 16294 16172 16346
rect 16196 16294 16226 16346
rect 16226 16294 16252 16346
rect 15956 16292 16012 16294
rect 16036 16292 16092 16294
rect 16116 16292 16172 16294
rect 16196 16292 16252 16294
rect 15106 12280 15162 12336
rect 15474 12416 15530 12472
rect 15474 12144 15530 12200
rect 15474 11192 15530 11248
rect 15382 10512 15438 10568
rect 15658 12144 15714 12200
rect 15658 10648 15714 10704
rect 15382 10240 15438 10296
rect 13910 8608 13966 8664
rect 14646 8880 14702 8936
rect 14370 7520 14426 7576
rect 14922 7148 14924 7168
rect 14924 7148 14976 7168
rect 14976 7148 14978 7168
rect 14922 7112 14978 7148
rect 15198 5208 15254 5264
rect 15658 10376 15714 10432
rect 15658 10124 15714 10160
rect 15658 10104 15660 10124
rect 15660 10104 15712 10124
rect 15712 10104 15714 10124
rect 15658 8880 15714 8936
rect 15566 8472 15622 8528
rect 15474 5616 15530 5672
rect 15956 15258 16012 15260
rect 16036 15258 16092 15260
rect 16116 15258 16172 15260
rect 16196 15258 16252 15260
rect 15956 15206 15982 15258
rect 15982 15206 16012 15258
rect 16036 15206 16046 15258
rect 16046 15206 16092 15258
rect 16116 15206 16162 15258
rect 16162 15206 16172 15258
rect 16196 15206 16226 15258
rect 16226 15206 16252 15258
rect 15956 15204 16012 15206
rect 16036 15204 16092 15206
rect 16116 15204 16172 15206
rect 16196 15204 16252 15206
rect 15956 14170 16012 14172
rect 16036 14170 16092 14172
rect 16116 14170 16172 14172
rect 16196 14170 16252 14172
rect 15956 14118 15982 14170
rect 15982 14118 16012 14170
rect 16036 14118 16046 14170
rect 16046 14118 16092 14170
rect 16116 14118 16162 14170
rect 16162 14118 16172 14170
rect 16196 14118 16226 14170
rect 16226 14118 16252 14170
rect 15956 14116 16012 14118
rect 16036 14116 16092 14118
rect 16116 14116 16172 14118
rect 16196 14116 16252 14118
rect 18602 16632 18658 16688
rect 18418 15408 18474 15464
rect 17958 14592 18014 14648
rect 20166 17720 20222 17776
rect 21638 19916 21694 19952
rect 21638 19896 21640 19916
rect 21640 19896 21692 19916
rect 21692 19896 21694 19916
rect 20956 19066 21012 19068
rect 21036 19066 21092 19068
rect 21116 19066 21172 19068
rect 21196 19066 21252 19068
rect 20956 19014 20982 19066
rect 20982 19014 21012 19066
rect 21036 19014 21046 19066
rect 21046 19014 21092 19066
rect 21116 19014 21162 19066
rect 21162 19014 21172 19066
rect 21196 19014 21226 19066
rect 21226 19014 21252 19066
rect 20956 19012 21012 19014
rect 21036 19012 21092 19014
rect 21116 19012 21172 19014
rect 21196 19012 21252 19014
rect 21178 18808 21234 18864
rect 20956 17978 21012 17980
rect 21036 17978 21092 17980
rect 21116 17978 21172 17980
rect 21196 17978 21252 17980
rect 20956 17926 20982 17978
rect 20982 17926 21012 17978
rect 21036 17926 21046 17978
rect 21046 17926 21092 17978
rect 21116 17926 21162 17978
rect 21162 17926 21172 17978
rect 21196 17926 21226 17978
rect 21226 17926 21252 17978
rect 20956 17924 21012 17926
rect 21036 17924 21092 17926
rect 21116 17924 21172 17926
rect 21196 17924 21252 17926
rect 23662 19896 23718 19952
rect 20956 16890 21012 16892
rect 21036 16890 21092 16892
rect 21116 16890 21172 16892
rect 21196 16890 21252 16892
rect 20956 16838 20982 16890
rect 20982 16838 21012 16890
rect 21036 16838 21046 16890
rect 21046 16838 21092 16890
rect 21116 16838 21162 16890
rect 21162 16838 21172 16890
rect 21196 16838 21226 16890
rect 21226 16838 21252 16890
rect 20956 16836 21012 16838
rect 21036 16836 21092 16838
rect 21116 16836 21172 16838
rect 21196 16836 21252 16838
rect 18694 14864 18750 14920
rect 16670 13912 16726 13968
rect 16854 13912 16910 13968
rect 16854 13368 16910 13424
rect 16302 13232 16358 13288
rect 15956 13082 16012 13084
rect 16036 13082 16092 13084
rect 16116 13082 16172 13084
rect 16196 13082 16252 13084
rect 15956 13030 15982 13082
rect 15982 13030 16012 13082
rect 16036 13030 16046 13082
rect 16046 13030 16092 13082
rect 16116 13030 16162 13082
rect 16162 13030 16172 13082
rect 16196 13030 16226 13082
rect 16226 13030 16252 13082
rect 15956 13028 16012 13030
rect 16036 13028 16092 13030
rect 16116 13028 16172 13030
rect 16196 13028 16252 13030
rect 15956 11994 16012 11996
rect 16036 11994 16092 11996
rect 16116 11994 16172 11996
rect 16196 11994 16252 11996
rect 15956 11942 15982 11994
rect 15982 11942 16012 11994
rect 16036 11942 16046 11994
rect 16046 11942 16092 11994
rect 16116 11942 16162 11994
rect 16162 11942 16172 11994
rect 16196 11942 16226 11994
rect 16226 11942 16252 11994
rect 15956 11940 16012 11942
rect 16036 11940 16092 11942
rect 16116 11940 16172 11942
rect 16196 11940 16252 11942
rect 18694 13912 18750 13968
rect 16394 11192 16450 11248
rect 15956 10906 16012 10908
rect 16036 10906 16092 10908
rect 16116 10906 16172 10908
rect 16196 10906 16252 10908
rect 15956 10854 15982 10906
rect 15982 10854 16012 10906
rect 16036 10854 16046 10906
rect 16046 10854 16092 10906
rect 16116 10854 16162 10906
rect 16162 10854 16172 10906
rect 16196 10854 16226 10906
rect 16226 10854 16252 10906
rect 15956 10852 16012 10854
rect 16036 10852 16092 10854
rect 16116 10852 16172 10854
rect 16196 10852 16252 10854
rect 15842 10240 15898 10296
rect 16486 10784 16542 10840
rect 15956 9818 16012 9820
rect 16036 9818 16092 9820
rect 16116 9818 16172 9820
rect 16196 9818 16252 9820
rect 15956 9766 15982 9818
rect 15982 9766 16012 9818
rect 16036 9766 16046 9818
rect 16046 9766 16092 9818
rect 16116 9766 16162 9818
rect 16162 9766 16172 9818
rect 16196 9766 16226 9818
rect 16226 9766 16252 9818
rect 15956 9764 16012 9766
rect 16036 9764 16092 9766
rect 16116 9764 16172 9766
rect 16196 9764 16252 9766
rect 16762 8916 16764 8936
rect 16764 8916 16816 8936
rect 16816 8916 16818 8936
rect 16762 8880 16818 8916
rect 15956 8730 16012 8732
rect 16036 8730 16092 8732
rect 16116 8730 16172 8732
rect 16196 8730 16252 8732
rect 15956 8678 15982 8730
rect 15982 8678 16012 8730
rect 16036 8678 16046 8730
rect 16046 8678 16092 8730
rect 16116 8678 16162 8730
rect 16162 8678 16172 8730
rect 16196 8678 16226 8730
rect 16226 8678 16252 8730
rect 15956 8676 16012 8678
rect 16036 8676 16092 8678
rect 16116 8676 16172 8678
rect 16196 8676 16252 8678
rect 15956 7642 16012 7644
rect 16036 7642 16092 7644
rect 16116 7642 16172 7644
rect 16196 7642 16252 7644
rect 15956 7590 15982 7642
rect 15982 7590 16012 7642
rect 16036 7590 16046 7642
rect 16046 7590 16092 7642
rect 16116 7590 16162 7642
rect 16162 7590 16172 7642
rect 16196 7590 16226 7642
rect 16226 7590 16252 7642
rect 15956 7588 16012 7590
rect 16036 7588 16092 7590
rect 16116 7588 16172 7590
rect 16196 7588 16252 7590
rect 16118 6740 16120 6760
rect 16120 6740 16172 6760
rect 16172 6740 16174 6760
rect 16118 6704 16174 6740
rect 15956 6554 16012 6556
rect 16036 6554 16092 6556
rect 16116 6554 16172 6556
rect 16196 6554 16252 6556
rect 15956 6502 15982 6554
rect 15982 6502 16012 6554
rect 16036 6502 16046 6554
rect 16046 6502 16092 6554
rect 16116 6502 16162 6554
rect 16162 6502 16172 6554
rect 16196 6502 16226 6554
rect 16226 6502 16252 6554
rect 15956 6500 16012 6502
rect 16036 6500 16092 6502
rect 16116 6500 16172 6502
rect 16196 6500 16252 6502
rect 15842 6296 15898 6352
rect 16670 7384 16726 7440
rect 15566 5072 15622 5128
rect 15956 5466 16012 5468
rect 16036 5466 16092 5468
rect 16116 5466 16172 5468
rect 16196 5466 16252 5468
rect 15956 5414 15982 5466
rect 15982 5414 16012 5466
rect 16036 5414 16046 5466
rect 16046 5414 16092 5466
rect 16116 5414 16162 5466
rect 16162 5414 16172 5466
rect 16196 5414 16226 5466
rect 16226 5414 16252 5466
rect 15956 5412 16012 5414
rect 16036 5412 16092 5414
rect 16116 5412 16172 5414
rect 16196 5412 16252 5414
rect 17958 6060 17960 6080
rect 17960 6060 18012 6080
rect 18012 6060 18014 6080
rect 17958 6024 18014 6060
rect 16486 5480 16542 5536
rect 16670 5344 16726 5400
rect 15956 4378 16012 4380
rect 16036 4378 16092 4380
rect 16116 4378 16172 4380
rect 16196 4378 16252 4380
rect 15956 4326 15982 4378
rect 15982 4326 16012 4378
rect 16036 4326 16046 4378
rect 16046 4326 16092 4378
rect 16116 4326 16162 4378
rect 16162 4326 16172 4378
rect 16196 4326 16226 4378
rect 16226 4326 16252 4378
rect 15956 4324 16012 4326
rect 16036 4324 16092 4326
rect 16116 4324 16172 4326
rect 16196 4324 16252 4326
rect 16670 4392 16726 4448
rect 16394 4120 16450 4176
rect 15956 3290 16012 3292
rect 16036 3290 16092 3292
rect 16116 3290 16172 3292
rect 16196 3290 16252 3292
rect 15956 3238 15982 3290
rect 15982 3238 16012 3290
rect 16036 3238 16046 3290
rect 16046 3238 16092 3290
rect 16116 3238 16162 3290
rect 16162 3238 16172 3290
rect 16196 3238 16226 3290
rect 16226 3238 16252 3290
rect 15956 3236 16012 3238
rect 16036 3236 16092 3238
rect 16116 3236 16172 3238
rect 16196 3236 16252 3238
rect 15956 2202 16012 2204
rect 16036 2202 16092 2204
rect 16116 2202 16172 2204
rect 16196 2202 16252 2204
rect 15956 2150 15982 2202
rect 15982 2150 16012 2202
rect 16036 2150 16046 2202
rect 16046 2150 16092 2202
rect 16116 2150 16162 2202
rect 16162 2150 16172 2202
rect 16196 2150 16226 2202
rect 16226 2150 16252 2202
rect 15956 2148 16012 2150
rect 16036 2148 16092 2150
rect 16116 2148 16172 2150
rect 16196 2148 16252 2150
rect 18142 12552 18198 12608
rect 20956 15802 21012 15804
rect 21036 15802 21092 15804
rect 21116 15802 21172 15804
rect 21196 15802 21252 15804
rect 20956 15750 20982 15802
rect 20982 15750 21012 15802
rect 21036 15750 21046 15802
rect 21046 15750 21092 15802
rect 21116 15750 21162 15802
rect 21162 15750 21172 15802
rect 21196 15750 21226 15802
rect 21226 15750 21252 15802
rect 20956 15748 21012 15750
rect 21036 15748 21092 15750
rect 21116 15748 21172 15750
rect 21196 15748 21252 15750
rect 20956 14714 21012 14716
rect 21036 14714 21092 14716
rect 21116 14714 21172 14716
rect 21196 14714 21252 14716
rect 20956 14662 20982 14714
rect 20982 14662 21012 14714
rect 21036 14662 21046 14714
rect 21046 14662 21092 14714
rect 21116 14662 21162 14714
rect 21162 14662 21172 14714
rect 21196 14662 21226 14714
rect 21226 14662 21252 14714
rect 20956 14660 21012 14662
rect 21036 14660 21092 14662
rect 21116 14660 21172 14662
rect 21196 14660 21252 14662
rect 19890 14612 19946 14648
rect 19890 14592 19892 14612
rect 19892 14592 19944 14612
rect 19944 14592 19946 14612
rect 20718 13912 20774 13968
rect 18510 7384 18566 7440
rect 18418 7248 18474 7304
rect 18510 6432 18566 6488
rect 19246 12688 19302 12744
rect 19154 12588 19156 12608
rect 19156 12588 19208 12608
rect 19208 12588 19210 12608
rect 19154 12552 19210 12588
rect 20956 13626 21012 13628
rect 21036 13626 21092 13628
rect 21116 13626 21172 13628
rect 21196 13626 21252 13628
rect 20956 13574 20982 13626
rect 20982 13574 21012 13626
rect 21036 13574 21046 13626
rect 21046 13574 21092 13626
rect 21116 13574 21162 13626
rect 21162 13574 21172 13626
rect 21196 13574 21226 13626
rect 21226 13574 21252 13626
rect 20956 13572 21012 13574
rect 21036 13572 21092 13574
rect 21116 13572 21172 13574
rect 21196 13572 21252 13574
rect 20718 12960 20774 13016
rect 20534 12280 20590 12336
rect 21730 12708 21786 12744
rect 21730 12688 21732 12708
rect 21732 12688 21784 12708
rect 21784 12688 21786 12708
rect 20718 12552 20774 12608
rect 19062 10648 19118 10704
rect 19522 10920 19578 10976
rect 19062 10260 19118 10296
rect 19062 10240 19064 10260
rect 19064 10240 19116 10260
rect 19116 10240 19118 10260
rect 19154 9968 19210 10024
rect 19154 9560 19210 9616
rect 19338 9424 19394 9480
rect 19246 8780 19248 8800
rect 19248 8780 19300 8800
rect 19300 8780 19302 8800
rect 19246 8744 19302 8780
rect 19062 7928 19118 7984
rect 18786 3168 18842 3224
rect 19062 7112 19118 7168
rect 19522 5752 19578 5808
rect 20956 12538 21012 12540
rect 21036 12538 21092 12540
rect 21116 12538 21172 12540
rect 21196 12538 21252 12540
rect 20956 12486 20982 12538
rect 20982 12486 21012 12538
rect 21036 12486 21046 12538
rect 21046 12486 21092 12538
rect 21116 12486 21162 12538
rect 21162 12486 21172 12538
rect 21196 12486 21226 12538
rect 21226 12486 21252 12538
rect 20956 12484 21012 12486
rect 21036 12484 21092 12486
rect 21116 12484 21172 12486
rect 21196 12484 21252 12486
rect 21730 12416 21786 12472
rect 21270 11636 21272 11656
rect 21272 11636 21324 11656
rect 21324 11636 21326 11656
rect 21270 11600 21326 11636
rect 20956 11450 21012 11452
rect 21036 11450 21092 11452
rect 21116 11450 21172 11452
rect 21196 11450 21252 11452
rect 20956 11398 20982 11450
rect 20982 11398 21012 11450
rect 21036 11398 21046 11450
rect 21046 11398 21092 11450
rect 21116 11398 21162 11450
rect 21162 11398 21172 11450
rect 21196 11398 21226 11450
rect 21226 11398 21252 11450
rect 20956 11396 21012 11398
rect 21036 11396 21092 11398
rect 21116 11396 21172 11398
rect 21196 11396 21252 11398
rect 21730 11056 21786 11112
rect 21454 10784 21510 10840
rect 20956 10362 21012 10364
rect 21036 10362 21092 10364
rect 21116 10362 21172 10364
rect 21196 10362 21252 10364
rect 20956 10310 20982 10362
rect 20982 10310 21012 10362
rect 21036 10310 21046 10362
rect 21046 10310 21092 10362
rect 21116 10310 21162 10362
rect 21162 10310 21172 10362
rect 21196 10310 21226 10362
rect 21226 10310 21252 10362
rect 20956 10308 21012 10310
rect 21036 10308 21092 10310
rect 21116 10308 21172 10310
rect 21196 10308 21252 10310
rect 21362 10240 21418 10296
rect 21546 9968 21602 10024
rect 20956 9274 21012 9276
rect 21036 9274 21092 9276
rect 21116 9274 21172 9276
rect 21196 9274 21252 9276
rect 20956 9222 20982 9274
rect 20982 9222 21012 9274
rect 21036 9222 21046 9274
rect 21046 9222 21092 9274
rect 21116 9222 21162 9274
rect 21162 9222 21172 9274
rect 21196 9222 21226 9274
rect 21226 9222 21252 9274
rect 20956 9220 21012 9222
rect 21036 9220 21092 9222
rect 21116 9220 21172 9222
rect 21196 9220 21252 9222
rect 20718 8744 20774 8800
rect 21362 8744 21418 8800
rect 20534 5752 20590 5808
rect 20350 5228 20406 5264
rect 20350 5208 20352 5228
rect 20352 5208 20404 5228
rect 20404 5208 20406 5228
rect 19246 4120 19302 4176
rect 19890 4564 19892 4584
rect 19892 4564 19944 4584
rect 19944 4564 19946 4584
rect 19890 4528 19946 4564
rect 19982 3168 20038 3224
rect 19154 2760 19210 2816
rect 20956 8186 21012 8188
rect 21036 8186 21092 8188
rect 21116 8186 21172 8188
rect 21196 8186 21252 8188
rect 20956 8134 20982 8186
rect 20982 8134 21012 8186
rect 21036 8134 21046 8186
rect 21046 8134 21092 8186
rect 21116 8134 21162 8186
rect 21162 8134 21172 8186
rect 21196 8134 21226 8186
rect 21226 8134 21252 8186
rect 20956 8132 21012 8134
rect 21036 8132 21092 8134
rect 21116 8132 21172 8134
rect 21196 8132 21252 8134
rect 20956 7098 21012 7100
rect 21036 7098 21092 7100
rect 21116 7098 21172 7100
rect 21196 7098 21252 7100
rect 20956 7046 20982 7098
rect 20982 7046 21012 7098
rect 21036 7046 21046 7098
rect 21046 7046 21092 7098
rect 21116 7046 21162 7098
rect 21162 7046 21172 7098
rect 21196 7046 21226 7098
rect 21226 7046 21252 7098
rect 20956 7044 21012 7046
rect 21036 7044 21092 7046
rect 21116 7044 21172 7046
rect 21196 7044 21252 7046
rect 20956 6010 21012 6012
rect 21036 6010 21092 6012
rect 21116 6010 21172 6012
rect 21196 6010 21252 6012
rect 20956 5958 20982 6010
rect 20982 5958 21012 6010
rect 21036 5958 21046 6010
rect 21046 5958 21092 6010
rect 21116 5958 21162 6010
rect 21162 5958 21172 6010
rect 21196 5958 21226 6010
rect 21226 5958 21252 6010
rect 20956 5956 21012 5958
rect 21036 5956 21092 5958
rect 21116 5956 21172 5958
rect 21196 5956 21252 5958
rect 20956 4922 21012 4924
rect 21036 4922 21092 4924
rect 21116 4922 21172 4924
rect 21196 4922 21252 4924
rect 20956 4870 20982 4922
rect 20982 4870 21012 4922
rect 21036 4870 21046 4922
rect 21046 4870 21092 4922
rect 21116 4870 21162 4922
rect 21162 4870 21172 4922
rect 21196 4870 21226 4922
rect 21226 4870 21252 4922
rect 20956 4868 21012 4870
rect 21036 4868 21092 4870
rect 21116 4868 21172 4870
rect 21196 4868 21252 4870
rect 20718 4392 20774 4448
rect 21822 9560 21878 9616
rect 24122 19216 24178 19272
rect 23570 18164 23572 18184
rect 23572 18164 23624 18184
rect 23624 18164 23626 18184
rect 23570 18128 23626 18164
rect 23478 17176 23534 17232
rect 23110 16088 23166 16144
rect 23478 14864 23534 14920
rect 22558 13912 22614 13968
rect 22098 12824 22154 12880
rect 23478 12416 23534 12472
rect 22006 11736 22062 11792
rect 22558 9580 22614 9616
rect 22558 9560 22560 9580
rect 22560 9560 22612 9580
rect 22612 9560 22614 9580
rect 21914 8508 21916 8528
rect 21916 8508 21968 8528
rect 21968 8508 21970 8528
rect 21914 8472 21970 8508
rect 23846 16632 23902 16688
rect 24030 17856 24086 17912
rect 23754 15408 23810 15464
rect 23570 9968 23626 10024
rect 20626 3984 20682 4040
rect 20956 3834 21012 3836
rect 21036 3834 21092 3836
rect 21116 3834 21172 3836
rect 21196 3834 21252 3836
rect 20956 3782 20982 3834
rect 20982 3782 21012 3834
rect 21036 3782 21046 3834
rect 21046 3782 21092 3834
rect 21116 3782 21162 3834
rect 21162 3782 21172 3834
rect 21196 3782 21226 3834
rect 21226 3782 21252 3834
rect 20956 3780 21012 3782
rect 21036 3780 21092 3782
rect 21116 3780 21172 3782
rect 21196 3780 21252 3782
rect 20626 2760 20682 2816
rect 22006 5616 22062 5672
rect 22006 5072 22062 5128
rect 22006 3848 22062 3904
rect 20956 2746 21012 2748
rect 21036 2746 21092 2748
rect 21116 2746 21172 2748
rect 21196 2746 21252 2748
rect 20956 2694 20982 2746
rect 20982 2694 21012 2746
rect 21036 2694 21046 2746
rect 21046 2694 21092 2746
rect 21116 2694 21162 2746
rect 21162 2694 21172 2746
rect 21196 2694 21226 2746
rect 21226 2694 21252 2746
rect 20956 2692 21012 2694
rect 21036 2692 21092 2694
rect 21116 2692 21172 2694
rect 21196 2692 21252 2694
rect 24858 19252 24860 19272
rect 24860 19252 24912 19272
rect 24912 19252 24914 19272
rect 24858 19216 24914 19252
rect 24214 18400 24270 18456
rect 24306 17584 24362 17640
rect 24490 15408 24546 15464
rect 24398 14592 24454 14648
rect 24214 10240 24270 10296
rect 24766 13368 24822 13424
rect 25134 21256 25190 21312
rect 25226 20032 25282 20088
rect 25134 18672 25190 18728
rect 25134 18300 25136 18320
rect 25136 18300 25188 18320
rect 25188 18300 25190 18320
rect 25134 18264 25190 18300
rect 25318 19352 25374 19408
rect 25318 18400 25374 18456
rect 25318 17584 25374 17640
rect 25594 22344 25650 22400
rect 25956 21786 26012 21788
rect 26036 21786 26092 21788
rect 26116 21786 26172 21788
rect 26196 21786 26252 21788
rect 25956 21734 25982 21786
rect 25982 21734 26012 21786
rect 26036 21734 26046 21786
rect 26046 21734 26092 21786
rect 26116 21734 26162 21786
rect 26162 21734 26172 21786
rect 26196 21734 26226 21786
rect 26226 21734 26252 21786
rect 25956 21732 26012 21734
rect 26036 21732 26092 21734
rect 26116 21732 26172 21734
rect 26196 21732 26252 21734
rect 25870 21528 25926 21584
rect 25778 20440 25834 20496
rect 25502 16088 25558 16144
rect 25042 14864 25098 14920
rect 25042 12960 25098 13016
rect 25134 12552 25190 12608
rect 25042 12144 25098 12200
rect 25226 12144 25282 12200
rect 25042 12008 25098 12064
rect 24950 10920 25006 10976
rect 24122 9016 24178 9072
rect 23846 6160 23902 6216
rect 23754 5616 23810 5672
rect 23938 5480 23994 5536
rect 23938 5072 23994 5128
rect 23846 4020 23848 4040
rect 23848 4020 23900 4040
rect 23900 4020 23902 4040
rect 23846 3984 23902 4020
rect 23846 2896 23902 2952
rect 24214 7420 24216 7440
rect 24216 7420 24268 7440
rect 24268 7420 24270 7440
rect 24214 7384 24270 7420
rect 24122 6432 24178 6488
rect 25226 11464 25282 11520
rect 25226 7928 25282 7984
rect 24766 5344 24822 5400
rect 24950 4548 25006 4584
rect 24950 4528 24952 4548
rect 24952 4528 25004 4548
rect 25004 4528 25006 4548
rect 24858 3712 24914 3768
rect 22006 1400 22062 1456
rect 24214 1400 24270 1456
rect 25502 11328 25558 11384
rect 25956 20698 26012 20700
rect 26036 20698 26092 20700
rect 26116 20698 26172 20700
rect 26196 20698 26252 20700
rect 25956 20646 25982 20698
rect 25982 20646 26012 20698
rect 26036 20646 26046 20698
rect 26046 20646 26092 20698
rect 26116 20646 26162 20698
rect 26162 20646 26172 20698
rect 26196 20646 26226 20698
rect 26226 20646 26252 20698
rect 25956 20644 26012 20646
rect 26036 20644 26092 20646
rect 26116 20644 26172 20646
rect 26196 20644 26252 20646
rect 26330 20304 26386 20360
rect 25956 19610 26012 19612
rect 26036 19610 26092 19612
rect 26116 19610 26172 19612
rect 26196 19610 26252 19612
rect 25956 19558 25982 19610
rect 25982 19558 26012 19610
rect 26036 19558 26046 19610
rect 26046 19558 26092 19610
rect 26116 19558 26162 19610
rect 26162 19558 26172 19610
rect 26196 19558 26226 19610
rect 26226 19558 26252 19610
rect 25956 19556 26012 19558
rect 26036 19556 26092 19558
rect 26116 19556 26172 19558
rect 26196 19556 26252 19558
rect 25956 18522 26012 18524
rect 26036 18522 26092 18524
rect 26116 18522 26172 18524
rect 26196 18522 26252 18524
rect 25956 18470 25982 18522
rect 25982 18470 26012 18522
rect 26036 18470 26046 18522
rect 26046 18470 26092 18522
rect 26116 18470 26162 18522
rect 26162 18470 26172 18522
rect 26196 18470 26226 18522
rect 26226 18470 26252 18522
rect 25956 18468 26012 18470
rect 26036 18468 26092 18470
rect 26116 18468 26172 18470
rect 26196 18468 26252 18470
rect 26514 17856 26570 17912
rect 26422 17720 26478 17776
rect 25956 17434 26012 17436
rect 26036 17434 26092 17436
rect 26116 17434 26172 17436
rect 26196 17434 26252 17436
rect 25956 17382 25982 17434
rect 25982 17382 26012 17434
rect 26036 17382 26046 17434
rect 26046 17382 26092 17434
rect 26116 17382 26162 17434
rect 26162 17382 26172 17434
rect 26196 17382 26226 17434
rect 26226 17382 26252 17434
rect 25956 17380 26012 17382
rect 26036 17380 26092 17382
rect 26116 17380 26172 17382
rect 26196 17380 26252 17382
rect 25778 15544 25834 15600
rect 25778 15408 25834 15464
rect 25778 13776 25834 13832
rect 25778 13640 25834 13696
rect 25778 12552 25834 12608
rect 25778 11736 25834 11792
rect 25502 6840 25558 6896
rect 25956 16346 26012 16348
rect 26036 16346 26092 16348
rect 26116 16346 26172 16348
rect 26196 16346 26252 16348
rect 25956 16294 25982 16346
rect 25982 16294 26012 16346
rect 26036 16294 26046 16346
rect 26046 16294 26092 16346
rect 26116 16294 26162 16346
rect 26162 16294 26172 16346
rect 26196 16294 26226 16346
rect 26226 16294 26252 16346
rect 25956 16292 26012 16294
rect 26036 16292 26092 16294
rect 26116 16292 26172 16294
rect 26196 16292 26252 16294
rect 25956 15258 26012 15260
rect 26036 15258 26092 15260
rect 26116 15258 26172 15260
rect 26196 15258 26252 15260
rect 25956 15206 25982 15258
rect 25982 15206 26012 15258
rect 26036 15206 26046 15258
rect 26046 15206 26092 15258
rect 26116 15206 26162 15258
rect 26162 15206 26172 15258
rect 26196 15206 26226 15258
rect 26226 15206 26252 15258
rect 25956 15204 26012 15206
rect 26036 15204 26092 15206
rect 26116 15204 26172 15206
rect 26196 15204 26252 15206
rect 25956 14170 26012 14172
rect 26036 14170 26092 14172
rect 26116 14170 26172 14172
rect 26196 14170 26252 14172
rect 25956 14118 25982 14170
rect 25982 14118 26012 14170
rect 26036 14118 26046 14170
rect 26046 14118 26092 14170
rect 26116 14118 26162 14170
rect 26162 14118 26172 14170
rect 26196 14118 26226 14170
rect 26226 14118 26252 14170
rect 25956 14116 26012 14118
rect 26036 14116 26092 14118
rect 26116 14116 26172 14118
rect 26196 14116 26252 14118
rect 26146 13912 26202 13968
rect 25956 13082 26012 13084
rect 26036 13082 26092 13084
rect 26116 13082 26172 13084
rect 26196 13082 26252 13084
rect 25956 13030 25982 13082
rect 25982 13030 26012 13082
rect 26036 13030 26046 13082
rect 26046 13030 26092 13082
rect 26116 13030 26162 13082
rect 26162 13030 26172 13082
rect 26196 13030 26226 13082
rect 26226 13030 26252 13082
rect 25956 13028 26012 13030
rect 26036 13028 26092 13030
rect 26116 13028 26172 13030
rect 26196 13028 26252 13030
rect 25956 11994 26012 11996
rect 26036 11994 26092 11996
rect 26116 11994 26172 11996
rect 26196 11994 26252 11996
rect 25956 11942 25982 11994
rect 25982 11942 26012 11994
rect 26036 11942 26046 11994
rect 26046 11942 26092 11994
rect 26116 11942 26162 11994
rect 26162 11942 26172 11994
rect 26196 11942 26226 11994
rect 26226 11942 26252 11994
rect 25956 11940 26012 11942
rect 26036 11940 26092 11942
rect 26116 11940 26172 11942
rect 26196 11940 26252 11942
rect 26698 11600 26754 11656
rect 25870 11056 25926 11112
rect 25956 10906 26012 10908
rect 26036 10906 26092 10908
rect 26116 10906 26172 10908
rect 26196 10906 26252 10908
rect 25956 10854 25982 10906
rect 25982 10854 26012 10906
rect 26036 10854 26046 10906
rect 26046 10854 26092 10906
rect 26116 10854 26162 10906
rect 26162 10854 26172 10906
rect 26196 10854 26226 10906
rect 26226 10854 26252 10906
rect 25956 10852 26012 10854
rect 26036 10852 26092 10854
rect 26116 10852 26172 10854
rect 26196 10852 26252 10854
rect 26606 10412 26608 10432
rect 26608 10412 26660 10432
rect 26660 10412 26662 10432
rect 26606 10376 26662 10412
rect 26514 10104 26570 10160
rect 26422 9968 26478 10024
rect 25956 9818 26012 9820
rect 26036 9818 26092 9820
rect 26116 9818 26172 9820
rect 26196 9818 26252 9820
rect 25956 9766 25982 9818
rect 25982 9766 26012 9818
rect 26036 9766 26046 9818
rect 26046 9766 26092 9818
rect 26116 9766 26162 9818
rect 26162 9766 26172 9818
rect 26196 9766 26226 9818
rect 26226 9766 26252 9818
rect 25956 9764 26012 9766
rect 26036 9764 26092 9766
rect 26116 9764 26172 9766
rect 26196 9764 26252 9766
rect 26698 9868 26700 9888
rect 26700 9868 26752 9888
rect 26752 9868 26754 9888
rect 26698 9832 26754 9868
rect 26698 9288 26754 9344
rect 25956 8730 26012 8732
rect 26036 8730 26092 8732
rect 26116 8730 26172 8732
rect 26196 8730 26252 8732
rect 25956 8678 25982 8730
rect 25982 8678 26012 8730
rect 26036 8678 26046 8730
rect 26046 8678 26092 8730
rect 26116 8678 26162 8730
rect 26162 8678 26172 8730
rect 26196 8678 26226 8730
rect 26226 8678 26252 8730
rect 25956 8676 26012 8678
rect 26036 8676 26092 8678
rect 26116 8676 26172 8678
rect 26196 8676 26252 8678
rect 26698 8608 26754 8664
rect 25956 7642 26012 7644
rect 26036 7642 26092 7644
rect 26116 7642 26172 7644
rect 26196 7642 26252 7644
rect 25956 7590 25982 7642
rect 25982 7590 26012 7642
rect 26036 7590 26046 7642
rect 26046 7590 26092 7642
rect 26116 7590 26162 7642
rect 26162 7590 26172 7642
rect 26196 7590 26226 7642
rect 26226 7590 26252 7642
rect 25956 7588 26012 7590
rect 26036 7588 26092 7590
rect 26116 7588 26172 7590
rect 26196 7588 26252 7590
rect 26330 7384 26386 7440
rect 25962 7284 25964 7304
rect 25964 7284 26016 7304
rect 26016 7284 26018 7304
rect 25962 7248 26018 7284
rect 25956 6554 26012 6556
rect 26036 6554 26092 6556
rect 26116 6554 26172 6556
rect 26196 6554 26252 6556
rect 25956 6502 25982 6554
rect 25982 6502 26012 6554
rect 26036 6502 26046 6554
rect 26046 6502 26092 6554
rect 26116 6502 26162 6554
rect 26162 6502 26172 6554
rect 26196 6502 26226 6554
rect 26226 6502 26252 6554
rect 25956 6500 26012 6502
rect 26036 6500 26092 6502
rect 26116 6500 26172 6502
rect 26196 6500 26252 6502
rect 26238 6316 26294 6352
rect 26238 6296 26240 6316
rect 26240 6296 26292 6316
rect 26292 6296 26294 6316
rect 25778 6160 25834 6216
rect 25956 5466 26012 5468
rect 26036 5466 26092 5468
rect 26116 5466 26172 5468
rect 26196 5466 26252 5468
rect 25956 5414 25982 5466
rect 25982 5414 26012 5466
rect 26036 5414 26046 5466
rect 26046 5414 26092 5466
rect 26116 5414 26162 5466
rect 26162 5414 26172 5466
rect 26196 5414 26226 5466
rect 26226 5414 26252 5466
rect 25956 5412 26012 5414
rect 26036 5412 26092 5414
rect 26116 5412 26172 5414
rect 26196 5412 26252 5414
rect 25956 4378 26012 4380
rect 26036 4378 26092 4380
rect 26116 4378 26172 4380
rect 26196 4378 26252 4380
rect 25956 4326 25982 4378
rect 25982 4326 26012 4378
rect 26036 4326 26046 4378
rect 26046 4326 26092 4378
rect 26116 4326 26162 4378
rect 26162 4326 26172 4378
rect 26196 4326 26226 4378
rect 26226 4326 26252 4378
rect 25956 4324 26012 4326
rect 26036 4324 26092 4326
rect 26116 4324 26172 4326
rect 26196 4324 26252 4326
rect 26698 7384 26754 7440
rect 26514 5772 26570 5808
rect 26514 5752 26516 5772
rect 26516 5752 26568 5772
rect 26568 5752 26570 5772
rect 26606 5616 26662 5672
rect 26422 5208 26478 5264
rect 26514 5072 26570 5128
rect 26698 5072 26754 5128
rect 26698 4120 26754 4176
rect 26974 18808 27030 18864
rect 26974 13504 27030 13560
rect 27434 15816 27490 15872
rect 27342 12280 27398 12336
rect 27618 12144 27674 12200
rect 27526 10648 27582 10704
rect 26974 9596 26976 9616
rect 26976 9596 27028 9616
rect 27028 9596 27030 9616
rect 26974 9560 27030 9596
rect 26882 3984 26938 4040
rect 26606 3848 26662 3904
rect 25502 3460 25558 3496
rect 25502 3440 25504 3460
rect 25504 3440 25556 3460
rect 25556 3440 25558 3460
rect 27710 8064 27766 8120
rect 27066 3712 27122 3768
rect 25956 3290 26012 3292
rect 26036 3290 26092 3292
rect 26116 3290 26172 3292
rect 26196 3290 26252 3292
rect 25956 3238 25982 3290
rect 25982 3238 26012 3290
rect 26036 3238 26046 3290
rect 26046 3238 26092 3290
rect 26116 3238 26162 3290
rect 26162 3238 26172 3290
rect 26196 3238 26226 3290
rect 26226 3238 26252 3290
rect 25956 3236 26012 3238
rect 26036 3236 26092 3238
rect 26116 3236 26172 3238
rect 26196 3236 26252 3238
rect 25318 3052 25374 3088
rect 25318 3032 25320 3052
rect 25320 3032 25372 3052
rect 25372 3032 25374 3052
rect 25956 2202 26012 2204
rect 26036 2202 26092 2204
rect 26116 2202 26172 2204
rect 26196 2202 26252 2204
rect 25956 2150 25982 2202
rect 25982 2150 26012 2202
rect 26036 2150 26046 2202
rect 26046 2150 26092 2202
rect 26116 2150 26162 2202
rect 26162 2150 26172 2202
rect 26196 2150 26226 2202
rect 26226 2150 26252 2202
rect 25956 2148 26012 2150
rect 26036 2148 26092 2150
rect 26116 2148 26172 2150
rect 26196 2148 26252 2150
rect 25870 1400 25926 1456
rect 26422 3032 26478 3088
rect 26698 2080 26754 2136
rect 26606 856 26662 912
rect 1398 312 1454 368
rect 27526 4392 27582 4448
rect 27618 3984 27674 4040
rect 27710 2796 27712 2816
rect 27712 2796 27764 2816
rect 27764 2796 27766 2816
rect 27710 2760 27766 2796
rect 26790 312 26846 368
<< metal3 >>
rect 0 23626 480 23656
rect 3325 23626 3391 23629
rect 0 23624 3391 23626
rect 0 23568 3330 23624
rect 3386 23568 3391 23624
rect 0 23566 3391 23568
rect 0 23536 480 23566
rect 3325 23563 3391 23566
rect 25405 23626 25471 23629
rect 29520 23626 30000 23656
rect 25405 23624 30000 23626
rect 25405 23568 25410 23624
rect 25466 23568 30000 23624
rect 25405 23566 30000 23568
rect 25405 23563 25471 23566
rect 29520 23536 30000 23566
rect 0 23082 480 23112
rect 4153 23082 4219 23085
rect 0 23080 4219 23082
rect 0 23024 4158 23080
rect 4214 23024 4219 23080
rect 0 23022 4219 23024
rect 0 22992 480 23022
rect 4153 23019 4219 23022
rect 24853 23082 24919 23085
rect 29520 23082 30000 23112
rect 24853 23080 30000 23082
rect 24853 23024 24858 23080
rect 24914 23024 30000 23080
rect 24853 23022 30000 23024
rect 24853 23019 24919 23022
rect 29520 22992 30000 23022
rect 0 22402 480 22432
rect 2773 22402 2839 22405
rect 0 22400 2839 22402
rect 0 22344 2778 22400
rect 2834 22344 2839 22400
rect 0 22342 2839 22344
rect 0 22312 480 22342
rect 2773 22339 2839 22342
rect 25589 22402 25655 22405
rect 29520 22402 30000 22432
rect 25589 22400 30000 22402
rect 25589 22344 25594 22400
rect 25650 22344 30000 22400
rect 25589 22342 30000 22344
rect 25589 22339 25655 22342
rect 29520 22312 30000 22342
rect 0 21858 480 21888
rect 4061 21858 4127 21861
rect 29520 21858 30000 21888
rect 0 21856 4127 21858
rect 0 21800 4066 21856
rect 4122 21800 4127 21856
rect 0 21798 4127 21800
rect 0 21768 480 21798
rect 4061 21795 4127 21798
rect 26374 21798 30000 21858
rect 5944 21792 6264 21793
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 21727 6264 21728
rect 15944 21792 16264 21793
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 21727 16264 21728
rect 25944 21792 26264 21793
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 21727 26264 21728
rect 25865 21586 25931 21589
rect 26374 21586 26434 21798
rect 29520 21768 30000 21798
rect 25865 21584 26434 21586
rect 25865 21528 25870 21584
rect 25926 21528 26434 21584
rect 25865 21526 26434 21528
rect 25865 21523 25931 21526
rect 0 21314 480 21344
rect 3969 21314 4035 21317
rect 0 21312 4035 21314
rect 0 21256 3974 21312
rect 4030 21256 4035 21312
rect 0 21254 4035 21256
rect 0 21224 480 21254
rect 3969 21251 4035 21254
rect 25129 21314 25195 21317
rect 29520 21314 30000 21344
rect 25129 21312 30000 21314
rect 25129 21256 25134 21312
rect 25190 21256 30000 21312
rect 25129 21254 30000 21256
rect 25129 21251 25195 21254
rect 10944 21248 11264 21249
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 21183 11264 21184
rect 20944 21248 21264 21249
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 29520 21224 30000 21254
rect 20944 21183 21264 21184
rect 5944 20704 6264 20705
rect 0 20634 480 20664
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 20639 6264 20640
rect 15944 20704 16264 20705
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 20639 16264 20640
rect 25944 20704 26264 20705
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 20639 26264 20640
rect 3785 20634 3851 20637
rect 29520 20634 30000 20664
rect 0 20632 3851 20634
rect 0 20576 3790 20632
rect 3846 20576 3851 20632
rect 0 20574 3851 20576
rect 0 20544 480 20574
rect 3785 20571 3851 20574
rect 26374 20574 30000 20634
rect 14917 20498 14983 20501
rect 20621 20498 20687 20501
rect 14917 20496 20687 20498
rect 14917 20440 14922 20496
rect 14978 20440 20626 20496
rect 20682 20440 20687 20496
rect 14917 20438 20687 20440
rect 14917 20435 14983 20438
rect 20621 20435 20687 20438
rect 25773 20498 25839 20501
rect 26374 20498 26434 20574
rect 29520 20544 30000 20574
rect 25773 20496 26434 20498
rect 25773 20440 25778 20496
rect 25834 20440 26434 20496
rect 25773 20438 26434 20440
rect 25773 20435 25839 20438
rect 4981 20362 5047 20365
rect 26325 20362 26391 20365
rect 4981 20360 26391 20362
rect 4981 20304 4986 20360
rect 5042 20304 26330 20360
rect 26386 20304 26391 20360
rect 4981 20302 26391 20304
rect 4981 20299 5047 20302
rect 26325 20299 26391 20302
rect 10944 20160 11264 20161
rect 0 20090 480 20120
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 20095 11264 20096
rect 20944 20160 21264 20161
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 20095 21264 20096
rect 3325 20090 3391 20093
rect 0 20088 3391 20090
rect 0 20032 3330 20088
rect 3386 20032 3391 20088
rect 0 20030 3391 20032
rect 0 20000 480 20030
rect 3325 20027 3391 20030
rect 4061 20090 4127 20093
rect 6637 20090 6703 20093
rect 4061 20088 6703 20090
rect 4061 20032 4066 20088
rect 4122 20032 6642 20088
rect 6698 20032 6703 20088
rect 4061 20030 6703 20032
rect 4061 20027 4127 20030
rect 6637 20027 6703 20030
rect 25221 20090 25287 20093
rect 29520 20090 30000 20120
rect 25221 20088 30000 20090
rect 25221 20032 25226 20088
rect 25282 20032 30000 20088
rect 25221 20030 30000 20032
rect 25221 20027 25287 20030
rect 29520 20000 30000 20030
rect 21633 19954 21699 19957
rect 23657 19954 23723 19957
rect 21633 19952 23723 19954
rect 21633 19896 21638 19952
rect 21694 19896 23662 19952
rect 23718 19896 23723 19952
rect 21633 19894 23723 19896
rect 21633 19891 21699 19894
rect 23657 19891 23723 19894
rect 7741 19818 7807 19821
rect 16665 19818 16731 19821
rect 7741 19816 16731 19818
rect 7741 19760 7746 19816
rect 7802 19760 16670 19816
rect 16726 19760 16731 19816
rect 7741 19758 16731 19760
rect 7741 19755 7807 19758
rect 16665 19755 16731 19758
rect 5944 19616 6264 19617
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 19551 6264 19552
rect 15944 19616 16264 19617
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 19551 16264 19552
rect 25944 19616 26264 19617
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 19551 26264 19552
rect 0 19410 480 19440
rect 11789 19410 11855 19413
rect 0 19408 11855 19410
rect 0 19352 11794 19408
rect 11850 19352 11855 19408
rect 0 19350 11855 19352
rect 0 19320 480 19350
rect 11789 19347 11855 19350
rect 25313 19410 25379 19413
rect 29520 19410 30000 19440
rect 25313 19408 30000 19410
rect 25313 19352 25318 19408
rect 25374 19352 30000 19408
rect 25313 19350 30000 19352
rect 25313 19347 25379 19350
rect 29520 19320 30000 19350
rect 8109 19274 8175 19277
rect 24117 19274 24183 19277
rect 24853 19274 24919 19277
rect 8109 19272 24919 19274
rect 8109 19216 8114 19272
rect 8170 19216 24122 19272
rect 24178 19216 24858 19272
rect 24914 19216 24919 19272
rect 8109 19214 24919 19216
rect 8109 19211 8175 19214
rect 24117 19211 24183 19214
rect 24853 19211 24919 19214
rect 10944 19072 11264 19073
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 19007 11264 19008
rect 20944 19072 21264 19073
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 19007 21264 19008
rect 0 18866 480 18896
rect 2957 18866 3023 18869
rect 0 18864 3023 18866
rect 0 18808 2962 18864
rect 3018 18808 3023 18864
rect 0 18806 3023 18808
rect 0 18776 480 18806
rect 2957 18803 3023 18806
rect 4429 18866 4495 18869
rect 12341 18866 12407 18869
rect 4429 18864 12407 18866
rect 4429 18808 4434 18864
rect 4490 18808 12346 18864
rect 12402 18808 12407 18864
rect 4429 18806 12407 18808
rect 4429 18803 4495 18806
rect 12341 18803 12407 18806
rect 14549 18866 14615 18869
rect 17309 18866 17375 18869
rect 21173 18866 21239 18869
rect 14549 18864 21239 18866
rect 14549 18808 14554 18864
rect 14610 18808 17314 18864
rect 17370 18808 21178 18864
rect 21234 18808 21239 18864
rect 14549 18806 21239 18808
rect 14549 18803 14615 18806
rect 17309 18803 17375 18806
rect 21173 18803 21239 18806
rect 26969 18866 27035 18869
rect 29520 18866 30000 18896
rect 26969 18864 30000 18866
rect 26969 18808 26974 18864
rect 27030 18808 30000 18864
rect 26969 18806 30000 18808
rect 26969 18803 27035 18806
rect 29520 18776 30000 18806
rect 2037 18730 2103 18733
rect 4521 18730 4587 18733
rect 7649 18730 7715 18733
rect 19333 18730 19399 18733
rect 25129 18730 25195 18733
rect 2037 18728 25195 18730
rect 2037 18672 2042 18728
rect 2098 18672 4526 18728
rect 4582 18672 7654 18728
rect 7710 18672 19338 18728
rect 19394 18672 25134 18728
rect 25190 18672 25195 18728
rect 2037 18670 25195 18672
rect 2037 18667 2103 18670
rect 4521 18667 4587 18670
rect 7649 18667 7715 18670
rect 19333 18667 19399 18670
rect 25129 18667 25195 18670
rect 5944 18528 6264 18529
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 18463 6264 18464
rect 15944 18528 16264 18529
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 18463 16264 18464
rect 25944 18528 26264 18529
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 18463 26264 18464
rect 17033 18458 17099 18461
rect 24209 18458 24275 18461
rect 25313 18458 25379 18461
rect 17033 18456 25379 18458
rect 17033 18400 17038 18456
rect 17094 18400 24214 18456
rect 24270 18400 25318 18456
rect 25374 18400 25379 18456
rect 17033 18398 25379 18400
rect 17033 18395 17099 18398
rect 24209 18395 24275 18398
rect 25313 18395 25379 18398
rect 0 18322 480 18352
rect 3601 18322 3667 18325
rect 14549 18322 14615 18325
rect 0 18262 2376 18322
rect 0 18232 480 18262
rect 2316 17917 2376 18262
rect 3601 18320 14615 18322
rect 3601 18264 3606 18320
rect 3662 18264 14554 18320
rect 14610 18264 14615 18320
rect 3601 18262 14615 18264
rect 3601 18259 3667 18262
rect 14549 18259 14615 18262
rect 14733 18322 14799 18325
rect 17125 18322 17191 18325
rect 14733 18320 17191 18322
rect 14733 18264 14738 18320
rect 14794 18264 17130 18320
rect 17186 18264 17191 18320
rect 14733 18262 17191 18264
rect 14733 18259 14799 18262
rect 17125 18259 17191 18262
rect 25129 18322 25195 18325
rect 29520 18322 30000 18352
rect 25129 18320 30000 18322
rect 25129 18264 25134 18320
rect 25190 18264 30000 18320
rect 25129 18262 30000 18264
rect 25129 18259 25195 18262
rect 29520 18232 30000 18262
rect 7557 18186 7623 18189
rect 23565 18186 23631 18189
rect 7557 18184 23631 18186
rect 7557 18128 7562 18184
rect 7618 18128 23570 18184
rect 23626 18128 23631 18184
rect 7557 18126 23631 18128
rect 7557 18123 7623 18126
rect 23565 18123 23631 18126
rect 3049 18050 3115 18053
rect 5625 18050 5691 18053
rect 3049 18048 5691 18050
rect 3049 17992 3054 18048
rect 3110 17992 5630 18048
rect 5686 17992 5691 18048
rect 3049 17990 5691 17992
rect 3049 17987 3115 17990
rect 5625 17987 5691 17990
rect 10944 17984 11264 17985
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 17919 11264 17920
rect 20944 17984 21264 17985
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 17919 21264 17920
rect 2313 17912 2379 17917
rect 2313 17856 2318 17912
rect 2374 17856 2379 17912
rect 2313 17851 2379 17856
rect 24025 17914 24091 17917
rect 26509 17914 26575 17917
rect 24025 17912 26575 17914
rect 24025 17856 24030 17912
rect 24086 17856 26514 17912
rect 26570 17856 26575 17912
rect 24025 17854 26575 17856
rect 24025 17851 24091 17854
rect 26509 17851 26575 17854
rect 8017 17778 8083 17781
rect 17769 17778 17835 17781
rect 8017 17776 17835 17778
rect 8017 17720 8022 17776
rect 8078 17720 17774 17776
rect 17830 17720 17835 17776
rect 8017 17718 17835 17720
rect 8017 17715 8083 17718
rect 17769 17715 17835 17718
rect 20161 17778 20227 17781
rect 26417 17778 26483 17781
rect 20161 17776 26483 17778
rect 20161 17720 20166 17776
rect 20222 17720 26422 17776
rect 26478 17720 26483 17776
rect 20161 17718 26483 17720
rect 20161 17715 20227 17718
rect 26417 17715 26483 17718
rect 0 17642 480 17672
rect 3601 17642 3667 17645
rect 0 17640 3667 17642
rect 0 17584 3606 17640
rect 3662 17584 3667 17640
rect 0 17582 3667 17584
rect 0 17552 480 17582
rect 3601 17579 3667 17582
rect 4521 17642 4587 17645
rect 10777 17642 10843 17645
rect 4521 17640 10843 17642
rect 4521 17584 4526 17640
rect 4582 17584 10782 17640
rect 10838 17584 10843 17640
rect 4521 17582 10843 17584
rect 4521 17579 4587 17582
rect 10777 17579 10843 17582
rect 14825 17642 14891 17645
rect 18229 17642 18295 17645
rect 24301 17642 24367 17645
rect 14825 17640 24367 17642
rect 14825 17584 14830 17640
rect 14886 17584 18234 17640
rect 18290 17584 24306 17640
rect 24362 17584 24367 17640
rect 14825 17582 24367 17584
rect 14825 17579 14891 17582
rect 18229 17579 18295 17582
rect 24301 17579 24367 17582
rect 25313 17642 25379 17645
rect 29520 17642 30000 17672
rect 25313 17640 30000 17642
rect 25313 17584 25318 17640
rect 25374 17584 30000 17640
rect 25313 17582 30000 17584
rect 25313 17579 25379 17582
rect 29520 17552 30000 17582
rect 10685 17506 10751 17509
rect 15745 17506 15811 17509
rect 10685 17504 15811 17506
rect 10685 17448 10690 17504
rect 10746 17448 15750 17504
rect 15806 17448 15811 17504
rect 10685 17446 15811 17448
rect 10685 17443 10751 17446
rect 15745 17443 15811 17446
rect 5944 17440 6264 17441
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 17375 6264 17376
rect 15944 17440 16264 17441
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 17375 16264 17376
rect 25944 17440 26264 17441
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 17375 26264 17376
rect 15745 17234 15811 17237
rect 2776 17232 15811 17234
rect 2776 17200 15750 17232
rect 2684 17176 15750 17200
rect 15806 17176 15811 17232
rect 2684 17174 15811 17176
rect 2684 17140 2836 17174
rect 15745 17171 15811 17174
rect 18505 17234 18571 17237
rect 23473 17234 23539 17237
rect 18505 17232 23539 17234
rect 18505 17176 18510 17232
rect 18566 17176 23478 17232
rect 23534 17176 23539 17232
rect 18505 17174 23539 17176
rect 18505 17171 18571 17174
rect 23473 17171 23539 17174
rect 0 17098 480 17128
rect 2684 17098 2744 17140
rect 0 17038 2744 17098
rect 4429 17098 4495 17101
rect 9489 17098 9555 17101
rect 4429 17096 9555 17098
rect 4429 17040 4434 17096
rect 4490 17040 9494 17096
rect 9550 17040 9555 17096
rect 4429 17038 9555 17040
rect 0 17008 480 17038
rect 4429 17035 4495 17038
rect 9489 17035 9555 17038
rect 15653 17098 15719 17101
rect 29520 17098 30000 17128
rect 15653 17096 30000 17098
rect 15653 17040 15658 17096
rect 15714 17040 30000 17096
rect 15653 17038 30000 17040
rect 15653 17035 15719 17038
rect 29520 17008 30000 17038
rect 2313 16962 2379 16965
rect 2681 16962 2747 16965
rect 8017 16962 8083 16965
rect 2313 16960 8083 16962
rect 2313 16904 2318 16960
rect 2374 16904 2686 16960
rect 2742 16904 8022 16960
rect 8078 16904 8083 16960
rect 2313 16902 8083 16904
rect 2313 16899 2379 16902
rect 2681 16899 2747 16902
rect 8017 16899 8083 16902
rect 10944 16896 11264 16897
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 16831 11264 16832
rect 20944 16896 21264 16897
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 16831 21264 16832
rect 4061 16826 4127 16829
rect 5717 16826 5783 16829
rect 4061 16824 5783 16826
rect 4061 16768 4066 16824
rect 4122 16768 5722 16824
rect 5778 16768 5783 16824
rect 4061 16766 5783 16768
rect 4061 16763 4127 16766
rect 5717 16763 5783 16766
rect 11329 16826 11395 16829
rect 14825 16826 14891 16829
rect 11329 16824 14891 16826
rect 11329 16768 11334 16824
rect 11390 16768 14830 16824
rect 14886 16768 14891 16824
rect 11329 16766 14891 16768
rect 11329 16763 11395 16766
rect 14825 16763 14891 16766
rect 2865 16690 2931 16693
rect 9857 16690 9923 16693
rect 2865 16688 9923 16690
rect 2865 16632 2870 16688
rect 2926 16632 9862 16688
rect 9918 16632 9923 16688
rect 2865 16630 9923 16632
rect 2865 16627 2931 16630
rect 9857 16627 9923 16630
rect 18597 16690 18663 16693
rect 23841 16690 23907 16693
rect 18597 16688 23907 16690
rect 18597 16632 18602 16688
rect 18658 16632 23846 16688
rect 23902 16632 23907 16688
rect 18597 16630 23907 16632
rect 18597 16627 18663 16630
rect 23841 16627 23907 16630
rect 0 16418 480 16448
rect 5533 16418 5599 16421
rect 29520 16418 30000 16448
rect 0 16416 5599 16418
rect 0 16360 5538 16416
rect 5594 16360 5599 16416
rect 0 16358 5599 16360
rect 0 16328 480 16358
rect 5533 16355 5599 16358
rect 26374 16358 30000 16418
rect 5944 16352 6264 16353
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 16287 6264 16288
rect 15944 16352 16264 16353
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 16287 16264 16288
rect 25944 16352 26264 16353
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 16287 26264 16288
rect 12709 16146 12775 16149
rect 23105 16146 23171 16149
rect 12709 16144 23171 16146
rect 12709 16088 12714 16144
rect 12770 16088 23110 16144
rect 23166 16088 23171 16144
rect 12709 16086 23171 16088
rect 12709 16083 12775 16086
rect 23105 16083 23171 16086
rect 25497 16146 25563 16149
rect 26374 16146 26434 16358
rect 29520 16328 30000 16358
rect 25497 16144 26434 16146
rect 25497 16088 25502 16144
rect 25558 16088 26434 16144
rect 25497 16086 26434 16088
rect 25497 16083 25563 16086
rect 4245 16010 4311 16013
rect 10961 16010 11027 16013
rect 14917 16010 14983 16013
rect 4245 16008 14983 16010
rect 4245 15952 4250 16008
rect 4306 15952 10966 16008
rect 11022 15952 14922 16008
rect 14978 15952 14983 16008
rect 4245 15950 14983 15952
rect 4245 15947 4311 15950
rect 10961 15947 11027 15950
rect 14917 15947 14983 15950
rect 0 15874 480 15904
rect 3877 15874 3943 15877
rect 0 15872 3943 15874
rect 0 15816 3882 15872
rect 3938 15816 3943 15872
rect 0 15814 3943 15816
rect 0 15784 480 15814
rect 3877 15811 3943 15814
rect 27429 15874 27495 15877
rect 29520 15874 30000 15904
rect 27429 15872 30000 15874
rect 27429 15816 27434 15872
rect 27490 15816 30000 15872
rect 27429 15814 30000 15816
rect 27429 15811 27495 15814
rect 10944 15808 11264 15809
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 15743 11264 15744
rect 20944 15808 21264 15809
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 29520 15784 30000 15814
rect 20944 15743 21264 15744
rect 25630 15540 25636 15604
rect 25700 15602 25706 15604
rect 25773 15602 25839 15605
rect 25700 15600 25839 15602
rect 25700 15544 25778 15600
rect 25834 15544 25839 15600
rect 25700 15542 25839 15544
rect 25700 15540 25706 15542
rect 25773 15539 25839 15542
rect 14917 15466 14983 15469
rect 18413 15466 18479 15469
rect 23749 15466 23815 15469
rect 24485 15466 24551 15469
rect 14917 15464 24551 15466
rect 14917 15408 14922 15464
rect 14978 15408 18418 15464
rect 18474 15408 23754 15464
rect 23810 15408 24490 15464
rect 24546 15408 24551 15464
rect 14917 15406 24551 15408
rect 14917 15403 14983 15406
rect 18413 15403 18479 15406
rect 23749 15403 23815 15406
rect 24485 15403 24551 15406
rect 25773 15466 25839 15469
rect 25773 15464 26434 15466
rect 25773 15408 25778 15464
rect 25834 15408 26434 15464
rect 25773 15406 26434 15408
rect 25773 15403 25839 15406
rect 0 15330 480 15360
rect 749 15330 815 15333
rect 0 15328 815 15330
rect 0 15272 754 15328
rect 810 15272 815 15328
rect 0 15270 815 15272
rect 26374 15330 26434 15406
rect 29520 15330 30000 15360
rect 26374 15270 30000 15330
rect 0 15240 480 15270
rect 749 15267 815 15270
rect 5944 15264 6264 15265
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 15199 6264 15200
rect 15944 15264 16264 15265
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 15199 16264 15200
rect 25944 15264 26264 15265
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 29520 15240 30000 15270
rect 25944 15199 26264 15200
rect 18689 14922 18755 14925
rect 23473 14922 23539 14925
rect 18689 14920 23539 14922
rect 18689 14864 18694 14920
rect 18750 14864 23478 14920
rect 23534 14864 23539 14920
rect 18689 14862 23539 14864
rect 18689 14859 18755 14862
rect 23473 14859 23539 14862
rect 25037 14924 25103 14925
rect 25037 14920 25084 14924
rect 25148 14922 25154 14924
rect 25037 14864 25042 14920
rect 25037 14860 25084 14864
rect 25148 14862 25194 14922
rect 25148 14860 25154 14862
rect 25037 14859 25103 14860
rect 10944 14720 11264 14721
rect 0 14650 480 14680
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 14655 11264 14656
rect 20944 14720 21264 14721
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 14655 21264 14656
rect 10225 14650 10291 14653
rect 0 14648 10291 14650
rect 0 14592 10230 14648
rect 10286 14592 10291 14648
rect 0 14590 10291 14592
rect 0 14560 480 14590
rect 10225 14587 10291 14590
rect 17953 14650 18019 14653
rect 19885 14650 19951 14653
rect 17953 14648 19951 14650
rect 17953 14592 17958 14648
rect 18014 14592 19890 14648
rect 19946 14592 19951 14648
rect 17953 14590 19951 14592
rect 17953 14587 18019 14590
rect 19885 14587 19951 14590
rect 24393 14650 24459 14653
rect 29520 14650 30000 14680
rect 24393 14648 30000 14650
rect 24393 14592 24398 14648
rect 24454 14592 30000 14648
rect 24393 14590 30000 14592
rect 24393 14587 24459 14590
rect 29520 14560 30000 14590
rect 5944 14176 6264 14177
rect 0 14106 480 14136
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 14111 6264 14112
rect 15944 14176 16264 14177
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 14111 16264 14112
rect 25944 14176 26264 14177
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 14111 26264 14112
rect 4061 14106 4127 14109
rect 29520 14106 30000 14136
rect 0 14104 4127 14106
rect 0 14048 4066 14104
rect 4122 14048 4127 14104
rect 0 14046 4127 14048
rect 0 14016 480 14046
rect 4061 14043 4127 14046
rect 26374 14046 30000 14106
rect 9673 13970 9739 13973
rect 11329 13970 11395 13973
rect 9673 13968 11395 13970
rect 9673 13912 9678 13968
rect 9734 13912 11334 13968
rect 11390 13912 11395 13968
rect 9673 13910 11395 13912
rect 9673 13907 9739 13910
rect 11329 13907 11395 13910
rect 14917 13970 14983 13973
rect 16665 13970 16731 13973
rect 14917 13968 16731 13970
rect 14917 13912 14922 13968
rect 14978 13912 16670 13968
rect 16726 13912 16731 13968
rect 14917 13910 16731 13912
rect 14917 13907 14983 13910
rect 16665 13907 16731 13910
rect 16849 13970 16915 13973
rect 18689 13970 18755 13973
rect 20713 13970 20779 13973
rect 16849 13968 20779 13970
rect 16849 13912 16854 13968
rect 16910 13912 18694 13968
rect 18750 13912 20718 13968
rect 20774 13912 20779 13968
rect 16849 13910 20779 13912
rect 16849 13907 16915 13910
rect 18689 13907 18755 13910
rect 20713 13907 20779 13910
rect 22553 13970 22619 13973
rect 26141 13970 26207 13973
rect 22553 13968 26207 13970
rect 22553 13912 22558 13968
rect 22614 13912 26146 13968
rect 26202 13912 26207 13968
rect 22553 13910 26207 13912
rect 22553 13907 22619 13910
rect 26141 13907 26207 13910
rect 9949 13834 10015 13837
rect 25773 13834 25839 13837
rect 26374 13834 26434 14046
rect 29520 14016 30000 14046
rect 9949 13832 25839 13834
rect 9949 13776 9954 13832
rect 10010 13776 25778 13832
rect 25834 13776 25839 13832
rect 9949 13774 25839 13776
rect 9949 13771 10015 13774
rect 25773 13771 25839 13774
rect 26006 13774 26434 13834
rect 25773 13698 25839 13701
rect 26006 13698 26066 13774
rect 25773 13696 26066 13698
rect 25773 13640 25778 13696
rect 25834 13640 26066 13696
rect 25773 13638 26066 13640
rect 25773 13635 25839 13638
rect 10944 13632 11264 13633
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 13567 11264 13568
rect 20944 13632 21264 13633
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 13567 21264 13568
rect 3325 13562 3391 13565
rect 10501 13562 10567 13565
rect 3325 13560 10567 13562
rect 3325 13504 3330 13560
rect 3386 13504 10506 13560
rect 10562 13504 10567 13560
rect 3325 13502 10567 13504
rect 3325 13499 3391 13502
rect 10501 13499 10567 13502
rect 12157 13562 12223 13565
rect 26969 13562 27035 13565
rect 12157 13560 17234 13562
rect 12157 13504 12162 13560
rect 12218 13504 17234 13560
rect 12157 13502 17234 13504
rect 12157 13499 12223 13502
rect 0 13426 480 13456
rect 3601 13426 3667 13429
rect 0 13424 3667 13426
rect 0 13368 3606 13424
rect 3662 13368 3667 13424
rect 0 13366 3667 13368
rect 0 13336 480 13366
rect 3601 13363 3667 13366
rect 4705 13426 4771 13429
rect 7557 13426 7623 13429
rect 13629 13426 13695 13429
rect 16849 13426 16915 13429
rect 4705 13424 16915 13426
rect 4705 13368 4710 13424
rect 4766 13368 7562 13424
rect 7618 13368 13634 13424
rect 13690 13368 16854 13424
rect 16910 13368 16915 13424
rect 4705 13366 16915 13368
rect 17174 13426 17234 13502
rect 21958 13560 27035 13562
rect 21958 13504 26974 13560
rect 27030 13504 27035 13560
rect 21958 13502 27035 13504
rect 21958 13426 22018 13502
rect 26969 13499 27035 13502
rect 17174 13366 22018 13426
rect 24761 13426 24827 13429
rect 29520 13426 30000 13456
rect 24761 13424 30000 13426
rect 24761 13368 24766 13424
rect 24822 13368 30000 13424
rect 24761 13366 30000 13368
rect 4705 13363 4771 13366
rect 7557 13363 7623 13366
rect 13629 13363 13695 13366
rect 16849 13363 16915 13366
rect 24761 13363 24827 13366
rect 29520 13336 30000 13366
rect 8569 13290 8635 13293
rect 10133 13290 10199 13293
rect 8569 13288 10199 13290
rect 8569 13232 8574 13288
rect 8630 13232 10138 13288
rect 10194 13232 10199 13288
rect 8569 13230 10199 13232
rect 8569 13227 8635 13230
rect 10133 13227 10199 13230
rect 16297 13290 16363 13293
rect 16297 13288 19304 13290
rect 16297 13232 16302 13288
rect 16358 13232 19304 13288
rect 16297 13230 19304 13232
rect 16297 13227 16363 13230
rect 7925 13154 7991 13157
rect 10041 13154 10107 13157
rect 7925 13152 10107 13154
rect 7925 13096 7930 13152
rect 7986 13096 10046 13152
rect 10102 13096 10107 13152
rect 7925 13094 10107 13096
rect 7925 13091 7991 13094
rect 10041 13091 10107 13094
rect 10317 13154 10383 13157
rect 15193 13154 15259 13157
rect 10317 13152 15259 13154
rect 10317 13096 10322 13152
rect 10378 13096 15198 13152
rect 15254 13096 15259 13152
rect 10317 13094 15259 13096
rect 10317 13091 10383 13094
rect 15193 13091 15259 13094
rect 5944 13088 6264 13089
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 13023 6264 13024
rect 15944 13088 16264 13089
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 13023 16264 13024
rect 19244 13018 19304 13230
rect 25944 13088 26264 13089
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 13023 26264 13024
rect 20713 13018 20779 13021
rect 25037 13018 25103 13021
rect 19244 13016 25103 13018
rect 19244 12960 20718 13016
rect 20774 12960 25042 13016
rect 25098 12960 25103 13016
rect 19244 12958 25103 12960
rect 20713 12955 20779 12958
rect 25037 12955 25103 12958
rect 0 12882 480 12912
rect 4705 12882 4771 12885
rect 0 12880 4771 12882
rect 0 12824 4710 12880
rect 4766 12824 4771 12880
rect 0 12822 4771 12824
rect 0 12792 480 12822
rect 4705 12819 4771 12822
rect 5073 12882 5139 12885
rect 7925 12882 7991 12885
rect 5073 12880 7991 12882
rect 5073 12824 5078 12880
rect 5134 12824 7930 12880
rect 7986 12824 7991 12880
rect 5073 12822 7991 12824
rect 5073 12819 5139 12822
rect 7925 12819 7991 12822
rect 8109 12882 8175 12885
rect 10317 12882 10383 12885
rect 8109 12880 10383 12882
rect 8109 12824 8114 12880
rect 8170 12824 10322 12880
rect 10378 12824 10383 12880
rect 8109 12822 10383 12824
rect 8109 12819 8175 12822
rect 10317 12819 10383 12822
rect 10501 12882 10567 12885
rect 11329 12882 11395 12885
rect 10501 12880 11395 12882
rect 10501 12824 10506 12880
rect 10562 12824 11334 12880
rect 11390 12824 11395 12880
rect 10501 12822 11395 12824
rect 10501 12819 10567 12822
rect 11329 12819 11395 12822
rect 13997 12882 14063 12885
rect 19006 12882 19012 12884
rect 13997 12880 19012 12882
rect 13997 12824 14002 12880
rect 14058 12824 19012 12880
rect 13997 12822 19012 12824
rect 13997 12819 14063 12822
rect 19006 12820 19012 12822
rect 19076 12820 19082 12884
rect 19190 12820 19196 12884
rect 19260 12882 19266 12884
rect 22093 12882 22159 12885
rect 29520 12882 30000 12912
rect 19260 12880 30000 12882
rect 19260 12824 22098 12880
rect 22154 12824 30000 12880
rect 19260 12822 30000 12824
rect 19260 12820 19266 12822
rect 22093 12819 22159 12822
rect 29520 12792 30000 12822
rect 3601 12746 3667 12749
rect 19241 12746 19307 12749
rect 21725 12746 21791 12749
rect 3601 12744 4032 12746
rect 3601 12688 3606 12744
rect 3662 12688 4032 12744
rect 3601 12686 4032 12688
rect 3601 12683 3667 12686
rect 1853 12610 1919 12613
rect 3049 12610 3115 12613
rect 3972 12610 4032 12686
rect 19241 12744 21791 12746
rect 19241 12688 19246 12744
rect 19302 12688 21730 12744
rect 21786 12688 21791 12744
rect 19241 12686 21791 12688
rect 19241 12683 19307 12686
rect 21725 12683 21791 12686
rect 4245 12610 4311 12613
rect 9673 12610 9739 12613
rect 10777 12610 10843 12613
rect 1853 12608 3802 12610
rect 1853 12552 1858 12608
rect 1914 12552 3054 12608
rect 3110 12552 3802 12608
rect 1853 12550 3802 12552
rect 3972 12608 4311 12610
rect 3972 12552 4250 12608
rect 4306 12552 4311 12608
rect 3972 12550 4311 12552
rect 1853 12547 1919 12550
rect 3049 12547 3115 12550
rect 3742 12474 3802 12550
rect 4245 12547 4311 12550
rect 5030 12608 10843 12610
rect 5030 12552 9678 12608
rect 9734 12552 10782 12608
rect 10838 12552 10843 12608
rect 5030 12550 10843 12552
rect 5030 12474 5090 12550
rect 9673 12547 9739 12550
rect 10777 12547 10843 12550
rect 11329 12610 11395 12613
rect 14641 12610 14707 12613
rect 18137 12610 18203 12613
rect 11329 12608 18203 12610
rect 11329 12552 11334 12608
rect 11390 12552 14646 12608
rect 14702 12552 18142 12608
rect 18198 12552 18203 12608
rect 11329 12550 18203 12552
rect 11329 12547 11395 12550
rect 14641 12547 14707 12550
rect 18137 12547 18203 12550
rect 19149 12610 19215 12613
rect 20713 12610 20779 12613
rect 19149 12608 20779 12610
rect 19149 12552 19154 12608
rect 19210 12552 20718 12608
rect 20774 12552 20779 12608
rect 19149 12550 20779 12552
rect 19149 12547 19215 12550
rect 20713 12547 20779 12550
rect 25129 12610 25195 12613
rect 25773 12610 25839 12613
rect 25129 12608 25839 12610
rect 25129 12552 25134 12608
rect 25190 12552 25778 12608
rect 25834 12552 25839 12608
rect 25129 12550 25839 12552
rect 25129 12547 25195 12550
rect 25773 12547 25839 12550
rect 10944 12544 11264 12545
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 12479 11264 12480
rect 20944 12544 21264 12545
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 12479 21264 12480
rect 3742 12414 5090 12474
rect 15469 12474 15535 12477
rect 21725 12474 21791 12477
rect 23473 12474 23539 12477
rect 15469 12472 20730 12474
rect 15469 12416 15474 12472
rect 15530 12416 20730 12472
rect 15469 12414 20730 12416
rect 15469 12411 15535 12414
rect 0 12338 480 12368
rect 3141 12338 3207 12341
rect 5625 12338 5691 12341
rect 0 12278 1410 12338
rect 0 12248 480 12278
rect 1350 11930 1410 12278
rect 3141 12336 5691 12338
rect 3141 12280 3146 12336
rect 3202 12280 5630 12336
rect 5686 12280 5691 12336
rect 3141 12278 5691 12280
rect 3141 12275 3207 12278
rect 5625 12275 5691 12278
rect 8845 12338 8911 12341
rect 15101 12338 15167 12341
rect 20529 12338 20595 12341
rect 8845 12336 20595 12338
rect 8845 12280 8850 12336
rect 8906 12280 15106 12336
rect 15162 12280 20534 12336
rect 20590 12280 20595 12336
rect 8845 12278 20595 12280
rect 20670 12338 20730 12414
rect 21406 12472 23539 12474
rect 21406 12416 21730 12472
rect 21786 12416 23478 12472
rect 23534 12416 23539 12472
rect 21406 12414 23539 12416
rect 21406 12338 21466 12414
rect 21725 12411 21791 12414
rect 23473 12411 23539 12414
rect 20670 12278 21466 12338
rect 27337 12338 27403 12341
rect 29520 12338 30000 12368
rect 27337 12336 30000 12338
rect 27337 12280 27342 12336
rect 27398 12280 30000 12336
rect 27337 12278 30000 12280
rect 8845 12275 8911 12278
rect 15101 12275 15167 12278
rect 20529 12275 20595 12278
rect 27337 12275 27403 12278
rect 29520 12248 30000 12278
rect 3969 12202 4035 12205
rect 12525 12202 12591 12205
rect 15469 12202 15535 12205
rect 3969 12200 15535 12202
rect 3969 12144 3974 12200
rect 4030 12144 12530 12200
rect 12586 12144 15474 12200
rect 15530 12144 15535 12200
rect 3969 12142 15535 12144
rect 3969 12139 4035 12142
rect 12525 12139 12591 12142
rect 15469 12139 15535 12142
rect 15653 12202 15719 12205
rect 25037 12202 25103 12205
rect 15653 12200 25103 12202
rect 15653 12144 15658 12200
rect 15714 12144 25042 12200
rect 25098 12144 25103 12200
rect 15653 12142 25103 12144
rect 15653 12139 15719 12142
rect 25037 12139 25103 12142
rect 25221 12202 25287 12205
rect 27613 12202 27679 12205
rect 25221 12200 27679 12202
rect 25221 12144 25226 12200
rect 25282 12144 27618 12200
rect 27674 12144 27679 12200
rect 25221 12142 27679 12144
rect 25221 12139 25287 12142
rect 27613 12139 27679 12142
rect 2313 12066 2379 12069
rect 4429 12066 4495 12069
rect 25037 12068 25103 12069
rect 25037 12066 25084 12068
rect 2313 12064 4495 12066
rect 2313 12008 2318 12064
rect 2374 12008 4434 12064
rect 4490 12008 4495 12064
rect 2313 12006 4495 12008
rect 24992 12064 25084 12066
rect 24992 12008 25042 12064
rect 24992 12006 25084 12008
rect 2313 12003 2379 12006
rect 4429 12003 4495 12006
rect 25037 12004 25084 12006
rect 25148 12004 25154 12068
rect 25037 12003 25103 12004
rect 5944 12000 6264 12001
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 11935 6264 11936
rect 15944 12000 16264 12001
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 11935 16264 11936
rect 25944 12000 26264 12001
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 11935 26264 11936
rect 4153 11930 4219 11933
rect 1350 11928 4219 11930
rect 1350 11872 4158 11928
rect 4214 11872 4219 11928
rect 1350 11870 4219 11872
rect 4153 11867 4219 11870
rect 2129 11794 2195 11797
rect 13629 11794 13695 11797
rect 2129 11792 13695 11794
rect 2129 11736 2134 11792
rect 2190 11736 13634 11792
rect 13690 11736 13695 11792
rect 2129 11734 13695 11736
rect 2129 11731 2195 11734
rect 13629 11731 13695 11734
rect 22001 11794 22067 11797
rect 25773 11794 25839 11797
rect 22001 11792 25839 11794
rect 22001 11736 22006 11792
rect 22062 11736 25778 11792
rect 25834 11736 25839 11792
rect 22001 11734 25839 11736
rect 22001 11731 22067 11734
rect 25773 11731 25839 11734
rect 0 11658 480 11688
rect 3509 11658 3575 11661
rect 21265 11658 21331 11661
rect 0 11656 3575 11658
rect 0 11600 3514 11656
rect 3570 11600 3575 11656
rect 0 11598 3575 11600
rect 0 11568 480 11598
rect 3509 11595 3575 11598
rect 4524 11656 21331 11658
rect 4524 11600 21270 11656
rect 21326 11600 21331 11656
rect 4524 11598 21331 11600
rect 2773 11522 2839 11525
rect 4524 11522 4584 11598
rect 21265 11595 21331 11598
rect 26693 11658 26759 11661
rect 29520 11658 30000 11688
rect 26693 11656 30000 11658
rect 26693 11600 26698 11656
rect 26754 11600 30000 11656
rect 26693 11598 30000 11600
rect 26693 11595 26759 11598
rect 29520 11568 30000 11598
rect 2773 11520 4584 11522
rect 2773 11464 2778 11520
rect 2834 11464 4584 11520
rect 2773 11462 4584 11464
rect 7189 11522 7255 11525
rect 9673 11522 9739 11525
rect 7189 11520 9739 11522
rect 7189 11464 7194 11520
rect 7250 11464 9678 11520
rect 9734 11464 9739 11520
rect 7189 11462 9739 11464
rect 2773 11459 2839 11462
rect 7189 11459 7255 11462
rect 9673 11459 9739 11462
rect 25221 11522 25287 11525
rect 25630 11522 25636 11524
rect 25221 11520 25636 11522
rect 25221 11464 25226 11520
rect 25282 11464 25636 11520
rect 25221 11462 25636 11464
rect 25221 11459 25287 11462
rect 25630 11460 25636 11462
rect 25700 11460 25706 11524
rect 10944 11456 11264 11457
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 11391 11264 11392
rect 20944 11456 21264 11457
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 11391 21264 11392
rect 25497 11386 25563 11389
rect 21958 11384 25563 11386
rect 21958 11328 25502 11384
rect 25558 11328 25563 11384
rect 21958 11326 25563 11328
rect 2773 11250 2839 11253
rect 12157 11250 12223 11253
rect 2773 11248 12223 11250
rect 2773 11192 2778 11248
rect 2834 11192 12162 11248
rect 12218 11192 12223 11248
rect 2773 11190 12223 11192
rect 2773 11187 2839 11190
rect 12157 11187 12223 11190
rect 15469 11250 15535 11253
rect 16389 11250 16455 11253
rect 21958 11250 22018 11326
rect 25497 11323 25563 11326
rect 15469 11248 22018 11250
rect 15469 11192 15474 11248
rect 15530 11192 16394 11248
rect 16450 11192 22018 11248
rect 15469 11190 22018 11192
rect 15469 11187 15535 11190
rect 16389 11187 16455 11190
rect 0 11114 480 11144
rect 1577 11114 1643 11117
rect 0 11112 1643 11114
rect 0 11056 1582 11112
rect 1638 11056 1643 11112
rect 0 11054 1643 11056
rect 0 11024 480 11054
rect 1577 11051 1643 11054
rect 2957 11114 3023 11117
rect 21725 11114 21791 11117
rect 2957 11112 21791 11114
rect 2957 11056 2962 11112
rect 3018 11056 21730 11112
rect 21786 11056 21791 11112
rect 2957 11054 21791 11056
rect 2957 11051 3023 11054
rect 21725 11051 21791 11054
rect 25865 11114 25931 11117
rect 29520 11114 30000 11144
rect 25865 11112 30000 11114
rect 25865 11056 25870 11112
rect 25926 11056 30000 11112
rect 25865 11054 30000 11056
rect 25865 11051 25931 11054
rect 29520 11024 30000 11054
rect 19517 10978 19583 10981
rect 24945 10978 25011 10981
rect 19517 10976 25011 10978
rect 19517 10920 19522 10976
rect 19578 10920 24950 10976
rect 25006 10920 25011 10976
rect 19517 10918 25011 10920
rect 19517 10915 19583 10918
rect 24945 10915 25011 10918
rect 5944 10912 6264 10913
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 10847 6264 10848
rect 15944 10912 16264 10913
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 10847 16264 10848
rect 25944 10912 26264 10913
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 10847 26264 10848
rect 16481 10842 16547 10845
rect 21449 10842 21515 10845
rect 16481 10840 21515 10842
rect 16481 10784 16486 10840
rect 16542 10784 21454 10840
rect 21510 10784 21515 10840
rect 16481 10782 21515 10784
rect 16481 10779 16547 10782
rect 21449 10779 21515 10782
rect 10593 10706 10659 10709
rect 15653 10706 15719 10709
rect 10593 10704 15719 10706
rect 10593 10648 10598 10704
rect 10654 10648 15658 10704
rect 15714 10648 15719 10704
rect 10593 10646 15719 10648
rect 10593 10643 10659 10646
rect 15653 10643 15719 10646
rect 19057 10706 19123 10709
rect 27521 10706 27587 10709
rect 19057 10704 27587 10706
rect 19057 10648 19062 10704
rect 19118 10648 27526 10704
rect 27582 10648 27587 10704
rect 19057 10646 27587 10648
rect 19057 10643 19123 10646
rect 27521 10643 27587 10646
rect 3693 10570 3759 10573
rect 7465 10570 7531 10573
rect 15377 10570 15443 10573
rect 3693 10568 15443 10570
rect 3693 10512 3698 10568
rect 3754 10512 7470 10568
rect 7526 10512 15382 10568
rect 15438 10512 15443 10568
rect 3693 10510 15443 10512
rect 3693 10507 3759 10510
rect 7465 10507 7531 10510
rect 15377 10507 15443 10510
rect 0 10434 480 10464
rect 1577 10434 1643 10437
rect 0 10432 1643 10434
rect 0 10376 1582 10432
rect 1638 10376 1643 10432
rect 0 10374 1643 10376
rect 0 10344 480 10374
rect 1577 10371 1643 10374
rect 7281 10434 7347 10437
rect 7925 10434 7991 10437
rect 9857 10434 9923 10437
rect 7281 10432 9923 10434
rect 7281 10376 7286 10432
rect 7342 10376 7930 10432
rect 7986 10376 9862 10432
rect 9918 10376 9923 10432
rect 7281 10374 9923 10376
rect 7281 10371 7347 10374
rect 7925 10371 7991 10374
rect 9857 10371 9923 10374
rect 11973 10434 12039 10437
rect 15653 10434 15719 10437
rect 11973 10432 15719 10434
rect 11973 10376 11978 10432
rect 12034 10376 15658 10432
rect 15714 10376 15719 10432
rect 11973 10374 15719 10376
rect 11973 10371 12039 10374
rect 15653 10371 15719 10374
rect 26601 10434 26667 10437
rect 29520 10434 30000 10464
rect 26601 10432 30000 10434
rect 26601 10376 26606 10432
rect 26662 10376 30000 10432
rect 26601 10374 30000 10376
rect 26601 10371 26667 10374
rect 10944 10368 11264 10369
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 10303 11264 10304
rect 20944 10368 21264 10369
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 29520 10344 30000 10374
rect 20944 10303 21264 10304
rect 15377 10298 15443 10301
rect 15837 10298 15903 10301
rect 19057 10300 19123 10301
rect 15377 10296 15903 10298
rect 15377 10240 15382 10296
rect 15438 10240 15842 10296
rect 15898 10240 15903 10296
rect 15377 10238 15903 10240
rect 15377 10235 15443 10238
rect 15837 10235 15903 10238
rect 19006 10236 19012 10300
rect 19076 10298 19123 10300
rect 21357 10298 21423 10301
rect 24209 10298 24275 10301
rect 19076 10296 19168 10298
rect 19118 10240 19168 10296
rect 19076 10238 19168 10240
rect 21357 10296 24275 10298
rect 21357 10240 21362 10296
rect 21418 10240 24214 10296
rect 24270 10240 24275 10296
rect 21357 10238 24275 10240
rect 19076 10236 19123 10238
rect 19057 10235 19123 10236
rect 21357 10235 21423 10238
rect 24209 10235 24275 10238
rect 7465 10162 7531 10165
rect 15653 10162 15719 10165
rect 26509 10162 26575 10165
rect 7465 10160 12266 10162
rect 7465 10104 7470 10160
rect 7526 10104 12266 10160
rect 7465 10102 12266 10104
rect 7465 10099 7531 10102
rect 12206 10060 12266 10102
rect 15653 10160 26575 10162
rect 15653 10104 15658 10160
rect 15714 10104 26514 10160
rect 26570 10104 26575 10160
rect 15653 10102 26575 10104
rect 15653 10099 15719 10102
rect 26509 10099 26575 10102
rect 12206 10026 12450 10060
rect 19149 10026 19215 10029
rect 21541 10026 21607 10029
rect 12206 10024 21607 10026
rect 12206 10000 19154 10024
rect 12390 9968 19154 10000
rect 19210 9968 21546 10024
rect 21602 9968 21607 10024
rect 12390 9966 21607 9968
rect 19149 9963 19215 9966
rect 21541 9963 21607 9966
rect 23565 10026 23631 10029
rect 26417 10026 26483 10029
rect 23565 10024 26483 10026
rect 23565 9968 23570 10024
rect 23626 9968 26422 10024
rect 26478 9968 26483 10024
rect 23565 9966 26483 9968
rect 23565 9963 23631 9966
rect 26417 9963 26483 9966
rect 0 9890 480 9920
rect 2681 9890 2747 9893
rect 0 9888 2747 9890
rect 0 9832 2686 9888
rect 2742 9832 2747 9888
rect 0 9830 2747 9832
rect 0 9800 480 9830
rect 2681 9827 2747 9830
rect 26693 9890 26759 9893
rect 29520 9890 30000 9920
rect 26693 9888 30000 9890
rect 26693 9832 26698 9888
rect 26754 9832 30000 9888
rect 26693 9830 30000 9832
rect 26693 9827 26759 9830
rect 5944 9824 6264 9825
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 9759 6264 9760
rect 15944 9824 16264 9825
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 9759 16264 9760
rect 25944 9824 26264 9825
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 29520 9800 30000 9830
rect 25944 9759 26264 9760
rect 8569 9754 8635 9757
rect 8158 9752 8635 9754
rect 8158 9696 8574 9752
rect 8630 9696 8635 9752
rect 8158 9694 8635 9696
rect 3141 9618 3207 9621
rect 6545 9618 6611 9621
rect 3141 9616 6611 9618
rect 3141 9560 3146 9616
rect 3202 9560 6550 9616
rect 6606 9560 6611 9616
rect 3141 9558 6611 9560
rect 8158 9618 8218 9694
rect 8569 9691 8635 9694
rect 8569 9618 8635 9621
rect 8158 9616 8635 9618
rect 8158 9560 8574 9616
rect 8630 9560 8635 9616
rect 8158 9558 8635 9560
rect 3141 9555 3207 9558
rect 6545 9555 6611 9558
rect 8569 9555 8635 9558
rect 19149 9618 19215 9621
rect 21817 9618 21883 9621
rect 19149 9616 21883 9618
rect 19149 9560 19154 9616
rect 19210 9560 21822 9616
rect 21878 9560 21883 9616
rect 19149 9558 21883 9560
rect 19149 9555 19215 9558
rect 21817 9555 21883 9558
rect 22553 9618 22619 9621
rect 26969 9618 27035 9621
rect 22553 9616 27035 9618
rect 22553 9560 22558 9616
rect 22614 9560 26974 9616
rect 27030 9560 27035 9616
rect 22553 9558 27035 9560
rect 22553 9555 22619 9558
rect 26969 9555 27035 9558
rect 2957 9482 3023 9485
rect 7833 9482 7899 9485
rect 10317 9482 10383 9485
rect 19333 9482 19399 9485
rect 2957 9480 19399 9482
rect 2957 9424 2962 9480
rect 3018 9424 7838 9480
rect 7894 9424 10322 9480
rect 10378 9424 19338 9480
rect 19394 9424 19399 9480
rect 2957 9422 19399 9424
rect 2957 9419 3023 9422
rect 7833 9419 7899 9422
rect 10317 9419 10383 9422
rect 19333 9419 19399 9422
rect 0 9346 480 9376
rect 1577 9346 1643 9349
rect 0 9344 1643 9346
rect 0 9288 1582 9344
rect 1638 9288 1643 9344
rect 0 9286 1643 9288
rect 0 9256 480 9286
rect 1577 9283 1643 9286
rect 5625 9346 5691 9349
rect 7557 9346 7623 9349
rect 5625 9344 7623 9346
rect 5625 9288 5630 9344
rect 5686 9288 7562 9344
rect 7618 9288 7623 9344
rect 5625 9286 7623 9288
rect 5625 9283 5691 9286
rect 7557 9283 7623 9286
rect 26693 9346 26759 9349
rect 29520 9346 30000 9376
rect 26693 9344 30000 9346
rect 26693 9288 26698 9344
rect 26754 9288 30000 9344
rect 26693 9286 30000 9288
rect 26693 9283 26759 9286
rect 10944 9280 11264 9281
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 9215 11264 9216
rect 20944 9280 21264 9281
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 29520 9256 30000 9286
rect 20944 9215 21264 9216
rect 2037 9074 2103 9077
rect 24117 9074 24183 9077
rect 2037 9072 24183 9074
rect 2037 9016 2042 9072
rect 2098 9016 24122 9072
rect 24178 9016 24183 9072
rect 2037 9014 24183 9016
rect 2037 9011 2103 9014
rect 24117 9011 24183 9014
rect 3049 8938 3115 8941
rect 9857 8938 9923 8941
rect 3049 8936 9923 8938
rect 3049 8880 3054 8936
rect 3110 8880 9862 8936
rect 9918 8880 9923 8936
rect 3049 8878 9923 8880
rect 3049 8875 3115 8878
rect 9857 8875 9923 8878
rect 14641 8938 14707 8941
rect 15653 8938 15719 8941
rect 16757 8938 16823 8941
rect 14641 8936 16823 8938
rect 14641 8880 14646 8936
rect 14702 8880 15658 8936
rect 15714 8880 16762 8936
rect 16818 8880 16823 8936
rect 14641 8878 16823 8880
rect 14641 8875 14707 8878
rect 15653 8875 15719 8878
rect 16757 8875 16823 8878
rect 19241 8802 19307 8805
rect 20713 8802 20779 8805
rect 21357 8802 21423 8805
rect 19241 8800 21423 8802
rect 19241 8744 19246 8800
rect 19302 8744 20718 8800
rect 20774 8744 21362 8800
rect 21418 8744 21423 8800
rect 19241 8742 21423 8744
rect 19241 8739 19307 8742
rect 20713 8739 20779 8742
rect 21357 8739 21423 8742
rect 5944 8736 6264 8737
rect 0 8666 480 8696
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 8671 6264 8672
rect 15944 8736 16264 8737
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 8671 16264 8672
rect 25944 8736 26264 8737
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 8671 26264 8672
rect 1485 8666 1551 8669
rect 0 8664 1551 8666
rect 0 8608 1490 8664
rect 1546 8608 1551 8664
rect 0 8606 1551 8608
rect 0 8576 480 8606
rect 1485 8603 1551 8606
rect 13905 8666 13971 8669
rect 26693 8666 26759 8669
rect 29520 8666 30000 8696
rect 13905 8664 15762 8666
rect 13905 8608 13910 8664
rect 13966 8608 15762 8664
rect 13905 8606 15762 8608
rect 13905 8603 13971 8606
rect 2405 8530 2471 8533
rect 15561 8530 15627 8533
rect 2405 8528 15627 8530
rect 2405 8472 2410 8528
rect 2466 8472 15566 8528
rect 15622 8472 15627 8528
rect 2405 8470 15627 8472
rect 15702 8530 15762 8606
rect 26693 8664 30000 8666
rect 26693 8608 26698 8664
rect 26754 8608 30000 8664
rect 26693 8606 30000 8608
rect 26693 8603 26759 8606
rect 29520 8576 30000 8606
rect 21909 8530 21975 8533
rect 15702 8528 21975 8530
rect 15702 8472 21914 8528
rect 21970 8472 21975 8528
rect 15702 8470 21975 8472
rect 2405 8467 2471 8470
rect 15561 8467 15627 8470
rect 21909 8467 21975 8470
rect 10944 8192 11264 8193
rect 0 8122 480 8152
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 8127 11264 8128
rect 20944 8192 21264 8193
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 8127 21264 8128
rect 1577 8122 1643 8125
rect 0 8120 1643 8122
rect 0 8064 1582 8120
rect 1638 8064 1643 8120
rect 0 8062 1643 8064
rect 0 8032 480 8062
rect 1577 8059 1643 8062
rect 27705 8122 27771 8125
rect 29520 8122 30000 8152
rect 27705 8120 30000 8122
rect 27705 8064 27710 8120
rect 27766 8064 30000 8120
rect 27705 8062 30000 8064
rect 27705 8059 27771 8062
rect 29520 8032 30000 8062
rect 19057 7986 19123 7989
rect 25221 7986 25287 7989
rect 19057 7984 25287 7986
rect 19057 7928 19062 7984
rect 19118 7928 25226 7984
rect 25282 7928 25287 7984
rect 19057 7926 25287 7928
rect 19057 7923 19123 7926
rect 25221 7923 25287 7926
rect 5944 7648 6264 7649
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 7583 6264 7584
rect 15944 7648 16264 7649
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 7583 16264 7584
rect 25944 7648 26264 7649
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 7583 26264 7584
rect 7281 7578 7347 7581
rect 14365 7578 14431 7581
rect 7281 7576 14431 7578
rect 7281 7520 7286 7576
rect 7342 7520 14370 7576
rect 14426 7520 14431 7576
rect 7281 7518 14431 7520
rect 7281 7515 7347 7518
rect 14365 7515 14431 7518
rect 0 7442 480 7472
rect 1393 7442 1459 7445
rect 0 7440 1459 7442
rect 0 7384 1398 7440
rect 1454 7384 1459 7440
rect 0 7382 1459 7384
rect 0 7352 480 7382
rect 1393 7379 1459 7382
rect 1945 7442 2011 7445
rect 6637 7442 6703 7445
rect 1945 7440 6703 7442
rect 1945 7384 1950 7440
rect 2006 7384 6642 7440
rect 6698 7384 6703 7440
rect 1945 7382 6703 7384
rect 1945 7379 2011 7382
rect 6637 7379 6703 7382
rect 16665 7442 16731 7445
rect 18505 7442 18571 7445
rect 24209 7442 24275 7445
rect 26325 7442 26391 7445
rect 16665 7440 26391 7442
rect 16665 7384 16670 7440
rect 16726 7384 18510 7440
rect 18566 7384 24214 7440
rect 24270 7384 26330 7440
rect 26386 7384 26391 7440
rect 16665 7382 26391 7384
rect 16665 7379 16731 7382
rect 18505 7379 18571 7382
rect 24209 7379 24275 7382
rect 26325 7379 26391 7382
rect 26693 7442 26759 7445
rect 29520 7442 30000 7472
rect 26693 7440 30000 7442
rect 26693 7384 26698 7440
rect 26754 7384 30000 7440
rect 26693 7382 30000 7384
rect 26693 7379 26759 7382
rect 29520 7352 30000 7382
rect 13445 7306 13511 7309
rect 18413 7306 18479 7309
rect 25957 7306 26023 7309
rect 7054 7304 26023 7306
rect 7054 7248 13450 7304
rect 13506 7248 18418 7304
rect 18474 7248 25962 7304
rect 26018 7248 26023 7304
rect 7054 7246 26023 7248
rect 3785 7034 3851 7037
rect 5809 7034 5875 7037
rect 6177 7034 6243 7037
rect 7054 7034 7114 7246
rect 13445 7243 13511 7246
rect 18413 7243 18479 7246
rect 25957 7243 26023 7246
rect 12157 7170 12223 7173
rect 13353 7170 13419 7173
rect 12157 7168 13419 7170
rect 12157 7112 12162 7168
rect 12218 7112 13358 7168
rect 13414 7112 13419 7168
rect 12157 7110 13419 7112
rect 12157 7107 12223 7110
rect 13353 7107 13419 7110
rect 14917 7170 14983 7173
rect 19057 7170 19123 7173
rect 14917 7168 19123 7170
rect 14917 7112 14922 7168
rect 14978 7112 19062 7168
rect 19118 7112 19123 7168
rect 14917 7110 19123 7112
rect 14917 7107 14983 7110
rect 19057 7107 19123 7110
rect 10944 7104 11264 7105
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 7039 11264 7040
rect 20944 7104 21264 7105
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 7039 21264 7040
rect 3785 7032 7114 7034
rect 3785 6976 3790 7032
rect 3846 6976 5814 7032
rect 5870 6976 6182 7032
rect 6238 6976 7114 7032
rect 3785 6974 7114 6976
rect 3785 6971 3851 6974
rect 5809 6971 5875 6974
rect 6177 6971 6243 6974
rect 0 6898 480 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 480 6838
rect 1577 6835 1643 6838
rect 10317 6898 10383 6901
rect 12341 6898 12407 6901
rect 10317 6896 12407 6898
rect 10317 6840 10322 6896
rect 10378 6840 12346 6896
rect 12402 6840 12407 6896
rect 10317 6838 12407 6840
rect 10317 6835 10383 6838
rect 12341 6835 12407 6838
rect 25497 6898 25563 6901
rect 29520 6898 30000 6928
rect 25497 6896 30000 6898
rect 25497 6840 25502 6896
rect 25558 6840 30000 6896
rect 25497 6838 30000 6840
rect 25497 6835 25563 6838
rect 29520 6808 30000 6838
rect 2037 6762 2103 6765
rect 4521 6762 4587 6765
rect 11789 6762 11855 6765
rect 16113 6762 16179 6765
rect 2037 6760 16179 6762
rect 2037 6704 2042 6760
rect 2098 6704 4526 6760
rect 4582 6704 11794 6760
rect 11850 6704 16118 6760
rect 16174 6704 16179 6760
rect 2037 6702 16179 6704
rect 2037 6699 2103 6702
rect 4521 6699 4587 6702
rect 11789 6699 11855 6702
rect 16113 6699 16179 6702
rect 5944 6560 6264 6561
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 6495 6264 6496
rect 15944 6560 16264 6561
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 6495 16264 6496
rect 25944 6560 26264 6561
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 6495 26264 6496
rect 18505 6490 18571 6493
rect 24117 6490 24183 6493
rect 18505 6488 24183 6490
rect 18505 6432 18510 6488
rect 18566 6432 24122 6488
rect 24178 6432 24183 6488
rect 18505 6430 24183 6432
rect 18505 6427 18571 6430
rect 24117 6427 24183 6430
rect 0 6354 480 6384
rect 1853 6354 1919 6357
rect 0 6352 1919 6354
rect 0 6296 1858 6352
rect 1914 6296 1919 6352
rect 0 6294 1919 6296
rect 0 6264 480 6294
rect 1853 6291 1919 6294
rect 15837 6354 15903 6357
rect 26233 6354 26299 6357
rect 29520 6354 30000 6384
rect 15837 6352 26299 6354
rect 15837 6296 15842 6352
rect 15898 6296 26238 6352
rect 26294 6296 26299 6352
rect 15837 6294 26299 6296
rect 15837 6291 15903 6294
rect 26233 6291 26299 6294
rect 26558 6294 30000 6354
rect 6269 6218 6335 6221
rect 12709 6218 12775 6221
rect 23841 6218 23907 6221
rect 6269 6216 12404 6218
rect 6269 6160 6274 6216
rect 6330 6184 12404 6216
rect 12709 6216 23907 6218
rect 6330 6160 12450 6184
rect 6269 6158 12450 6160
rect 6269 6155 6335 6158
rect 12344 6124 12450 6158
rect 12709 6160 12714 6216
rect 12770 6160 23846 6216
rect 23902 6160 23907 6216
rect 12709 6158 23907 6160
rect 12709 6155 12775 6158
rect 23841 6155 23907 6158
rect 25773 6218 25839 6221
rect 26558 6218 26618 6294
rect 29520 6264 30000 6294
rect 25773 6216 26618 6218
rect 25773 6160 25778 6216
rect 25834 6160 26618 6216
rect 25773 6158 26618 6160
rect 25773 6155 25839 6158
rect 12390 6082 12450 6124
rect 17953 6082 18019 6085
rect 12390 6080 18019 6082
rect 12390 6024 17958 6080
rect 18014 6024 18019 6080
rect 12390 6022 18019 6024
rect 17953 6019 18019 6022
rect 10944 6016 11264 6017
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 5951 11264 5952
rect 20944 6016 21264 6017
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 5951 21264 5952
rect 7465 5810 7531 5813
rect 19517 5810 19583 5813
rect 20529 5810 20595 5813
rect 26509 5810 26575 5813
rect 7465 5808 20595 5810
rect 7465 5752 7470 5808
rect 7526 5752 19522 5808
rect 19578 5752 20534 5808
rect 20590 5752 20595 5808
rect 7465 5750 20595 5752
rect 7465 5747 7531 5750
rect 19517 5747 19583 5750
rect 20529 5747 20595 5750
rect 20670 5808 26575 5810
rect 20670 5752 26514 5808
rect 26570 5752 26575 5808
rect 20670 5750 26575 5752
rect 0 5674 480 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 480 5614
rect 1577 5611 1643 5614
rect 10961 5674 11027 5677
rect 15469 5674 15535 5677
rect 20670 5674 20730 5750
rect 26509 5747 26575 5750
rect 10961 5672 20730 5674
rect 10961 5616 10966 5672
rect 11022 5616 15474 5672
rect 15530 5616 20730 5672
rect 10961 5614 20730 5616
rect 22001 5674 22067 5677
rect 23749 5674 23815 5677
rect 22001 5672 23815 5674
rect 22001 5616 22006 5672
rect 22062 5616 23754 5672
rect 23810 5616 23815 5672
rect 22001 5614 23815 5616
rect 10961 5611 11027 5614
rect 15469 5611 15535 5614
rect 22001 5611 22067 5614
rect 23749 5611 23815 5614
rect 26601 5674 26667 5677
rect 29520 5674 30000 5704
rect 26601 5672 30000 5674
rect 26601 5616 26606 5672
rect 26662 5616 30000 5672
rect 26601 5614 30000 5616
rect 26601 5611 26667 5614
rect 29520 5584 30000 5614
rect 2221 5538 2287 5541
rect 4705 5538 4771 5541
rect 2221 5536 4771 5538
rect 2221 5480 2226 5536
rect 2282 5480 4710 5536
rect 4766 5480 4771 5536
rect 2221 5478 4771 5480
rect 2221 5475 2287 5478
rect 4705 5475 4771 5478
rect 16481 5538 16547 5541
rect 23933 5538 23999 5541
rect 16481 5536 23999 5538
rect 16481 5480 16486 5536
rect 16542 5480 23938 5536
rect 23994 5480 23999 5536
rect 16481 5478 23999 5480
rect 16481 5475 16547 5478
rect 23933 5475 23999 5478
rect 5944 5472 6264 5473
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 5407 6264 5408
rect 15944 5472 16264 5473
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 5407 16264 5408
rect 25944 5472 26264 5473
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 5407 26264 5408
rect 7741 5402 7807 5405
rect 16665 5402 16731 5405
rect 24761 5402 24827 5405
rect 7741 5400 15762 5402
rect 7741 5344 7746 5400
rect 7802 5344 15762 5400
rect 7741 5342 15762 5344
rect 7741 5339 7807 5342
rect 4337 5266 4403 5269
rect 15193 5266 15259 5269
rect 4337 5264 15259 5266
rect 4337 5208 4342 5264
rect 4398 5208 15198 5264
rect 15254 5208 15259 5264
rect 4337 5206 15259 5208
rect 15702 5266 15762 5342
rect 16665 5400 24827 5402
rect 16665 5344 16670 5400
rect 16726 5344 24766 5400
rect 24822 5344 24827 5400
rect 16665 5342 24827 5344
rect 16665 5339 16731 5342
rect 24761 5339 24827 5342
rect 20345 5266 20411 5269
rect 26417 5266 26483 5269
rect 15702 5264 26483 5266
rect 15702 5208 20350 5264
rect 20406 5208 26422 5264
rect 26478 5208 26483 5264
rect 15702 5206 26483 5208
rect 4337 5203 4403 5206
rect 15193 5203 15259 5206
rect 20345 5203 20411 5206
rect 26417 5203 26483 5206
rect 0 5130 480 5160
rect 1577 5130 1643 5133
rect 0 5128 1643 5130
rect 0 5072 1582 5128
rect 1638 5072 1643 5128
rect 0 5070 1643 5072
rect 0 5040 480 5070
rect 1577 5067 1643 5070
rect 4705 5130 4771 5133
rect 13445 5130 13511 5133
rect 15561 5130 15627 5133
rect 22001 5130 22067 5133
rect 4705 5128 13511 5130
rect 4705 5072 4710 5128
rect 4766 5072 13450 5128
rect 13506 5072 13511 5128
rect 4705 5070 13511 5072
rect 4705 5067 4771 5070
rect 13445 5067 13511 5070
rect 13678 5128 22067 5130
rect 13678 5072 15566 5128
rect 15622 5072 22006 5128
rect 22062 5072 22067 5128
rect 13678 5070 22067 5072
rect 13537 4994 13603 4997
rect 13678 4994 13738 5070
rect 15561 5067 15627 5070
rect 22001 5067 22067 5070
rect 23933 5130 23999 5133
rect 26509 5130 26575 5133
rect 23933 5128 26575 5130
rect 23933 5072 23938 5128
rect 23994 5072 26514 5128
rect 26570 5072 26575 5128
rect 23933 5070 26575 5072
rect 23933 5067 23999 5070
rect 26509 5067 26575 5070
rect 26693 5130 26759 5133
rect 29520 5130 30000 5160
rect 26693 5128 30000 5130
rect 26693 5072 26698 5128
rect 26754 5072 30000 5128
rect 26693 5070 30000 5072
rect 26693 5067 26759 5070
rect 29520 5040 30000 5070
rect 13537 4992 13738 4994
rect 13537 4936 13542 4992
rect 13598 4936 13738 4992
rect 13537 4934 13738 4936
rect 13537 4931 13603 4934
rect 10944 4928 11264 4929
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 4863 11264 4864
rect 20944 4928 21264 4929
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 4863 21264 4864
rect 2037 4722 2103 4725
rect 12157 4722 12223 4725
rect 2037 4720 12223 4722
rect 2037 4664 2042 4720
rect 2098 4664 12162 4720
rect 12218 4664 12223 4720
rect 2037 4662 12223 4664
rect 2037 4659 2103 4662
rect 12157 4659 12223 4662
rect 19885 4586 19951 4589
rect 24945 4586 25011 4589
rect 19885 4584 25011 4586
rect 19885 4528 19890 4584
rect 19946 4528 24950 4584
rect 25006 4528 25011 4584
rect 19885 4526 25011 4528
rect 19885 4523 19951 4526
rect 24945 4523 25011 4526
rect 0 4450 480 4480
rect 1485 4450 1551 4453
rect 0 4448 1551 4450
rect 0 4392 1490 4448
rect 1546 4392 1551 4448
rect 0 4390 1551 4392
rect 0 4360 480 4390
rect 1485 4387 1551 4390
rect 16665 4450 16731 4453
rect 20713 4450 20779 4453
rect 16665 4448 20779 4450
rect 16665 4392 16670 4448
rect 16726 4392 20718 4448
rect 20774 4392 20779 4448
rect 16665 4390 20779 4392
rect 16665 4387 16731 4390
rect 20713 4387 20779 4390
rect 27521 4450 27587 4453
rect 29520 4450 30000 4480
rect 27521 4448 30000 4450
rect 27521 4392 27526 4448
rect 27582 4392 30000 4448
rect 27521 4390 30000 4392
rect 27521 4387 27587 4390
rect 5944 4384 6264 4385
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 4319 6264 4320
rect 15944 4384 16264 4385
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 4319 16264 4320
rect 25944 4384 26264 4385
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 29520 4360 30000 4390
rect 25944 4319 26264 4320
rect 2129 4178 2195 4181
rect 10041 4178 10107 4181
rect 2129 4176 10107 4178
rect 2129 4120 2134 4176
rect 2190 4120 10046 4176
rect 10102 4120 10107 4176
rect 2129 4118 10107 4120
rect 2129 4115 2195 4118
rect 10041 4115 10107 4118
rect 16389 4178 16455 4181
rect 19241 4178 19307 4181
rect 16389 4176 19307 4178
rect 16389 4120 16394 4176
rect 16450 4120 19246 4176
rect 19302 4120 19307 4176
rect 16389 4118 19307 4120
rect 16389 4115 16455 4118
rect 19241 4115 19307 4118
rect 26693 4178 26759 4181
rect 26693 4176 26802 4178
rect 26693 4120 26698 4176
rect 26754 4120 26802 4176
rect 26693 4115 26802 4120
rect 2037 4042 2103 4045
rect 6637 4042 6703 4045
rect 2037 4040 6703 4042
rect 2037 3984 2042 4040
rect 2098 3984 6642 4040
rect 6698 3984 6703 4040
rect 2037 3982 6703 3984
rect 2037 3979 2103 3982
rect 6637 3979 6703 3982
rect 20621 4042 20687 4045
rect 23841 4042 23907 4045
rect 20621 4040 23907 4042
rect 20621 3984 20626 4040
rect 20682 3984 23846 4040
rect 23902 3984 23907 4040
rect 20621 3982 23907 3984
rect 20621 3979 20687 3982
rect 23841 3979 23907 3982
rect 0 3906 480 3936
rect 1577 3906 1643 3909
rect 0 3904 1643 3906
rect 0 3848 1582 3904
rect 1638 3848 1643 3904
rect 0 3846 1643 3848
rect 0 3816 480 3846
rect 1577 3843 1643 3846
rect 22001 3906 22067 3909
rect 26601 3906 26667 3909
rect 22001 3904 26667 3906
rect 22001 3848 22006 3904
rect 22062 3848 26606 3904
rect 26662 3848 26667 3904
rect 22001 3846 26667 3848
rect 26742 3906 26802 4115
rect 26877 4042 26943 4045
rect 27613 4042 27679 4045
rect 26877 4040 27679 4042
rect 26877 3984 26882 4040
rect 26938 3984 27618 4040
rect 27674 3984 27679 4040
rect 26877 3982 27679 3984
rect 26877 3979 26943 3982
rect 27613 3979 27679 3982
rect 29520 3906 30000 3936
rect 26742 3846 30000 3906
rect 22001 3843 22067 3846
rect 26601 3843 26667 3846
rect 10944 3840 11264 3841
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 3775 11264 3776
rect 20944 3840 21264 3841
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 29520 3816 30000 3846
rect 20944 3775 21264 3776
rect 24853 3770 24919 3773
rect 27061 3770 27127 3773
rect 24853 3768 27127 3770
rect 24853 3712 24858 3768
rect 24914 3712 27066 3768
rect 27122 3712 27127 3768
rect 24853 3710 27127 3712
rect 24853 3707 24919 3710
rect 27061 3707 27127 3710
rect 657 3634 723 3637
rect 9397 3634 9463 3637
rect 657 3632 9463 3634
rect 657 3576 662 3632
rect 718 3576 9402 3632
rect 9458 3576 9463 3632
rect 657 3574 9463 3576
rect 657 3571 723 3574
rect 9397 3571 9463 3574
rect 2497 3498 2563 3501
rect 12525 3498 12591 3501
rect 2497 3496 12591 3498
rect 2497 3440 2502 3496
rect 2558 3440 12530 3496
rect 12586 3440 12591 3496
rect 2497 3438 12591 3440
rect 2497 3435 2563 3438
rect 12525 3435 12591 3438
rect 25497 3498 25563 3501
rect 25497 3496 27538 3498
rect 25497 3440 25502 3496
rect 25558 3440 27538 3496
rect 25497 3438 27538 3440
rect 25497 3435 25563 3438
rect 0 3362 480 3392
rect 2773 3362 2839 3365
rect 0 3360 2839 3362
rect 0 3304 2778 3360
rect 2834 3304 2839 3360
rect 0 3302 2839 3304
rect 27478 3362 27538 3438
rect 29520 3362 30000 3392
rect 27478 3302 30000 3362
rect 0 3272 480 3302
rect 2773 3299 2839 3302
rect 5944 3296 6264 3297
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 3231 6264 3232
rect 15944 3296 16264 3297
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 3231 16264 3232
rect 25944 3296 26264 3297
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 29520 3272 30000 3302
rect 25944 3231 26264 3232
rect 18781 3226 18847 3229
rect 19977 3226 20043 3229
rect 18781 3224 25882 3226
rect 18781 3168 18786 3224
rect 18842 3168 19982 3224
rect 20038 3168 25882 3224
rect 18781 3166 25882 3168
rect 18781 3163 18847 3166
rect 19977 3163 20043 3166
rect 9857 3090 9923 3093
rect 25313 3090 25379 3093
rect 9857 3088 25379 3090
rect 9857 3032 9862 3088
rect 9918 3032 25318 3088
rect 25374 3032 25379 3088
rect 9857 3030 25379 3032
rect 25822 3090 25882 3166
rect 26417 3090 26483 3093
rect 25822 3088 26483 3090
rect 25822 3032 26422 3088
rect 26478 3032 26483 3088
rect 25822 3030 26483 3032
rect 9857 3027 9923 3030
rect 25313 3027 25379 3030
rect 26417 3027 26483 3030
rect 5717 2954 5783 2957
rect 9213 2954 9279 2957
rect 5717 2952 9279 2954
rect 5717 2896 5722 2952
rect 5778 2896 9218 2952
rect 9274 2896 9279 2952
rect 5717 2894 9279 2896
rect 5717 2891 5783 2894
rect 9213 2891 9279 2894
rect 9397 2954 9463 2957
rect 23841 2954 23907 2957
rect 9397 2952 23907 2954
rect 9397 2896 9402 2952
rect 9458 2896 23846 2952
rect 23902 2896 23907 2952
rect 9397 2894 23907 2896
rect 9397 2891 9463 2894
rect 23841 2891 23907 2894
rect 4061 2818 4127 2821
rect 6821 2818 6887 2821
rect 4061 2816 6887 2818
rect 4061 2760 4066 2816
rect 4122 2760 6826 2816
rect 6882 2760 6887 2816
rect 4061 2758 6887 2760
rect 4061 2755 4127 2758
rect 6821 2755 6887 2758
rect 19149 2818 19215 2821
rect 20621 2818 20687 2821
rect 19149 2816 20687 2818
rect 19149 2760 19154 2816
rect 19210 2760 20626 2816
rect 20682 2760 20687 2816
rect 19149 2758 20687 2760
rect 19149 2755 19215 2758
rect 20621 2755 20687 2758
rect 27705 2818 27771 2821
rect 27705 2816 27906 2818
rect 27705 2760 27710 2816
rect 27766 2760 27906 2816
rect 27705 2758 27906 2760
rect 27705 2755 27771 2758
rect 10944 2752 11264 2753
rect 0 2682 480 2712
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2687 11264 2688
rect 20944 2752 21264 2753
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2687 21264 2688
rect 2865 2682 2931 2685
rect 0 2680 2931 2682
rect 0 2624 2870 2680
rect 2926 2624 2931 2680
rect 0 2622 2931 2624
rect 27846 2682 27906 2758
rect 29520 2682 30000 2712
rect 27846 2622 30000 2682
rect 0 2592 480 2622
rect 2865 2619 2931 2622
rect 29520 2592 30000 2622
rect 9765 2546 9831 2549
rect 11053 2546 11119 2549
rect 9765 2544 11119 2546
rect 9765 2488 9770 2544
rect 9826 2488 11058 2544
rect 11114 2488 11119 2544
rect 9765 2486 11119 2488
rect 9765 2483 9831 2486
rect 11053 2483 11119 2486
rect 5944 2208 6264 2209
rect 0 2138 480 2168
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2143 6264 2144
rect 15944 2208 16264 2209
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2143 16264 2144
rect 25944 2208 26264 2209
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2143 26264 2144
rect 2773 2138 2839 2141
rect 0 2136 2839 2138
rect 0 2080 2778 2136
rect 2834 2080 2839 2136
rect 0 2078 2839 2080
rect 0 2048 480 2078
rect 2773 2075 2839 2078
rect 26693 2138 26759 2141
rect 29520 2138 30000 2168
rect 26693 2136 30000 2138
rect 26693 2080 26698 2136
rect 26754 2080 30000 2136
rect 26693 2078 30000 2080
rect 26693 2075 26759 2078
rect 29520 2048 30000 2078
rect 0 1458 480 1488
rect 1577 1458 1643 1461
rect 0 1456 1643 1458
rect 0 1400 1582 1456
rect 1638 1400 1643 1456
rect 0 1398 1643 1400
rect 0 1368 480 1398
rect 1577 1395 1643 1398
rect 6361 1458 6427 1461
rect 9949 1458 10015 1461
rect 6361 1456 10015 1458
rect 6361 1400 6366 1456
rect 6422 1400 9954 1456
rect 10010 1400 10015 1456
rect 6361 1398 10015 1400
rect 6361 1395 6427 1398
rect 9949 1395 10015 1398
rect 22001 1458 22067 1461
rect 24209 1458 24275 1461
rect 22001 1456 24275 1458
rect 22001 1400 22006 1456
rect 22062 1400 24214 1456
rect 24270 1400 24275 1456
rect 22001 1398 24275 1400
rect 22001 1395 22067 1398
rect 24209 1395 24275 1398
rect 25865 1458 25931 1461
rect 29520 1458 30000 1488
rect 25865 1456 30000 1458
rect 25865 1400 25870 1456
rect 25926 1400 30000 1456
rect 25865 1398 30000 1400
rect 25865 1395 25931 1398
rect 29520 1368 30000 1398
rect 0 914 480 944
rect 3969 914 4035 917
rect 0 912 4035 914
rect 0 856 3974 912
rect 4030 856 4035 912
rect 0 854 4035 856
rect 0 824 480 854
rect 3969 851 4035 854
rect 26601 914 26667 917
rect 29520 914 30000 944
rect 26601 912 30000 914
rect 26601 856 26606 912
rect 26662 856 30000 912
rect 26601 854 30000 856
rect 26601 851 26667 854
rect 29520 824 30000 854
rect 0 370 480 400
rect 1393 370 1459 373
rect 0 368 1459 370
rect 0 312 1398 368
rect 1454 312 1459 368
rect 0 310 1459 312
rect 0 280 480 310
rect 1393 307 1459 310
rect 26785 370 26851 373
rect 29520 370 30000 400
rect 26785 368 30000 370
rect 26785 312 26790 368
rect 26846 312 30000 368
rect 26785 310 30000 312
rect 26785 307 26851 310
rect 29520 280 30000 310
<< via3 >>
rect 5952 21788 6016 21792
rect 5952 21732 5956 21788
rect 5956 21732 6012 21788
rect 6012 21732 6016 21788
rect 5952 21728 6016 21732
rect 6032 21788 6096 21792
rect 6032 21732 6036 21788
rect 6036 21732 6092 21788
rect 6092 21732 6096 21788
rect 6032 21728 6096 21732
rect 6112 21788 6176 21792
rect 6112 21732 6116 21788
rect 6116 21732 6172 21788
rect 6172 21732 6176 21788
rect 6112 21728 6176 21732
rect 6192 21788 6256 21792
rect 6192 21732 6196 21788
rect 6196 21732 6252 21788
rect 6252 21732 6256 21788
rect 6192 21728 6256 21732
rect 15952 21788 16016 21792
rect 15952 21732 15956 21788
rect 15956 21732 16012 21788
rect 16012 21732 16016 21788
rect 15952 21728 16016 21732
rect 16032 21788 16096 21792
rect 16032 21732 16036 21788
rect 16036 21732 16092 21788
rect 16092 21732 16096 21788
rect 16032 21728 16096 21732
rect 16112 21788 16176 21792
rect 16112 21732 16116 21788
rect 16116 21732 16172 21788
rect 16172 21732 16176 21788
rect 16112 21728 16176 21732
rect 16192 21788 16256 21792
rect 16192 21732 16196 21788
rect 16196 21732 16252 21788
rect 16252 21732 16256 21788
rect 16192 21728 16256 21732
rect 25952 21788 26016 21792
rect 25952 21732 25956 21788
rect 25956 21732 26012 21788
rect 26012 21732 26016 21788
rect 25952 21728 26016 21732
rect 26032 21788 26096 21792
rect 26032 21732 26036 21788
rect 26036 21732 26092 21788
rect 26092 21732 26096 21788
rect 26032 21728 26096 21732
rect 26112 21788 26176 21792
rect 26112 21732 26116 21788
rect 26116 21732 26172 21788
rect 26172 21732 26176 21788
rect 26112 21728 26176 21732
rect 26192 21788 26256 21792
rect 26192 21732 26196 21788
rect 26196 21732 26252 21788
rect 26252 21732 26256 21788
rect 26192 21728 26256 21732
rect 10952 21244 11016 21248
rect 10952 21188 10956 21244
rect 10956 21188 11012 21244
rect 11012 21188 11016 21244
rect 10952 21184 11016 21188
rect 11032 21244 11096 21248
rect 11032 21188 11036 21244
rect 11036 21188 11092 21244
rect 11092 21188 11096 21244
rect 11032 21184 11096 21188
rect 11112 21244 11176 21248
rect 11112 21188 11116 21244
rect 11116 21188 11172 21244
rect 11172 21188 11176 21244
rect 11112 21184 11176 21188
rect 11192 21244 11256 21248
rect 11192 21188 11196 21244
rect 11196 21188 11252 21244
rect 11252 21188 11256 21244
rect 11192 21184 11256 21188
rect 20952 21244 21016 21248
rect 20952 21188 20956 21244
rect 20956 21188 21012 21244
rect 21012 21188 21016 21244
rect 20952 21184 21016 21188
rect 21032 21244 21096 21248
rect 21032 21188 21036 21244
rect 21036 21188 21092 21244
rect 21092 21188 21096 21244
rect 21032 21184 21096 21188
rect 21112 21244 21176 21248
rect 21112 21188 21116 21244
rect 21116 21188 21172 21244
rect 21172 21188 21176 21244
rect 21112 21184 21176 21188
rect 21192 21244 21256 21248
rect 21192 21188 21196 21244
rect 21196 21188 21252 21244
rect 21252 21188 21256 21244
rect 21192 21184 21256 21188
rect 5952 20700 6016 20704
rect 5952 20644 5956 20700
rect 5956 20644 6012 20700
rect 6012 20644 6016 20700
rect 5952 20640 6016 20644
rect 6032 20700 6096 20704
rect 6032 20644 6036 20700
rect 6036 20644 6092 20700
rect 6092 20644 6096 20700
rect 6032 20640 6096 20644
rect 6112 20700 6176 20704
rect 6112 20644 6116 20700
rect 6116 20644 6172 20700
rect 6172 20644 6176 20700
rect 6112 20640 6176 20644
rect 6192 20700 6256 20704
rect 6192 20644 6196 20700
rect 6196 20644 6252 20700
rect 6252 20644 6256 20700
rect 6192 20640 6256 20644
rect 15952 20700 16016 20704
rect 15952 20644 15956 20700
rect 15956 20644 16012 20700
rect 16012 20644 16016 20700
rect 15952 20640 16016 20644
rect 16032 20700 16096 20704
rect 16032 20644 16036 20700
rect 16036 20644 16092 20700
rect 16092 20644 16096 20700
rect 16032 20640 16096 20644
rect 16112 20700 16176 20704
rect 16112 20644 16116 20700
rect 16116 20644 16172 20700
rect 16172 20644 16176 20700
rect 16112 20640 16176 20644
rect 16192 20700 16256 20704
rect 16192 20644 16196 20700
rect 16196 20644 16252 20700
rect 16252 20644 16256 20700
rect 16192 20640 16256 20644
rect 25952 20700 26016 20704
rect 25952 20644 25956 20700
rect 25956 20644 26012 20700
rect 26012 20644 26016 20700
rect 25952 20640 26016 20644
rect 26032 20700 26096 20704
rect 26032 20644 26036 20700
rect 26036 20644 26092 20700
rect 26092 20644 26096 20700
rect 26032 20640 26096 20644
rect 26112 20700 26176 20704
rect 26112 20644 26116 20700
rect 26116 20644 26172 20700
rect 26172 20644 26176 20700
rect 26112 20640 26176 20644
rect 26192 20700 26256 20704
rect 26192 20644 26196 20700
rect 26196 20644 26252 20700
rect 26252 20644 26256 20700
rect 26192 20640 26256 20644
rect 10952 20156 11016 20160
rect 10952 20100 10956 20156
rect 10956 20100 11012 20156
rect 11012 20100 11016 20156
rect 10952 20096 11016 20100
rect 11032 20156 11096 20160
rect 11032 20100 11036 20156
rect 11036 20100 11092 20156
rect 11092 20100 11096 20156
rect 11032 20096 11096 20100
rect 11112 20156 11176 20160
rect 11112 20100 11116 20156
rect 11116 20100 11172 20156
rect 11172 20100 11176 20156
rect 11112 20096 11176 20100
rect 11192 20156 11256 20160
rect 11192 20100 11196 20156
rect 11196 20100 11252 20156
rect 11252 20100 11256 20156
rect 11192 20096 11256 20100
rect 20952 20156 21016 20160
rect 20952 20100 20956 20156
rect 20956 20100 21012 20156
rect 21012 20100 21016 20156
rect 20952 20096 21016 20100
rect 21032 20156 21096 20160
rect 21032 20100 21036 20156
rect 21036 20100 21092 20156
rect 21092 20100 21096 20156
rect 21032 20096 21096 20100
rect 21112 20156 21176 20160
rect 21112 20100 21116 20156
rect 21116 20100 21172 20156
rect 21172 20100 21176 20156
rect 21112 20096 21176 20100
rect 21192 20156 21256 20160
rect 21192 20100 21196 20156
rect 21196 20100 21252 20156
rect 21252 20100 21256 20156
rect 21192 20096 21256 20100
rect 5952 19612 6016 19616
rect 5952 19556 5956 19612
rect 5956 19556 6012 19612
rect 6012 19556 6016 19612
rect 5952 19552 6016 19556
rect 6032 19612 6096 19616
rect 6032 19556 6036 19612
rect 6036 19556 6092 19612
rect 6092 19556 6096 19612
rect 6032 19552 6096 19556
rect 6112 19612 6176 19616
rect 6112 19556 6116 19612
rect 6116 19556 6172 19612
rect 6172 19556 6176 19612
rect 6112 19552 6176 19556
rect 6192 19612 6256 19616
rect 6192 19556 6196 19612
rect 6196 19556 6252 19612
rect 6252 19556 6256 19612
rect 6192 19552 6256 19556
rect 15952 19612 16016 19616
rect 15952 19556 15956 19612
rect 15956 19556 16012 19612
rect 16012 19556 16016 19612
rect 15952 19552 16016 19556
rect 16032 19612 16096 19616
rect 16032 19556 16036 19612
rect 16036 19556 16092 19612
rect 16092 19556 16096 19612
rect 16032 19552 16096 19556
rect 16112 19612 16176 19616
rect 16112 19556 16116 19612
rect 16116 19556 16172 19612
rect 16172 19556 16176 19612
rect 16112 19552 16176 19556
rect 16192 19612 16256 19616
rect 16192 19556 16196 19612
rect 16196 19556 16252 19612
rect 16252 19556 16256 19612
rect 16192 19552 16256 19556
rect 25952 19612 26016 19616
rect 25952 19556 25956 19612
rect 25956 19556 26012 19612
rect 26012 19556 26016 19612
rect 25952 19552 26016 19556
rect 26032 19612 26096 19616
rect 26032 19556 26036 19612
rect 26036 19556 26092 19612
rect 26092 19556 26096 19612
rect 26032 19552 26096 19556
rect 26112 19612 26176 19616
rect 26112 19556 26116 19612
rect 26116 19556 26172 19612
rect 26172 19556 26176 19612
rect 26112 19552 26176 19556
rect 26192 19612 26256 19616
rect 26192 19556 26196 19612
rect 26196 19556 26252 19612
rect 26252 19556 26256 19612
rect 26192 19552 26256 19556
rect 10952 19068 11016 19072
rect 10952 19012 10956 19068
rect 10956 19012 11012 19068
rect 11012 19012 11016 19068
rect 10952 19008 11016 19012
rect 11032 19068 11096 19072
rect 11032 19012 11036 19068
rect 11036 19012 11092 19068
rect 11092 19012 11096 19068
rect 11032 19008 11096 19012
rect 11112 19068 11176 19072
rect 11112 19012 11116 19068
rect 11116 19012 11172 19068
rect 11172 19012 11176 19068
rect 11112 19008 11176 19012
rect 11192 19068 11256 19072
rect 11192 19012 11196 19068
rect 11196 19012 11252 19068
rect 11252 19012 11256 19068
rect 11192 19008 11256 19012
rect 20952 19068 21016 19072
rect 20952 19012 20956 19068
rect 20956 19012 21012 19068
rect 21012 19012 21016 19068
rect 20952 19008 21016 19012
rect 21032 19068 21096 19072
rect 21032 19012 21036 19068
rect 21036 19012 21092 19068
rect 21092 19012 21096 19068
rect 21032 19008 21096 19012
rect 21112 19068 21176 19072
rect 21112 19012 21116 19068
rect 21116 19012 21172 19068
rect 21172 19012 21176 19068
rect 21112 19008 21176 19012
rect 21192 19068 21256 19072
rect 21192 19012 21196 19068
rect 21196 19012 21252 19068
rect 21252 19012 21256 19068
rect 21192 19008 21256 19012
rect 5952 18524 6016 18528
rect 5952 18468 5956 18524
rect 5956 18468 6012 18524
rect 6012 18468 6016 18524
rect 5952 18464 6016 18468
rect 6032 18524 6096 18528
rect 6032 18468 6036 18524
rect 6036 18468 6092 18524
rect 6092 18468 6096 18524
rect 6032 18464 6096 18468
rect 6112 18524 6176 18528
rect 6112 18468 6116 18524
rect 6116 18468 6172 18524
rect 6172 18468 6176 18524
rect 6112 18464 6176 18468
rect 6192 18524 6256 18528
rect 6192 18468 6196 18524
rect 6196 18468 6252 18524
rect 6252 18468 6256 18524
rect 6192 18464 6256 18468
rect 15952 18524 16016 18528
rect 15952 18468 15956 18524
rect 15956 18468 16012 18524
rect 16012 18468 16016 18524
rect 15952 18464 16016 18468
rect 16032 18524 16096 18528
rect 16032 18468 16036 18524
rect 16036 18468 16092 18524
rect 16092 18468 16096 18524
rect 16032 18464 16096 18468
rect 16112 18524 16176 18528
rect 16112 18468 16116 18524
rect 16116 18468 16172 18524
rect 16172 18468 16176 18524
rect 16112 18464 16176 18468
rect 16192 18524 16256 18528
rect 16192 18468 16196 18524
rect 16196 18468 16252 18524
rect 16252 18468 16256 18524
rect 16192 18464 16256 18468
rect 25952 18524 26016 18528
rect 25952 18468 25956 18524
rect 25956 18468 26012 18524
rect 26012 18468 26016 18524
rect 25952 18464 26016 18468
rect 26032 18524 26096 18528
rect 26032 18468 26036 18524
rect 26036 18468 26092 18524
rect 26092 18468 26096 18524
rect 26032 18464 26096 18468
rect 26112 18524 26176 18528
rect 26112 18468 26116 18524
rect 26116 18468 26172 18524
rect 26172 18468 26176 18524
rect 26112 18464 26176 18468
rect 26192 18524 26256 18528
rect 26192 18468 26196 18524
rect 26196 18468 26252 18524
rect 26252 18468 26256 18524
rect 26192 18464 26256 18468
rect 10952 17980 11016 17984
rect 10952 17924 10956 17980
rect 10956 17924 11012 17980
rect 11012 17924 11016 17980
rect 10952 17920 11016 17924
rect 11032 17980 11096 17984
rect 11032 17924 11036 17980
rect 11036 17924 11092 17980
rect 11092 17924 11096 17980
rect 11032 17920 11096 17924
rect 11112 17980 11176 17984
rect 11112 17924 11116 17980
rect 11116 17924 11172 17980
rect 11172 17924 11176 17980
rect 11112 17920 11176 17924
rect 11192 17980 11256 17984
rect 11192 17924 11196 17980
rect 11196 17924 11252 17980
rect 11252 17924 11256 17980
rect 11192 17920 11256 17924
rect 20952 17980 21016 17984
rect 20952 17924 20956 17980
rect 20956 17924 21012 17980
rect 21012 17924 21016 17980
rect 20952 17920 21016 17924
rect 21032 17980 21096 17984
rect 21032 17924 21036 17980
rect 21036 17924 21092 17980
rect 21092 17924 21096 17980
rect 21032 17920 21096 17924
rect 21112 17980 21176 17984
rect 21112 17924 21116 17980
rect 21116 17924 21172 17980
rect 21172 17924 21176 17980
rect 21112 17920 21176 17924
rect 21192 17980 21256 17984
rect 21192 17924 21196 17980
rect 21196 17924 21252 17980
rect 21252 17924 21256 17980
rect 21192 17920 21256 17924
rect 5952 17436 6016 17440
rect 5952 17380 5956 17436
rect 5956 17380 6012 17436
rect 6012 17380 6016 17436
rect 5952 17376 6016 17380
rect 6032 17436 6096 17440
rect 6032 17380 6036 17436
rect 6036 17380 6092 17436
rect 6092 17380 6096 17436
rect 6032 17376 6096 17380
rect 6112 17436 6176 17440
rect 6112 17380 6116 17436
rect 6116 17380 6172 17436
rect 6172 17380 6176 17436
rect 6112 17376 6176 17380
rect 6192 17436 6256 17440
rect 6192 17380 6196 17436
rect 6196 17380 6252 17436
rect 6252 17380 6256 17436
rect 6192 17376 6256 17380
rect 15952 17436 16016 17440
rect 15952 17380 15956 17436
rect 15956 17380 16012 17436
rect 16012 17380 16016 17436
rect 15952 17376 16016 17380
rect 16032 17436 16096 17440
rect 16032 17380 16036 17436
rect 16036 17380 16092 17436
rect 16092 17380 16096 17436
rect 16032 17376 16096 17380
rect 16112 17436 16176 17440
rect 16112 17380 16116 17436
rect 16116 17380 16172 17436
rect 16172 17380 16176 17436
rect 16112 17376 16176 17380
rect 16192 17436 16256 17440
rect 16192 17380 16196 17436
rect 16196 17380 16252 17436
rect 16252 17380 16256 17436
rect 16192 17376 16256 17380
rect 25952 17436 26016 17440
rect 25952 17380 25956 17436
rect 25956 17380 26012 17436
rect 26012 17380 26016 17436
rect 25952 17376 26016 17380
rect 26032 17436 26096 17440
rect 26032 17380 26036 17436
rect 26036 17380 26092 17436
rect 26092 17380 26096 17436
rect 26032 17376 26096 17380
rect 26112 17436 26176 17440
rect 26112 17380 26116 17436
rect 26116 17380 26172 17436
rect 26172 17380 26176 17436
rect 26112 17376 26176 17380
rect 26192 17436 26256 17440
rect 26192 17380 26196 17436
rect 26196 17380 26252 17436
rect 26252 17380 26256 17436
rect 26192 17376 26256 17380
rect 10952 16892 11016 16896
rect 10952 16836 10956 16892
rect 10956 16836 11012 16892
rect 11012 16836 11016 16892
rect 10952 16832 11016 16836
rect 11032 16892 11096 16896
rect 11032 16836 11036 16892
rect 11036 16836 11092 16892
rect 11092 16836 11096 16892
rect 11032 16832 11096 16836
rect 11112 16892 11176 16896
rect 11112 16836 11116 16892
rect 11116 16836 11172 16892
rect 11172 16836 11176 16892
rect 11112 16832 11176 16836
rect 11192 16892 11256 16896
rect 11192 16836 11196 16892
rect 11196 16836 11252 16892
rect 11252 16836 11256 16892
rect 11192 16832 11256 16836
rect 20952 16892 21016 16896
rect 20952 16836 20956 16892
rect 20956 16836 21012 16892
rect 21012 16836 21016 16892
rect 20952 16832 21016 16836
rect 21032 16892 21096 16896
rect 21032 16836 21036 16892
rect 21036 16836 21092 16892
rect 21092 16836 21096 16892
rect 21032 16832 21096 16836
rect 21112 16892 21176 16896
rect 21112 16836 21116 16892
rect 21116 16836 21172 16892
rect 21172 16836 21176 16892
rect 21112 16832 21176 16836
rect 21192 16892 21256 16896
rect 21192 16836 21196 16892
rect 21196 16836 21252 16892
rect 21252 16836 21256 16892
rect 21192 16832 21256 16836
rect 5952 16348 6016 16352
rect 5952 16292 5956 16348
rect 5956 16292 6012 16348
rect 6012 16292 6016 16348
rect 5952 16288 6016 16292
rect 6032 16348 6096 16352
rect 6032 16292 6036 16348
rect 6036 16292 6092 16348
rect 6092 16292 6096 16348
rect 6032 16288 6096 16292
rect 6112 16348 6176 16352
rect 6112 16292 6116 16348
rect 6116 16292 6172 16348
rect 6172 16292 6176 16348
rect 6112 16288 6176 16292
rect 6192 16348 6256 16352
rect 6192 16292 6196 16348
rect 6196 16292 6252 16348
rect 6252 16292 6256 16348
rect 6192 16288 6256 16292
rect 15952 16348 16016 16352
rect 15952 16292 15956 16348
rect 15956 16292 16012 16348
rect 16012 16292 16016 16348
rect 15952 16288 16016 16292
rect 16032 16348 16096 16352
rect 16032 16292 16036 16348
rect 16036 16292 16092 16348
rect 16092 16292 16096 16348
rect 16032 16288 16096 16292
rect 16112 16348 16176 16352
rect 16112 16292 16116 16348
rect 16116 16292 16172 16348
rect 16172 16292 16176 16348
rect 16112 16288 16176 16292
rect 16192 16348 16256 16352
rect 16192 16292 16196 16348
rect 16196 16292 16252 16348
rect 16252 16292 16256 16348
rect 16192 16288 16256 16292
rect 25952 16348 26016 16352
rect 25952 16292 25956 16348
rect 25956 16292 26012 16348
rect 26012 16292 26016 16348
rect 25952 16288 26016 16292
rect 26032 16348 26096 16352
rect 26032 16292 26036 16348
rect 26036 16292 26092 16348
rect 26092 16292 26096 16348
rect 26032 16288 26096 16292
rect 26112 16348 26176 16352
rect 26112 16292 26116 16348
rect 26116 16292 26172 16348
rect 26172 16292 26176 16348
rect 26112 16288 26176 16292
rect 26192 16348 26256 16352
rect 26192 16292 26196 16348
rect 26196 16292 26252 16348
rect 26252 16292 26256 16348
rect 26192 16288 26256 16292
rect 10952 15804 11016 15808
rect 10952 15748 10956 15804
rect 10956 15748 11012 15804
rect 11012 15748 11016 15804
rect 10952 15744 11016 15748
rect 11032 15804 11096 15808
rect 11032 15748 11036 15804
rect 11036 15748 11092 15804
rect 11092 15748 11096 15804
rect 11032 15744 11096 15748
rect 11112 15804 11176 15808
rect 11112 15748 11116 15804
rect 11116 15748 11172 15804
rect 11172 15748 11176 15804
rect 11112 15744 11176 15748
rect 11192 15804 11256 15808
rect 11192 15748 11196 15804
rect 11196 15748 11252 15804
rect 11252 15748 11256 15804
rect 11192 15744 11256 15748
rect 20952 15804 21016 15808
rect 20952 15748 20956 15804
rect 20956 15748 21012 15804
rect 21012 15748 21016 15804
rect 20952 15744 21016 15748
rect 21032 15804 21096 15808
rect 21032 15748 21036 15804
rect 21036 15748 21092 15804
rect 21092 15748 21096 15804
rect 21032 15744 21096 15748
rect 21112 15804 21176 15808
rect 21112 15748 21116 15804
rect 21116 15748 21172 15804
rect 21172 15748 21176 15804
rect 21112 15744 21176 15748
rect 21192 15804 21256 15808
rect 21192 15748 21196 15804
rect 21196 15748 21252 15804
rect 21252 15748 21256 15804
rect 21192 15744 21256 15748
rect 25636 15540 25700 15604
rect 5952 15260 6016 15264
rect 5952 15204 5956 15260
rect 5956 15204 6012 15260
rect 6012 15204 6016 15260
rect 5952 15200 6016 15204
rect 6032 15260 6096 15264
rect 6032 15204 6036 15260
rect 6036 15204 6092 15260
rect 6092 15204 6096 15260
rect 6032 15200 6096 15204
rect 6112 15260 6176 15264
rect 6112 15204 6116 15260
rect 6116 15204 6172 15260
rect 6172 15204 6176 15260
rect 6112 15200 6176 15204
rect 6192 15260 6256 15264
rect 6192 15204 6196 15260
rect 6196 15204 6252 15260
rect 6252 15204 6256 15260
rect 6192 15200 6256 15204
rect 15952 15260 16016 15264
rect 15952 15204 15956 15260
rect 15956 15204 16012 15260
rect 16012 15204 16016 15260
rect 15952 15200 16016 15204
rect 16032 15260 16096 15264
rect 16032 15204 16036 15260
rect 16036 15204 16092 15260
rect 16092 15204 16096 15260
rect 16032 15200 16096 15204
rect 16112 15260 16176 15264
rect 16112 15204 16116 15260
rect 16116 15204 16172 15260
rect 16172 15204 16176 15260
rect 16112 15200 16176 15204
rect 16192 15260 16256 15264
rect 16192 15204 16196 15260
rect 16196 15204 16252 15260
rect 16252 15204 16256 15260
rect 16192 15200 16256 15204
rect 25952 15260 26016 15264
rect 25952 15204 25956 15260
rect 25956 15204 26012 15260
rect 26012 15204 26016 15260
rect 25952 15200 26016 15204
rect 26032 15260 26096 15264
rect 26032 15204 26036 15260
rect 26036 15204 26092 15260
rect 26092 15204 26096 15260
rect 26032 15200 26096 15204
rect 26112 15260 26176 15264
rect 26112 15204 26116 15260
rect 26116 15204 26172 15260
rect 26172 15204 26176 15260
rect 26112 15200 26176 15204
rect 26192 15260 26256 15264
rect 26192 15204 26196 15260
rect 26196 15204 26252 15260
rect 26252 15204 26256 15260
rect 26192 15200 26256 15204
rect 25084 14920 25148 14924
rect 25084 14864 25098 14920
rect 25098 14864 25148 14920
rect 25084 14860 25148 14864
rect 10952 14716 11016 14720
rect 10952 14660 10956 14716
rect 10956 14660 11012 14716
rect 11012 14660 11016 14716
rect 10952 14656 11016 14660
rect 11032 14716 11096 14720
rect 11032 14660 11036 14716
rect 11036 14660 11092 14716
rect 11092 14660 11096 14716
rect 11032 14656 11096 14660
rect 11112 14716 11176 14720
rect 11112 14660 11116 14716
rect 11116 14660 11172 14716
rect 11172 14660 11176 14716
rect 11112 14656 11176 14660
rect 11192 14716 11256 14720
rect 11192 14660 11196 14716
rect 11196 14660 11252 14716
rect 11252 14660 11256 14716
rect 11192 14656 11256 14660
rect 20952 14716 21016 14720
rect 20952 14660 20956 14716
rect 20956 14660 21012 14716
rect 21012 14660 21016 14716
rect 20952 14656 21016 14660
rect 21032 14716 21096 14720
rect 21032 14660 21036 14716
rect 21036 14660 21092 14716
rect 21092 14660 21096 14716
rect 21032 14656 21096 14660
rect 21112 14716 21176 14720
rect 21112 14660 21116 14716
rect 21116 14660 21172 14716
rect 21172 14660 21176 14716
rect 21112 14656 21176 14660
rect 21192 14716 21256 14720
rect 21192 14660 21196 14716
rect 21196 14660 21252 14716
rect 21252 14660 21256 14716
rect 21192 14656 21256 14660
rect 5952 14172 6016 14176
rect 5952 14116 5956 14172
rect 5956 14116 6012 14172
rect 6012 14116 6016 14172
rect 5952 14112 6016 14116
rect 6032 14172 6096 14176
rect 6032 14116 6036 14172
rect 6036 14116 6092 14172
rect 6092 14116 6096 14172
rect 6032 14112 6096 14116
rect 6112 14172 6176 14176
rect 6112 14116 6116 14172
rect 6116 14116 6172 14172
rect 6172 14116 6176 14172
rect 6112 14112 6176 14116
rect 6192 14172 6256 14176
rect 6192 14116 6196 14172
rect 6196 14116 6252 14172
rect 6252 14116 6256 14172
rect 6192 14112 6256 14116
rect 15952 14172 16016 14176
rect 15952 14116 15956 14172
rect 15956 14116 16012 14172
rect 16012 14116 16016 14172
rect 15952 14112 16016 14116
rect 16032 14172 16096 14176
rect 16032 14116 16036 14172
rect 16036 14116 16092 14172
rect 16092 14116 16096 14172
rect 16032 14112 16096 14116
rect 16112 14172 16176 14176
rect 16112 14116 16116 14172
rect 16116 14116 16172 14172
rect 16172 14116 16176 14172
rect 16112 14112 16176 14116
rect 16192 14172 16256 14176
rect 16192 14116 16196 14172
rect 16196 14116 16252 14172
rect 16252 14116 16256 14172
rect 16192 14112 16256 14116
rect 25952 14172 26016 14176
rect 25952 14116 25956 14172
rect 25956 14116 26012 14172
rect 26012 14116 26016 14172
rect 25952 14112 26016 14116
rect 26032 14172 26096 14176
rect 26032 14116 26036 14172
rect 26036 14116 26092 14172
rect 26092 14116 26096 14172
rect 26032 14112 26096 14116
rect 26112 14172 26176 14176
rect 26112 14116 26116 14172
rect 26116 14116 26172 14172
rect 26172 14116 26176 14172
rect 26112 14112 26176 14116
rect 26192 14172 26256 14176
rect 26192 14116 26196 14172
rect 26196 14116 26252 14172
rect 26252 14116 26256 14172
rect 26192 14112 26256 14116
rect 10952 13628 11016 13632
rect 10952 13572 10956 13628
rect 10956 13572 11012 13628
rect 11012 13572 11016 13628
rect 10952 13568 11016 13572
rect 11032 13628 11096 13632
rect 11032 13572 11036 13628
rect 11036 13572 11092 13628
rect 11092 13572 11096 13628
rect 11032 13568 11096 13572
rect 11112 13628 11176 13632
rect 11112 13572 11116 13628
rect 11116 13572 11172 13628
rect 11172 13572 11176 13628
rect 11112 13568 11176 13572
rect 11192 13628 11256 13632
rect 11192 13572 11196 13628
rect 11196 13572 11252 13628
rect 11252 13572 11256 13628
rect 11192 13568 11256 13572
rect 20952 13628 21016 13632
rect 20952 13572 20956 13628
rect 20956 13572 21012 13628
rect 21012 13572 21016 13628
rect 20952 13568 21016 13572
rect 21032 13628 21096 13632
rect 21032 13572 21036 13628
rect 21036 13572 21092 13628
rect 21092 13572 21096 13628
rect 21032 13568 21096 13572
rect 21112 13628 21176 13632
rect 21112 13572 21116 13628
rect 21116 13572 21172 13628
rect 21172 13572 21176 13628
rect 21112 13568 21176 13572
rect 21192 13628 21256 13632
rect 21192 13572 21196 13628
rect 21196 13572 21252 13628
rect 21252 13572 21256 13628
rect 21192 13568 21256 13572
rect 5952 13084 6016 13088
rect 5952 13028 5956 13084
rect 5956 13028 6012 13084
rect 6012 13028 6016 13084
rect 5952 13024 6016 13028
rect 6032 13084 6096 13088
rect 6032 13028 6036 13084
rect 6036 13028 6092 13084
rect 6092 13028 6096 13084
rect 6032 13024 6096 13028
rect 6112 13084 6176 13088
rect 6112 13028 6116 13084
rect 6116 13028 6172 13084
rect 6172 13028 6176 13084
rect 6112 13024 6176 13028
rect 6192 13084 6256 13088
rect 6192 13028 6196 13084
rect 6196 13028 6252 13084
rect 6252 13028 6256 13084
rect 6192 13024 6256 13028
rect 15952 13084 16016 13088
rect 15952 13028 15956 13084
rect 15956 13028 16012 13084
rect 16012 13028 16016 13084
rect 15952 13024 16016 13028
rect 16032 13084 16096 13088
rect 16032 13028 16036 13084
rect 16036 13028 16092 13084
rect 16092 13028 16096 13084
rect 16032 13024 16096 13028
rect 16112 13084 16176 13088
rect 16112 13028 16116 13084
rect 16116 13028 16172 13084
rect 16172 13028 16176 13084
rect 16112 13024 16176 13028
rect 16192 13084 16256 13088
rect 16192 13028 16196 13084
rect 16196 13028 16252 13084
rect 16252 13028 16256 13084
rect 16192 13024 16256 13028
rect 25952 13084 26016 13088
rect 25952 13028 25956 13084
rect 25956 13028 26012 13084
rect 26012 13028 26016 13084
rect 25952 13024 26016 13028
rect 26032 13084 26096 13088
rect 26032 13028 26036 13084
rect 26036 13028 26092 13084
rect 26092 13028 26096 13084
rect 26032 13024 26096 13028
rect 26112 13084 26176 13088
rect 26112 13028 26116 13084
rect 26116 13028 26172 13084
rect 26172 13028 26176 13084
rect 26112 13024 26176 13028
rect 26192 13084 26256 13088
rect 26192 13028 26196 13084
rect 26196 13028 26252 13084
rect 26252 13028 26256 13084
rect 26192 13024 26256 13028
rect 19012 12820 19076 12884
rect 19196 12820 19260 12884
rect 10952 12540 11016 12544
rect 10952 12484 10956 12540
rect 10956 12484 11012 12540
rect 11012 12484 11016 12540
rect 10952 12480 11016 12484
rect 11032 12540 11096 12544
rect 11032 12484 11036 12540
rect 11036 12484 11092 12540
rect 11092 12484 11096 12540
rect 11032 12480 11096 12484
rect 11112 12540 11176 12544
rect 11112 12484 11116 12540
rect 11116 12484 11172 12540
rect 11172 12484 11176 12540
rect 11112 12480 11176 12484
rect 11192 12540 11256 12544
rect 11192 12484 11196 12540
rect 11196 12484 11252 12540
rect 11252 12484 11256 12540
rect 11192 12480 11256 12484
rect 20952 12540 21016 12544
rect 20952 12484 20956 12540
rect 20956 12484 21012 12540
rect 21012 12484 21016 12540
rect 20952 12480 21016 12484
rect 21032 12540 21096 12544
rect 21032 12484 21036 12540
rect 21036 12484 21092 12540
rect 21092 12484 21096 12540
rect 21032 12480 21096 12484
rect 21112 12540 21176 12544
rect 21112 12484 21116 12540
rect 21116 12484 21172 12540
rect 21172 12484 21176 12540
rect 21112 12480 21176 12484
rect 21192 12540 21256 12544
rect 21192 12484 21196 12540
rect 21196 12484 21252 12540
rect 21252 12484 21256 12540
rect 21192 12480 21256 12484
rect 25084 12064 25148 12068
rect 25084 12008 25098 12064
rect 25098 12008 25148 12064
rect 25084 12004 25148 12008
rect 5952 11996 6016 12000
rect 5952 11940 5956 11996
rect 5956 11940 6012 11996
rect 6012 11940 6016 11996
rect 5952 11936 6016 11940
rect 6032 11996 6096 12000
rect 6032 11940 6036 11996
rect 6036 11940 6092 11996
rect 6092 11940 6096 11996
rect 6032 11936 6096 11940
rect 6112 11996 6176 12000
rect 6112 11940 6116 11996
rect 6116 11940 6172 11996
rect 6172 11940 6176 11996
rect 6112 11936 6176 11940
rect 6192 11996 6256 12000
rect 6192 11940 6196 11996
rect 6196 11940 6252 11996
rect 6252 11940 6256 11996
rect 6192 11936 6256 11940
rect 15952 11996 16016 12000
rect 15952 11940 15956 11996
rect 15956 11940 16012 11996
rect 16012 11940 16016 11996
rect 15952 11936 16016 11940
rect 16032 11996 16096 12000
rect 16032 11940 16036 11996
rect 16036 11940 16092 11996
rect 16092 11940 16096 11996
rect 16032 11936 16096 11940
rect 16112 11996 16176 12000
rect 16112 11940 16116 11996
rect 16116 11940 16172 11996
rect 16172 11940 16176 11996
rect 16112 11936 16176 11940
rect 16192 11996 16256 12000
rect 16192 11940 16196 11996
rect 16196 11940 16252 11996
rect 16252 11940 16256 11996
rect 16192 11936 16256 11940
rect 25952 11996 26016 12000
rect 25952 11940 25956 11996
rect 25956 11940 26012 11996
rect 26012 11940 26016 11996
rect 25952 11936 26016 11940
rect 26032 11996 26096 12000
rect 26032 11940 26036 11996
rect 26036 11940 26092 11996
rect 26092 11940 26096 11996
rect 26032 11936 26096 11940
rect 26112 11996 26176 12000
rect 26112 11940 26116 11996
rect 26116 11940 26172 11996
rect 26172 11940 26176 11996
rect 26112 11936 26176 11940
rect 26192 11996 26256 12000
rect 26192 11940 26196 11996
rect 26196 11940 26252 11996
rect 26252 11940 26256 11996
rect 26192 11936 26256 11940
rect 25636 11460 25700 11524
rect 10952 11452 11016 11456
rect 10952 11396 10956 11452
rect 10956 11396 11012 11452
rect 11012 11396 11016 11452
rect 10952 11392 11016 11396
rect 11032 11452 11096 11456
rect 11032 11396 11036 11452
rect 11036 11396 11092 11452
rect 11092 11396 11096 11452
rect 11032 11392 11096 11396
rect 11112 11452 11176 11456
rect 11112 11396 11116 11452
rect 11116 11396 11172 11452
rect 11172 11396 11176 11452
rect 11112 11392 11176 11396
rect 11192 11452 11256 11456
rect 11192 11396 11196 11452
rect 11196 11396 11252 11452
rect 11252 11396 11256 11452
rect 11192 11392 11256 11396
rect 20952 11452 21016 11456
rect 20952 11396 20956 11452
rect 20956 11396 21012 11452
rect 21012 11396 21016 11452
rect 20952 11392 21016 11396
rect 21032 11452 21096 11456
rect 21032 11396 21036 11452
rect 21036 11396 21092 11452
rect 21092 11396 21096 11452
rect 21032 11392 21096 11396
rect 21112 11452 21176 11456
rect 21112 11396 21116 11452
rect 21116 11396 21172 11452
rect 21172 11396 21176 11452
rect 21112 11392 21176 11396
rect 21192 11452 21256 11456
rect 21192 11396 21196 11452
rect 21196 11396 21252 11452
rect 21252 11396 21256 11452
rect 21192 11392 21256 11396
rect 5952 10908 6016 10912
rect 5952 10852 5956 10908
rect 5956 10852 6012 10908
rect 6012 10852 6016 10908
rect 5952 10848 6016 10852
rect 6032 10908 6096 10912
rect 6032 10852 6036 10908
rect 6036 10852 6092 10908
rect 6092 10852 6096 10908
rect 6032 10848 6096 10852
rect 6112 10908 6176 10912
rect 6112 10852 6116 10908
rect 6116 10852 6172 10908
rect 6172 10852 6176 10908
rect 6112 10848 6176 10852
rect 6192 10908 6256 10912
rect 6192 10852 6196 10908
rect 6196 10852 6252 10908
rect 6252 10852 6256 10908
rect 6192 10848 6256 10852
rect 15952 10908 16016 10912
rect 15952 10852 15956 10908
rect 15956 10852 16012 10908
rect 16012 10852 16016 10908
rect 15952 10848 16016 10852
rect 16032 10908 16096 10912
rect 16032 10852 16036 10908
rect 16036 10852 16092 10908
rect 16092 10852 16096 10908
rect 16032 10848 16096 10852
rect 16112 10908 16176 10912
rect 16112 10852 16116 10908
rect 16116 10852 16172 10908
rect 16172 10852 16176 10908
rect 16112 10848 16176 10852
rect 16192 10908 16256 10912
rect 16192 10852 16196 10908
rect 16196 10852 16252 10908
rect 16252 10852 16256 10908
rect 16192 10848 16256 10852
rect 25952 10908 26016 10912
rect 25952 10852 25956 10908
rect 25956 10852 26012 10908
rect 26012 10852 26016 10908
rect 25952 10848 26016 10852
rect 26032 10908 26096 10912
rect 26032 10852 26036 10908
rect 26036 10852 26092 10908
rect 26092 10852 26096 10908
rect 26032 10848 26096 10852
rect 26112 10908 26176 10912
rect 26112 10852 26116 10908
rect 26116 10852 26172 10908
rect 26172 10852 26176 10908
rect 26112 10848 26176 10852
rect 26192 10908 26256 10912
rect 26192 10852 26196 10908
rect 26196 10852 26252 10908
rect 26252 10852 26256 10908
rect 26192 10848 26256 10852
rect 10952 10364 11016 10368
rect 10952 10308 10956 10364
rect 10956 10308 11012 10364
rect 11012 10308 11016 10364
rect 10952 10304 11016 10308
rect 11032 10364 11096 10368
rect 11032 10308 11036 10364
rect 11036 10308 11092 10364
rect 11092 10308 11096 10364
rect 11032 10304 11096 10308
rect 11112 10364 11176 10368
rect 11112 10308 11116 10364
rect 11116 10308 11172 10364
rect 11172 10308 11176 10364
rect 11112 10304 11176 10308
rect 11192 10364 11256 10368
rect 11192 10308 11196 10364
rect 11196 10308 11252 10364
rect 11252 10308 11256 10364
rect 11192 10304 11256 10308
rect 20952 10364 21016 10368
rect 20952 10308 20956 10364
rect 20956 10308 21012 10364
rect 21012 10308 21016 10364
rect 20952 10304 21016 10308
rect 21032 10364 21096 10368
rect 21032 10308 21036 10364
rect 21036 10308 21092 10364
rect 21092 10308 21096 10364
rect 21032 10304 21096 10308
rect 21112 10364 21176 10368
rect 21112 10308 21116 10364
rect 21116 10308 21172 10364
rect 21172 10308 21176 10364
rect 21112 10304 21176 10308
rect 21192 10364 21256 10368
rect 21192 10308 21196 10364
rect 21196 10308 21252 10364
rect 21252 10308 21256 10364
rect 21192 10304 21256 10308
rect 19012 10296 19076 10300
rect 19012 10240 19062 10296
rect 19062 10240 19076 10296
rect 19012 10236 19076 10240
rect 5952 9820 6016 9824
rect 5952 9764 5956 9820
rect 5956 9764 6012 9820
rect 6012 9764 6016 9820
rect 5952 9760 6016 9764
rect 6032 9820 6096 9824
rect 6032 9764 6036 9820
rect 6036 9764 6092 9820
rect 6092 9764 6096 9820
rect 6032 9760 6096 9764
rect 6112 9820 6176 9824
rect 6112 9764 6116 9820
rect 6116 9764 6172 9820
rect 6172 9764 6176 9820
rect 6112 9760 6176 9764
rect 6192 9820 6256 9824
rect 6192 9764 6196 9820
rect 6196 9764 6252 9820
rect 6252 9764 6256 9820
rect 6192 9760 6256 9764
rect 15952 9820 16016 9824
rect 15952 9764 15956 9820
rect 15956 9764 16012 9820
rect 16012 9764 16016 9820
rect 15952 9760 16016 9764
rect 16032 9820 16096 9824
rect 16032 9764 16036 9820
rect 16036 9764 16092 9820
rect 16092 9764 16096 9820
rect 16032 9760 16096 9764
rect 16112 9820 16176 9824
rect 16112 9764 16116 9820
rect 16116 9764 16172 9820
rect 16172 9764 16176 9820
rect 16112 9760 16176 9764
rect 16192 9820 16256 9824
rect 16192 9764 16196 9820
rect 16196 9764 16252 9820
rect 16252 9764 16256 9820
rect 16192 9760 16256 9764
rect 25952 9820 26016 9824
rect 25952 9764 25956 9820
rect 25956 9764 26012 9820
rect 26012 9764 26016 9820
rect 25952 9760 26016 9764
rect 26032 9820 26096 9824
rect 26032 9764 26036 9820
rect 26036 9764 26092 9820
rect 26092 9764 26096 9820
rect 26032 9760 26096 9764
rect 26112 9820 26176 9824
rect 26112 9764 26116 9820
rect 26116 9764 26172 9820
rect 26172 9764 26176 9820
rect 26112 9760 26176 9764
rect 26192 9820 26256 9824
rect 26192 9764 26196 9820
rect 26196 9764 26252 9820
rect 26252 9764 26256 9820
rect 26192 9760 26256 9764
rect 10952 9276 11016 9280
rect 10952 9220 10956 9276
rect 10956 9220 11012 9276
rect 11012 9220 11016 9276
rect 10952 9216 11016 9220
rect 11032 9276 11096 9280
rect 11032 9220 11036 9276
rect 11036 9220 11092 9276
rect 11092 9220 11096 9276
rect 11032 9216 11096 9220
rect 11112 9276 11176 9280
rect 11112 9220 11116 9276
rect 11116 9220 11172 9276
rect 11172 9220 11176 9276
rect 11112 9216 11176 9220
rect 11192 9276 11256 9280
rect 11192 9220 11196 9276
rect 11196 9220 11252 9276
rect 11252 9220 11256 9276
rect 11192 9216 11256 9220
rect 20952 9276 21016 9280
rect 20952 9220 20956 9276
rect 20956 9220 21012 9276
rect 21012 9220 21016 9276
rect 20952 9216 21016 9220
rect 21032 9276 21096 9280
rect 21032 9220 21036 9276
rect 21036 9220 21092 9276
rect 21092 9220 21096 9276
rect 21032 9216 21096 9220
rect 21112 9276 21176 9280
rect 21112 9220 21116 9276
rect 21116 9220 21172 9276
rect 21172 9220 21176 9276
rect 21112 9216 21176 9220
rect 21192 9276 21256 9280
rect 21192 9220 21196 9276
rect 21196 9220 21252 9276
rect 21252 9220 21256 9276
rect 21192 9216 21256 9220
rect 5952 8732 6016 8736
rect 5952 8676 5956 8732
rect 5956 8676 6012 8732
rect 6012 8676 6016 8732
rect 5952 8672 6016 8676
rect 6032 8732 6096 8736
rect 6032 8676 6036 8732
rect 6036 8676 6092 8732
rect 6092 8676 6096 8732
rect 6032 8672 6096 8676
rect 6112 8732 6176 8736
rect 6112 8676 6116 8732
rect 6116 8676 6172 8732
rect 6172 8676 6176 8732
rect 6112 8672 6176 8676
rect 6192 8732 6256 8736
rect 6192 8676 6196 8732
rect 6196 8676 6252 8732
rect 6252 8676 6256 8732
rect 6192 8672 6256 8676
rect 15952 8732 16016 8736
rect 15952 8676 15956 8732
rect 15956 8676 16012 8732
rect 16012 8676 16016 8732
rect 15952 8672 16016 8676
rect 16032 8732 16096 8736
rect 16032 8676 16036 8732
rect 16036 8676 16092 8732
rect 16092 8676 16096 8732
rect 16032 8672 16096 8676
rect 16112 8732 16176 8736
rect 16112 8676 16116 8732
rect 16116 8676 16172 8732
rect 16172 8676 16176 8732
rect 16112 8672 16176 8676
rect 16192 8732 16256 8736
rect 16192 8676 16196 8732
rect 16196 8676 16252 8732
rect 16252 8676 16256 8732
rect 16192 8672 16256 8676
rect 25952 8732 26016 8736
rect 25952 8676 25956 8732
rect 25956 8676 26012 8732
rect 26012 8676 26016 8732
rect 25952 8672 26016 8676
rect 26032 8732 26096 8736
rect 26032 8676 26036 8732
rect 26036 8676 26092 8732
rect 26092 8676 26096 8732
rect 26032 8672 26096 8676
rect 26112 8732 26176 8736
rect 26112 8676 26116 8732
rect 26116 8676 26172 8732
rect 26172 8676 26176 8732
rect 26112 8672 26176 8676
rect 26192 8732 26256 8736
rect 26192 8676 26196 8732
rect 26196 8676 26252 8732
rect 26252 8676 26256 8732
rect 26192 8672 26256 8676
rect 10952 8188 11016 8192
rect 10952 8132 10956 8188
rect 10956 8132 11012 8188
rect 11012 8132 11016 8188
rect 10952 8128 11016 8132
rect 11032 8188 11096 8192
rect 11032 8132 11036 8188
rect 11036 8132 11092 8188
rect 11092 8132 11096 8188
rect 11032 8128 11096 8132
rect 11112 8188 11176 8192
rect 11112 8132 11116 8188
rect 11116 8132 11172 8188
rect 11172 8132 11176 8188
rect 11112 8128 11176 8132
rect 11192 8188 11256 8192
rect 11192 8132 11196 8188
rect 11196 8132 11252 8188
rect 11252 8132 11256 8188
rect 11192 8128 11256 8132
rect 20952 8188 21016 8192
rect 20952 8132 20956 8188
rect 20956 8132 21012 8188
rect 21012 8132 21016 8188
rect 20952 8128 21016 8132
rect 21032 8188 21096 8192
rect 21032 8132 21036 8188
rect 21036 8132 21092 8188
rect 21092 8132 21096 8188
rect 21032 8128 21096 8132
rect 21112 8188 21176 8192
rect 21112 8132 21116 8188
rect 21116 8132 21172 8188
rect 21172 8132 21176 8188
rect 21112 8128 21176 8132
rect 21192 8188 21256 8192
rect 21192 8132 21196 8188
rect 21196 8132 21252 8188
rect 21252 8132 21256 8188
rect 21192 8128 21256 8132
rect 5952 7644 6016 7648
rect 5952 7588 5956 7644
rect 5956 7588 6012 7644
rect 6012 7588 6016 7644
rect 5952 7584 6016 7588
rect 6032 7644 6096 7648
rect 6032 7588 6036 7644
rect 6036 7588 6092 7644
rect 6092 7588 6096 7644
rect 6032 7584 6096 7588
rect 6112 7644 6176 7648
rect 6112 7588 6116 7644
rect 6116 7588 6172 7644
rect 6172 7588 6176 7644
rect 6112 7584 6176 7588
rect 6192 7644 6256 7648
rect 6192 7588 6196 7644
rect 6196 7588 6252 7644
rect 6252 7588 6256 7644
rect 6192 7584 6256 7588
rect 15952 7644 16016 7648
rect 15952 7588 15956 7644
rect 15956 7588 16012 7644
rect 16012 7588 16016 7644
rect 15952 7584 16016 7588
rect 16032 7644 16096 7648
rect 16032 7588 16036 7644
rect 16036 7588 16092 7644
rect 16092 7588 16096 7644
rect 16032 7584 16096 7588
rect 16112 7644 16176 7648
rect 16112 7588 16116 7644
rect 16116 7588 16172 7644
rect 16172 7588 16176 7644
rect 16112 7584 16176 7588
rect 16192 7644 16256 7648
rect 16192 7588 16196 7644
rect 16196 7588 16252 7644
rect 16252 7588 16256 7644
rect 16192 7584 16256 7588
rect 25952 7644 26016 7648
rect 25952 7588 25956 7644
rect 25956 7588 26012 7644
rect 26012 7588 26016 7644
rect 25952 7584 26016 7588
rect 26032 7644 26096 7648
rect 26032 7588 26036 7644
rect 26036 7588 26092 7644
rect 26092 7588 26096 7644
rect 26032 7584 26096 7588
rect 26112 7644 26176 7648
rect 26112 7588 26116 7644
rect 26116 7588 26172 7644
rect 26172 7588 26176 7644
rect 26112 7584 26176 7588
rect 26192 7644 26256 7648
rect 26192 7588 26196 7644
rect 26196 7588 26252 7644
rect 26252 7588 26256 7644
rect 26192 7584 26256 7588
rect 10952 7100 11016 7104
rect 10952 7044 10956 7100
rect 10956 7044 11012 7100
rect 11012 7044 11016 7100
rect 10952 7040 11016 7044
rect 11032 7100 11096 7104
rect 11032 7044 11036 7100
rect 11036 7044 11092 7100
rect 11092 7044 11096 7100
rect 11032 7040 11096 7044
rect 11112 7100 11176 7104
rect 11112 7044 11116 7100
rect 11116 7044 11172 7100
rect 11172 7044 11176 7100
rect 11112 7040 11176 7044
rect 11192 7100 11256 7104
rect 11192 7044 11196 7100
rect 11196 7044 11252 7100
rect 11252 7044 11256 7100
rect 11192 7040 11256 7044
rect 20952 7100 21016 7104
rect 20952 7044 20956 7100
rect 20956 7044 21012 7100
rect 21012 7044 21016 7100
rect 20952 7040 21016 7044
rect 21032 7100 21096 7104
rect 21032 7044 21036 7100
rect 21036 7044 21092 7100
rect 21092 7044 21096 7100
rect 21032 7040 21096 7044
rect 21112 7100 21176 7104
rect 21112 7044 21116 7100
rect 21116 7044 21172 7100
rect 21172 7044 21176 7100
rect 21112 7040 21176 7044
rect 21192 7100 21256 7104
rect 21192 7044 21196 7100
rect 21196 7044 21252 7100
rect 21252 7044 21256 7100
rect 21192 7040 21256 7044
rect 5952 6556 6016 6560
rect 5952 6500 5956 6556
rect 5956 6500 6012 6556
rect 6012 6500 6016 6556
rect 5952 6496 6016 6500
rect 6032 6556 6096 6560
rect 6032 6500 6036 6556
rect 6036 6500 6092 6556
rect 6092 6500 6096 6556
rect 6032 6496 6096 6500
rect 6112 6556 6176 6560
rect 6112 6500 6116 6556
rect 6116 6500 6172 6556
rect 6172 6500 6176 6556
rect 6112 6496 6176 6500
rect 6192 6556 6256 6560
rect 6192 6500 6196 6556
rect 6196 6500 6252 6556
rect 6252 6500 6256 6556
rect 6192 6496 6256 6500
rect 15952 6556 16016 6560
rect 15952 6500 15956 6556
rect 15956 6500 16012 6556
rect 16012 6500 16016 6556
rect 15952 6496 16016 6500
rect 16032 6556 16096 6560
rect 16032 6500 16036 6556
rect 16036 6500 16092 6556
rect 16092 6500 16096 6556
rect 16032 6496 16096 6500
rect 16112 6556 16176 6560
rect 16112 6500 16116 6556
rect 16116 6500 16172 6556
rect 16172 6500 16176 6556
rect 16112 6496 16176 6500
rect 16192 6556 16256 6560
rect 16192 6500 16196 6556
rect 16196 6500 16252 6556
rect 16252 6500 16256 6556
rect 16192 6496 16256 6500
rect 25952 6556 26016 6560
rect 25952 6500 25956 6556
rect 25956 6500 26012 6556
rect 26012 6500 26016 6556
rect 25952 6496 26016 6500
rect 26032 6556 26096 6560
rect 26032 6500 26036 6556
rect 26036 6500 26092 6556
rect 26092 6500 26096 6556
rect 26032 6496 26096 6500
rect 26112 6556 26176 6560
rect 26112 6500 26116 6556
rect 26116 6500 26172 6556
rect 26172 6500 26176 6556
rect 26112 6496 26176 6500
rect 26192 6556 26256 6560
rect 26192 6500 26196 6556
rect 26196 6500 26252 6556
rect 26252 6500 26256 6556
rect 26192 6496 26256 6500
rect 10952 6012 11016 6016
rect 10952 5956 10956 6012
rect 10956 5956 11012 6012
rect 11012 5956 11016 6012
rect 10952 5952 11016 5956
rect 11032 6012 11096 6016
rect 11032 5956 11036 6012
rect 11036 5956 11092 6012
rect 11092 5956 11096 6012
rect 11032 5952 11096 5956
rect 11112 6012 11176 6016
rect 11112 5956 11116 6012
rect 11116 5956 11172 6012
rect 11172 5956 11176 6012
rect 11112 5952 11176 5956
rect 11192 6012 11256 6016
rect 11192 5956 11196 6012
rect 11196 5956 11252 6012
rect 11252 5956 11256 6012
rect 11192 5952 11256 5956
rect 20952 6012 21016 6016
rect 20952 5956 20956 6012
rect 20956 5956 21012 6012
rect 21012 5956 21016 6012
rect 20952 5952 21016 5956
rect 21032 6012 21096 6016
rect 21032 5956 21036 6012
rect 21036 5956 21092 6012
rect 21092 5956 21096 6012
rect 21032 5952 21096 5956
rect 21112 6012 21176 6016
rect 21112 5956 21116 6012
rect 21116 5956 21172 6012
rect 21172 5956 21176 6012
rect 21112 5952 21176 5956
rect 21192 6012 21256 6016
rect 21192 5956 21196 6012
rect 21196 5956 21252 6012
rect 21252 5956 21256 6012
rect 21192 5952 21256 5956
rect 5952 5468 6016 5472
rect 5952 5412 5956 5468
rect 5956 5412 6012 5468
rect 6012 5412 6016 5468
rect 5952 5408 6016 5412
rect 6032 5468 6096 5472
rect 6032 5412 6036 5468
rect 6036 5412 6092 5468
rect 6092 5412 6096 5468
rect 6032 5408 6096 5412
rect 6112 5468 6176 5472
rect 6112 5412 6116 5468
rect 6116 5412 6172 5468
rect 6172 5412 6176 5468
rect 6112 5408 6176 5412
rect 6192 5468 6256 5472
rect 6192 5412 6196 5468
rect 6196 5412 6252 5468
rect 6252 5412 6256 5468
rect 6192 5408 6256 5412
rect 15952 5468 16016 5472
rect 15952 5412 15956 5468
rect 15956 5412 16012 5468
rect 16012 5412 16016 5468
rect 15952 5408 16016 5412
rect 16032 5468 16096 5472
rect 16032 5412 16036 5468
rect 16036 5412 16092 5468
rect 16092 5412 16096 5468
rect 16032 5408 16096 5412
rect 16112 5468 16176 5472
rect 16112 5412 16116 5468
rect 16116 5412 16172 5468
rect 16172 5412 16176 5468
rect 16112 5408 16176 5412
rect 16192 5468 16256 5472
rect 16192 5412 16196 5468
rect 16196 5412 16252 5468
rect 16252 5412 16256 5468
rect 16192 5408 16256 5412
rect 25952 5468 26016 5472
rect 25952 5412 25956 5468
rect 25956 5412 26012 5468
rect 26012 5412 26016 5468
rect 25952 5408 26016 5412
rect 26032 5468 26096 5472
rect 26032 5412 26036 5468
rect 26036 5412 26092 5468
rect 26092 5412 26096 5468
rect 26032 5408 26096 5412
rect 26112 5468 26176 5472
rect 26112 5412 26116 5468
rect 26116 5412 26172 5468
rect 26172 5412 26176 5468
rect 26112 5408 26176 5412
rect 26192 5468 26256 5472
rect 26192 5412 26196 5468
rect 26196 5412 26252 5468
rect 26252 5412 26256 5468
rect 26192 5408 26256 5412
rect 10952 4924 11016 4928
rect 10952 4868 10956 4924
rect 10956 4868 11012 4924
rect 11012 4868 11016 4924
rect 10952 4864 11016 4868
rect 11032 4924 11096 4928
rect 11032 4868 11036 4924
rect 11036 4868 11092 4924
rect 11092 4868 11096 4924
rect 11032 4864 11096 4868
rect 11112 4924 11176 4928
rect 11112 4868 11116 4924
rect 11116 4868 11172 4924
rect 11172 4868 11176 4924
rect 11112 4864 11176 4868
rect 11192 4924 11256 4928
rect 11192 4868 11196 4924
rect 11196 4868 11252 4924
rect 11252 4868 11256 4924
rect 11192 4864 11256 4868
rect 20952 4924 21016 4928
rect 20952 4868 20956 4924
rect 20956 4868 21012 4924
rect 21012 4868 21016 4924
rect 20952 4864 21016 4868
rect 21032 4924 21096 4928
rect 21032 4868 21036 4924
rect 21036 4868 21092 4924
rect 21092 4868 21096 4924
rect 21032 4864 21096 4868
rect 21112 4924 21176 4928
rect 21112 4868 21116 4924
rect 21116 4868 21172 4924
rect 21172 4868 21176 4924
rect 21112 4864 21176 4868
rect 21192 4924 21256 4928
rect 21192 4868 21196 4924
rect 21196 4868 21252 4924
rect 21252 4868 21256 4924
rect 21192 4864 21256 4868
rect 5952 4380 6016 4384
rect 5952 4324 5956 4380
rect 5956 4324 6012 4380
rect 6012 4324 6016 4380
rect 5952 4320 6016 4324
rect 6032 4380 6096 4384
rect 6032 4324 6036 4380
rect 6036 4324 6092 4380
rect 6092 4324 6096 4380
rect 6032 4320 6096 4324
rect 6112 4380 6176 4384
rect 6112 4324 6116 4380
rect 6116 4324 6172 4380
rect 6172 4324 6176 4380
rect 6112 4320 6176 4324
rect 6192 4380 6256 4384
rect 6192 4324 6196 4380
rect 6196 4324 6252 4380
rect 6252 4324 6256 4380
rect 6192 4320 6256 4324
rect 15952 4380 16016 4384
rect 15952 4324 15956 4380
rect 15956 4324 16012 4380
rect 16012 4324 16016 4380
rect 15952 4320 16016 4324
rect 16032 4380 16096 4384
rect 16032 4324 16036 4380
rect 16036 4324 16092 4380
rect 16092 4324 16096 4380
rect 16032 4320 16096 4324
rect 16112 4380 16176 4384
rect 16112 4324 16116 4380
rect 16116 4324 16172 4380
rect 16172 4324 16176 4380
rect 16112 4320 16176 4324
rect 16192 4380 16256 4384
rect 16192 4324 16196 4380
rect 16196 4324 16252 4380
rect 16252 4324 16256 4380
rect 16192 4320 16256 4324
rect 25952 4380 26016 4384
rect 25952 4324 25956 4380
rect 25956 4324 26012 4380
rect 26012 4324 26016 4380
rect 25952 4320 26016 4324
rect 26032 4380 26096 4384
rect 26032 4324 26036 4380
rect 26036 4324 26092 4380
rect 26092 4324 26096 4380
rect 26032 4320 26096 4324
rect 26112 4380 26176 4384
rect 26112 4324 26116 4380
rect 26116 4324 26172 4380
rect 26172 4324 26176 4380
rect 26112 4320 26176 4324
rect 26192 4380 26256 4384
rect 26192 4324 26196 4380
rect 26196 4324 26252 4380
rect 26252 4324 26256 4380
rect 26192 4320 26256 4324
rect 10952 3836 11016 3840
rect 10952 3780 10956 3836
rect 10956 3780 11012 3836
rect 11012 3780 11016 3836
rect 10952 3776 11016 3780
rect 11032 3836 11096 3840
rect 11032 3780 11036 3836
rect 11036 3780 11092 3836
rect 11092 3780 11096 3836
rect 11032 3776 11096 3780
rect 11112 3836 11176 3840
rect 11112 3780 11116 3836
rect 11116 3780 11172 3836
rect 11172 3780 11176 3836
rect 11112 3776 11176 3780
rect 11192 3836 11256 3840
rect 11192 3780 11196 3836
rect 11196 3780 11252 3836
rect 11252 3780 11256 3836
rect 11192 3776 11256 3780
rect 20952 3836 21016 3840
rect 20952 3780 20956 3836
rect 20956 3780 21012 3836
rect 21012 3780 21016 3836
rect 20952 3776 21016 3780
rect 21032 3836 21096 3840
rect 21032 3780 21036 3836
rect 21036 3780 21092 3836
rect 21092 3780 21096 3836
rect 21032 3776 21096 3780
rect 21112 3836 21176 3840
rect 21112 3780 21116 3836
rect 21116 3780 21172 3836
rect 21172 3780 21176 3836
rect 21112 3776 21176 3780
rect 21192 3836 21256 3840
rect 21192 3780 21196 3836
rect 21196 3780 21252 3836
rect 21252 3780 21256 3836
rect 21192 3776 21256 3780
rect 5952 3292 6016 3296
rect 5952 3236 5956 3292
rect 5956 3236 6012 3292
rect 6012 3236 6016 3292
rect 5952 3232 6016 3236
rect 6032 3292 6096 3296
rect 6032 3236 6036 3292
rect 6036 3236 6092 3292
rect 6092 3236 6096 3292
rect 6032 3232 6096 3236
rect 6112 3292 6176 3296
rect 6112 3236 6116 3292
rect 6116 3236 6172 3292
rect 6172 3236 6176 3292
rect 6112 3232 6176 3236
rect 6192 3292 6256 3296
rect 6192 3236 6196 3292
rect 6196 3236 6252 3292
rect 6252 3236 6256 3292
rect 6192 3232 6256 3236
rect 15952 3292 16016 3296
rect 15952 3236 15956 3292
rect 15956 3236 16012 3292
rect 16012 3236 16016 3292
rect 15952 3232 16016 3236
rect 16032 3292 16096 3296
rect 16032 3236 16036 3292
rect 16036 3236 16092 3292
rect 16092 3236 16096 3292
rect 16032 3232 16096 3236
rect 16112 3292 16176 3296
rect 16112 3236 16116 3292
rect 16116 3236 16172 3292
rect 16172 3236 16176 3292
rect 16112 3232 16176 3236
rect 16192 3292 16256 3296
rect 16192 3236 16196 3292
rect 16196 3236 16252 3292
rect 16252 3236 16256 3292
rect 16192 3232 16256 3236
rect 25952 3292 26016 3296
rect 25952 3236 25956 3292
rect 25956 3236 26012 3292
rect 26012 3236 26016 3292
rect 25952 3232 26016 3236
rect 26032 3292 26096 3296
rect 26032 3236 26036 3292
rect 26036 3236 26092 3292
rect 26092 3236 26096 3292
rect 26032 3232 26096 3236
rect 26112 3292 26176 3296
rect 26112 3236 26116 3292
rect 26116 3236 26172 3292
rect 26172 3236 26176 3292
rect 26112 3232 26176 3236
rect 26192 3292 26256 3296
rect 26192 3236 26196 3292
rect 26196 3236 26252 3292
rect 26252 3236 26256 3292
rect 26192 3232 26256 3236
rect 10952 2748 11016 2752
rect 10952 2692 10956 2748
rect 10956 2692 11012 2748
rect 11012 2692 11016 2748
rect 10952 2688 11016 2692
rect 11032 2748 11096 2752
rect 11032 2692 11036 2748
rect 11036 2692 11092 2748
rect 11092 2692 11096 2748
rect 11032 2688 11096 2692
rect 11112 2748 11176 2752
rect 11112 2692 11116 2748
rect 11116 2692 11172 2748
rect 11172 2692 11176 2748
rect 11112 2688 11176 2692
rect 11192 2748 11256 2752
rect 11192 2692 11196 2748
rect 11196 2692 11252 2748
rect 11252 2692 11256 2748
rect 11192 2688 11256 2692
rect 20952 2748 21016 2752
rect 20952 2692 20956 2748
rect 20956 2692 21012 2748
rect 21012 2692 21016 2748
rect 20952 2688 21016 2692
rect 21032 2748 21096 2752
rect 21032 2692 21036 2748
rect 21036 2692 21092 2748
rect 21092 2692 21096 2748
rect 21032 2688 21096 2692
rect 21112 2748 21176 2752
rect 21112 2692 21116 2748
rect 21116 2692 21172 2748
rect 21172 2692 21176 2748
rect 21112 2688 21176 2692
rect 21192 2748 21256 2752
rect 21192 2692 21196 2748
rect 21196 2692 21252 2748
rect 21252 2692 21256 2748
rect 21192 2688 21256 2692
rect 5952 2204 6016 2208
rect 5952 2148 5956 2204
rect 5956 2148 6012 2204
rect 6012 2148 6016 2204
rect 5952 2144 6016 2148
rect 6032 2204 6096 2208
rect 6032 2148 6036 2204
rect 6036 2148 6092 2204
rect 6092 2148 6096 2204
rect 6032 2144 6096 2148
rect 6112 2204 6176 2208
rect 6112 2148 6116 2204
rect 6116 2148 6172 2204
rect 6172 2148 6176 2204
rect 6112 2144 6176 2148
rect 6192 2204 6256 2208
rect 6192 2148 6196 2204
rect 6196 2148 6252 2204
rect 6252 2148 6256 2204
rect 6192 2144 6256 2148
rect 15952 2204 16016 2208
rect 15952 2148 15956 2204
rect 15956 2148 16012 2204
rect 16012 2148 16016 2204
rect 15952 2144 16016 2148
rect 16032 2204 16096 2208
rect 16032 2148 16036 2204
rect 16036 2148 16092 2204
rect 16092 2148 16096 2204
rect 16032 2144 16096 2148
rect 16112 2204 16176 2208
rect 16112 2148 16116 2204
rect 16116 2148 16172 2204
rect 16172 2148 16176 2204
rect 16112 2144 16176 2148
rect 16192 2204 16256 2208
rect 16192 2148 16196 2204
rect 16196 2148 16252 2204
rect 16252 2148 16256 2204
rect 16192 2144 16256 2148
rect 25952 2204 26016 2208
rect 25952 2148 25956 2204
rect 25956 2148 26012 2204
rect 26012 2148 26016 2204
rect 25952 2144 26016 2148
rect 26032 2204 26096 2208
rect 26032 2148 26036 2204
rect 26036 2148 26092 2204
rect 26092 2148 26096 2204
rect 26032 2144 26096 2148
rect 26112 2204 26176 2208
rect 26112 2148 26116 2204
rect 26116 2148 26172 2204
rect 26172 2148 26176 2204
rect 26112 2144 26176 2148
rect 26192 2204 26256 2208
rect 26192 2148 26196 2204
rect 26196 2148 26252 2204
rect 26252 2148 26256 2204
rect 26192 2144 26256 2148
<< metal4 >>
rect 5944 21792 6264 21808
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 20704 6264 21728
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 19616 6264 20640
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 18528 6264 19552
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 17440 6264 18464
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 16352 6264 17376
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 15264 6264 16288
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 14176 6264 15200
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 13088 6264 14112
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 12000 6264 13024
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 10912 6264 11936
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 9824 6264 10848
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 8736 6264 9760
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 7648 6264 8672
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 6560 6264 7584
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 5472 6264 6496
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 4384 6264 5408
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 3296 6264 4320
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 2208 6264 3232
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2128 6264 2144
rect 10944 21248 11264 21808
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 20160 11264 21184
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 19072 11264 20096
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 17984 11264 19008
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 16896 11264 17920
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 15808 11264 16832
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 14720 11264 15744
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 13632 11264 14656
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 12544 11264 13568
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 11456 11264 12480
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 10368 11264 11392
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 9280 11264 10304
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 8192 11264 9216
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 7104 11264 8128
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 6016 11264 7040
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 4928 11264 5952
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 3840 11264 4864
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 2752 11264 3776
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2128 11264 2688
rect 15944 21792 16264 21808
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 20704 16264 21728
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 19616 16264 20640
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 18528 16264 19552
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 17440 16264 18464
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 16352 16264 17376
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 15264 16264 16288
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 14176 16264 15200
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 13088 16264 14112
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 12000 16264 13024
rect 20944 21248 21264 21808
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 20160 21264 21184
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 19072 21264 20096
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 17984 21264 19008
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 16896 21264 17920
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 15808 21264 16832
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 14720 21264 15744
rect 25944 21792 26264 21808
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 20704 26264 21728
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 19616 26264 20640
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 18528 26264 19552
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 17440 26264 18464
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 16352 26264 17376
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25635 15604 25701 15605
rect 25635 15540 25636 15604
rect 25700 15540 25701 15604
rect 25635 15539 25701 15540
rect 25083 14924 25149 14925
rect 25083 14860 25084 14924
rect 25148 14860 25149 14924
rect 25083 14859 25149 14860
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 13632 21264 14656
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 19011 12884 19077 12885
rect 19011 12820 19012 12884
rect 19076 12820 19077 12884
rect 19011 12819 19077 12820
rect 19195 12884 19261 12885
rect 19195 12820 19196 12884
rect 19260 12820 19261 12884
rect 19195 12819 19261 12820
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 10912 16264 11936
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 9824 16264 10848
rect 19014 12610 19074 12819
rect 19198 12610 19258 12819
rect 19014 12550 19258 12610
rect 19014 10301 19074 12550
rect 20944 12544 21264 13568
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 11456 21264 12480
rect 25086 12069 25146 14859
rect 25083 12068 25149 12069
rect 25083 12004 25084 12068
rect 25148 12004 25149 12068
rect 25083 12003 25149 12004
rect 25638 11525 25698 15539
rect 25944 15264 26264 16288
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 14176 26264 15200
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 13088 26264 14112
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 12000 26264 13024
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25635 11524 25701 11525
rect 25635 11460 25636 11524
rect 25700 11460 25701 11524
rect 25635 11459 25701 11460
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 10368 21264 11392
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 19011 10300 19077 10301
rect 19011 10236 19012 10300
rect 19076 10236 19077 10300
rect 19011 10235 19077 10236
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 8736 16264 9760
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 7648 16264 8672
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 6560 16264 7584
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 5472 16264 6496
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 4384 16264 5408
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 3296 16264 4320
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 2208 16264 3232
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2128 16264 2144
rect 20944 9280 21264 10304
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 20944 8192 21264 9216
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 7104 21264 8128
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 6016 21264 7040
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 4928 21264 5952
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 3840 21264 4864
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 2752 21264 3776
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2128 21264 2688
rect 25944 10912 26264 11936
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 9824 26264 10848
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 8736 26264 9760
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 7648 26264 8672
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 6560 26264 7584
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 5472 26264 6496
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 4384 26264 5408
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 3296 26264 4320
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 25944 2208 26264 3232
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2128 26264 2144
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _56_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_13 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9
timestamp 1604681595
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11
timestamp 1604681595
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7
timestamp 1604681595
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2300 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 2668 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1604681595
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_21
timestamp 1604681595
transform 1 0 3036 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21
timestamp 1604681595
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3312 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3864 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_39
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1604681595
transform 1 0 4600 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_45
timestamp 1604681595
transform 1 0 5244 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45
timestamp 1604681595
transform 1 0 5244 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4968 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5428 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5520 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_71
timestamp 1604681595
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1604681595
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_1_83
timestamp 1604681595
transform 1 0 8740 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_79
timestamp 1604681595
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_75
timestamp 1604681595
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_76 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8096 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9200 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10488 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 9200 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_90
timestamp 1604681595
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100
timestamp 1604681595
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104
timestamp 1604681595
transform 1 0 10672 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_111
timestamp 1604681595
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_107
timestamp 1604681595
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11132 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_115 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 11684 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1604681595
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1604681595
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12788 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14352 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13156 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_133
timestamp 1604681595
transform 1 0 13340 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1604681595
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1604681595
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_133 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13340 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_141
timestamp 1604681595
transform 1 0 14076 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_150
timestamp 1604681595
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_166
timestamp 1604681595
transform 1 0 16376 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_164
timestamp 1604681595
transform 1 0 16192 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15640 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_154
timestamp 1604681595
transform 1 0 15272 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_175
timestamp 1604681595
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_168
timestamp 1604681595
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16928 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_179
timestamp 1604681595
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1604681595
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1604681595
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_192
timestamp 1604681595
transform 1 0 18768 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_196
timestamp 1604681595
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_192
timestamp 1604681595
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18584 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18952 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18860 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_203
timestamp 1604681595
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_199
timestamp 1604681595
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19596 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19504 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20148 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1604681595
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1604681595
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_226
timestamp 1604681595
transform 1 0 21896 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_222
timestamp 1604681595
transform 1 0 21528 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21344 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22080 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_236
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_249
timestamp 1604681595
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_242
timestamp 1604681595
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_240
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_230
timestamp 1604681595
transform 1 0 22264 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_253
timestamp 1604681595
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_255
timestamp 1604681595
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604681595
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604681595
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_265
timestamp 1604681595
transform 1 0 25484 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_261
timestamp 1604681595
transform 1 0 25116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_259
timestamp 1604681595
transform 1 0 24932 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 25300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 25668 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_279
timestamp 1604681595
transform 1 0 26772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_273
timestamp 1604681595
transform 1 0 26220 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1604681595
transform 1 0 26404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 1604681595
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 26956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 26404 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604681595
transform 1 0 26864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_291
timestamp 1604681595
transform 1 0 27876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_283
timestamp 1604681595
transform 1 0 27140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 27324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 27508 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_284
timestamp 1604681595
transform 1 0 27232 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 28888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 28060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_296
timestamp 1604681595
transform 1 0 28336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_295
timestamp 1604681595
transform 1 0 28244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604681595
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_7
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_11
timestamp 1604681595
transform 1 0 2116 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_19
timestamp 1604681595
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3036 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_40
timestamp 1604681595
transform 1 0 4784 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_36
timestamp 1604681595
transform 1 0 4416 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5060 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6072 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6440 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_52
timestamp 1604681595
transform 1 0 5888 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_60
timestamp 1604681595
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6992 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_2_73
timestamp 1604681595
transform 1 0 7820 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_85
timestamp 1604681595
transform 1 0 8924 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1604681595
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_2_124
timestamp 1604681595
transform 1 0 12512 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_136
timestamp 1604681595
transform 1 0 13616 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 15916 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1604681595
transform 1 0 14720 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1604681595
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_160
timestamp 1604681595
transform 1 0 15824 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1604681595
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 17204 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_2_167
timestamp 1604681595
transform 1 0 16468 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_194
timestamp 1604681595
transform 1 0 18952 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_199
timestamp 1604681595
transform 1 0 19412 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_207
timestamp 1604681595
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_211
timestamp 1604681595
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_224
timestamp 1604681595
transform 1 0 21712 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_236
timestamp 1604681595
transform 1 0 22816 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_248
timestamp 1604681595
transform 1 0 23920 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_260
timestamp 1604681595
transform 1 0 25024 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_267
timestamp 1604681595
transform 1 0 25668 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_280
timestamp 1604681595
transform 1 0 26864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_292
timestamp 1604681595
transform 1 0 27968 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1604681595
transform 1 0 28520 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 2760 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1604681595
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_11
timestamp 1604681595
transform 1 0 2116 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_17
timestamp 1604681595
transform 1 0 2668 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_37
timestamp 1604681595
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_41
timestamp 1604681595
transform 1 0 4876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 5244 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5060 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_49
timestamp 1604681595
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_53
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_67
timestamp 1604681595
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_71
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_75
timestamp 1604681595
transform 1 0 8004 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_87
timestamp 1604681595
transform 1 0 9108 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_99
timestamp 1604681595
transform 1 0 10212 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1604681595
transform 1 0 11316 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13708 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_131
timestamp 1604681595
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_139
timestamp 1604681595
transform 1 0 13892 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15916 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_151
timestamp 1604681595
transform 1 0 14996 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_157
timestamp 1604681595
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_170
timestamp 1604681595
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_174
timestamp 1604681595
transform 1 0 17112 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1604681595
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19964 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_192
timestamp 1604681595
transform 1 0 18768 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_195
timestamp 1604681595
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_199
timestamp 1604681595
transform 1 0 19412 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21528 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 21344 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_214
timestamp 1604681595
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_218
timestamp 1604681595
transform 1 0 21160 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 23828 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_231
timestamp 1604681595
transform 1 0 22356 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_243
timestamp 1604681595
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_249
timestamp 1604681595
transform 1 0 24012 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 24196 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_253
timestamp 1604681595
transform 1 0 24380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_265
timestamp 1604681595
transform 1 0 25484 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 27324 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 26220 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 26772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 27140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 27876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_277
timestamp 1604681595
transform 1 0 26588 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1604681595
transform 1 0 26956 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_289
timestamp 1604681595
transform 1 0 27692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 28888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1604681595
transform 1 0 28060 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604681595
transform 1 0 1932 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 2300 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_7
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_11
timestamp 1604681595
transform 1 0 2116 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_19
timestamp 1604681595
transform 1 0 2852 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4600 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_57
timestamp 1604681595
transform 1 0 6348 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 7084 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_74
timestamp 1604681595
transform 1 0 7912 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_78
timestamp 1604681595
transform 1 0 8280 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_103
timestamp 1604681595
transform 1 0 10580 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11408 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11132 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_107
timestamp 1604681595
transform 1 0 10948 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_111
timestamp 1604681595
transform 1 0 11316 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_121
timestamp 1604681595
transform 1 0 12236 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_138
timestamp 1604681595
transform 1 0 13800 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 16192 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16008 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp 1604681595
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_183
timestamp 1604681595
transform 1 0 17940 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_195
timestamp 1604681595
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_206
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 21528 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 20516 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_210
timestamp 1604681595
transform 1 0 20424 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1604681595
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_221
timestamp 1604681595
transform 1 0 21436 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_224
timestamp 1604681595
transform 1 0 21712 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 23552 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_4_236
timestamp 1604681595
transform 1 0 22816 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1604681595
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_280
timestamp 1604681595
transform 1 0 26864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 28888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_292
timestamp 1604681595
transform 1 0 27968 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_298
timestamp 1604681595
transform 1 0 28520 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2852 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604681595
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_7
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_11
timestamp 1604681595
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_28
timestamp 1604681595
transform 1 0 3680 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_32
timestamp 1604681595
transform 1 0 4048 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_44
timestamp 1604681595
transform 1 0 5152 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_52
timestamp 1604681595
transform 1 0 5888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604681595
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7084 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8096 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_68
timestamp 1604681595
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_72
timestamp 1604681595
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_95
timestamp 1604681595
transform 1 0 9844 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1604681595
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13248 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 1604681595
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_131
timestamp 1604681595
transform 1 0 13156 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16008 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_151
timestamp 1604681595
transform 1 0 14996 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_155
timestamp 1604681595
transform 1 0 15364 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_158
timestamp 1604681595
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_171
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_179
timestamp 1604681595
transform 1 0 17572 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_192
timestamp 1604681595
transform 1 0 18768 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_195
timestamp 1604681595
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_199
timestamp 1604681595
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_203
timestamp 1604681595
transform 1 0 19780 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_207
timestamp 1604681595
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1604681595
transform 1 0 20516 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_220
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_228
timestamp 1604681595
transform 1 0 22080 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 22724 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_233
timestamp 1604681595
transform 1 0 22540 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_237
timestamp 1604681595
transform 1 0 22908 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_243
timestamp 1604681595
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 25392 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 25208 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_257
timestamp 1604681595
transform 1 0 24748 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_261
timestamp 1604681595
transform 1 0 25116 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 27324 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_283
timestamp 1604681595
transform 1 0 27140 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_287
timestamp 1604681595
transform 1 0 27508 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1604681595
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1604681595
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp 1604681595
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604681595
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 1472 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3220 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_40
timestamp 1604681595
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_36
timestamp 1604681595
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_32
timestamp 1604681595
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_36
timestamp 1604681595
transform 1 0 4416 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_48
timestamp 1604681595
transform 1 0 5520 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4968 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4968 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_55
timestamp 1604681595
transform 1 0 6164 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_57
timestamp 1604681595
transform 1 0 6348 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_53
timestamp 1604681595
transform 1 0 5980 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6164 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 6992 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6992 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_63
timestamp 1604681595
transform 1 0 6900 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_73
timestamp 1604681595
transform 1 0 7820 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_73
timestamp 1604681595
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_77
timestamp 1604681595
transform 1 0 8188 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_91
timestamp 1604681595
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_87
timestamp 1604681595
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1604681595
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1604681595
transform 1 0 8924 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_95
timestamp 1604681595
transform 1 0 9844 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_102
timestamp 1604681595
transform 1 0 10488 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_98
timestamp 1604681595
transform 1 0 10120 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10304 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9936 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9936 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10580 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_7_109
timestamp 1604681595
transform 1 0 11132 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_105
timestamp 1604681595
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_112
timestamp 1604681595
transform 1 0 11408 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_117
timestamp 1604681595
transform 1 0 11868 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12144 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13616 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_129
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_134
timestamp 1604681595
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_138
timestamp 1604681595
transform 1 0 13800 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_127
timestamp 1604681595
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_131
timestamp 1604681595
transform 1 0 13156 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_143
timestamp 1604681595
transform 1 0 14260 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_156
timestamp 1604681595
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_152
timestamp 1604681595
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_149
timestamp 1604681595
transform 1 0 14812 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_6_150
timestamp 1604681595
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15824 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15824 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1604681595
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_169
timestamp 1604681595
transform 1 0 16652 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604681595
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_186
timestamp 1604681595
transform 1 0 18216 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_183
timestamp 1604681595
transform 1 0 17940 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_179
timestamp 1604681595
transform 1 0 17572 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1604681595
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1604681595
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_196
timestamp 1604681595
transform 1 0 19136 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1604681595
transform 1 0 18768 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_7_201
timestamp 1604681595
transform 1 0 19596 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_206
timestamp 1604681595
transform 1 0 20056 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1604681595
transform 1 0 20516 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 20332 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 20516 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_210
timestamp 1604681595
transform 1 0 20424 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1604681595
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_218
timestamp 1604681595
transform 1 0 21160 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1604681595
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_238
timestamp 1604681595
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_234
timestamp 1604681595
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_230
timestamp 1604681595
transform 1 0 22264 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 22448 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_242
timestamp 1604681595
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_250
timestamp 1604681595
transform 1 0 24104 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 22356 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 24380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 25116 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_262
timestamp 1604681595
transform 1 0 25208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_266
timestamp 1604681595
transform 1 0 25576 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_255
timestamp 1604681595
transform 1 0 24564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_259
timestamp 1604681595
transform 1 0 24932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_263
timestamp 1604681595
transform 1 0 25300 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_279
timestamp 1604681595
transform 1 0 26772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_271
timestamp 1604681595
transform 1 0 26036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_274
timestamp 1604681595
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 26220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 26956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 26404 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_283
timestamp 1604681595
transform 1 0 27140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_280
timestamp 1604681595
transform 1 0 26864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 28888 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_292
timestamp 1604681595
transform 1 0 27968 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_298
timestamp 1604681595
transform 1 0 28520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_295
timestamp 1604681595
transform 1 0 28244 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604681595
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 2300 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_7
timestamp 1604681595
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1604681595
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_25
timestamp 1604681595
transform 1 0 3404 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_41
timestamp 1604681595
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5796 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_45
timestamp 1604681595
transform 1 0 5244 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_60
timestamp 1604681595
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_64
timestamp 1604681595
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_71
timestamp 1604681595
transform 1 0 7636 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1604681595
transform 1 0 8924 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1604681595
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_102
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12144 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_114
timestamp 1604681595
transform 1 0 11592 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 13708 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_133
timestamp 1604681595
transform 1 0 13340 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_140
timestamp 1604681595
transform 1 0 13984 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_144
timestamp 1604681595
transform 1 0 14352 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_147
timestamp 1604681595
transform 1 0 14628 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_162
timestamp 1604681595
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_165
timestamp 1604681595
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 17020 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16836 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_169
timestamp 1604681595
transform 1 0 16652 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_182
timestamp 1604681595
transform 1 0 17848 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_186
timestamp 1604681595
transform 1 0 18216 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18584 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_199
timestamp 1604681595
transform 1 0 19412 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_203
timestamp 1604681595
transform 1 0 19780 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_206
timestamp 1604681595
transform 1 0 20056 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 20516 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 21160 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 21528 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_210
timestamp 1604681595
transform 1 0 20424 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604681595
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_220
timestamp 1604681595
transform 1 0 21344 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_224
timestamp 1604681595
transform 1 0 21712 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1604681595
transform 1 0 22448 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 24012 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_241
timestamp 1604681595
transform 1 0 23276 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24380 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_251
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_262
timestamp 1604681595
transform 1 0 25208 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_270
timestamp 1604681595
transform 1 0 25944 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 26128 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_274
timestamp 1604681595
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_280
timestamp 1604681595
transform 1 0 26864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_292
timestamp 1604681595
transform 1 0 27968 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1604681595
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1472 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_23
timestamp 1604681595
transform 1 0 3220 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_31
timestamp 1604681595
transform 1 0 3956 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_34
timestamp 1604681595
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_38
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_48
timestamp 1604681595
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_42
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5704 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604681595
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_52
timestamp 1604681595
transform 1 0 5888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 8740 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_71
timestamp 1604681595
transform 1 0 7636 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_79
timestamp 1604681595
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_102
timestamp 1604681595
transform 1 0 10488 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1604681595
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12880 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 14444 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_137
timestamp 1604681595
transform 1 0 13708 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16100 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_154
timestamp 1604681595
transform 1 0 15272 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_159
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1604681595
transform 1 0 18124 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_172
timestamp 1604681595
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_176
timestamp 1604681595
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_180
timestamp 1604681595
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 19872 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 19688 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_188
timestamp 1604681595
transform 1 0 18400 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_200
timestamp 1604681595
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_223
timestamp 1604681595
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_227
timestamp 1604681595
transform 1 0 21988 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 23828 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_239
timestamp 1604681595
transform 1 0 23092 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_249
timestamp 1604681595
transform 1 0 24012 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24380 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24196 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 25944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 25392 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_262
timestamp 1604681595
transform 1 0 25208 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_266
timestamp 1604681595
transform 1 0 25576 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 26128 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_9_291
timestamp 1604681595
transform 1 0 27876 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 28888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_7
timestamp 1604681595
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_11
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_41
timestamp 1604681595
transform 1 0 4876 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5704 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp 1604681595
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_69
timestamp 1604681595
transform 1 0 7452 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_81
timestamp 1604681595
transform 1 0 8556 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_89
timestamp 1604681595
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_103
timestamp 1604681595
transform 1 0 10580 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11408 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_10_111
timestamp 1604681595
transform 1 0 11316 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_131
timestamp 1604681595
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_143
timestamp 1604681595
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15916 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_147
timestamp 1604681595
transform 1 0 14628 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_160
timestamp 1604681595
transform 1 0 15824 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_170
timestamp 1604681595
transform 1 0 16744 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_182
timestamp 1604681595
transform 1 0 17848 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_194
timestamp 1604681595
transform 1 0 18952 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_208
timestamp 1604681595
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1604681595
transform 1 0 21160 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1604681595
transform 1 0 24012 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23184 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_239
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_242
timestamp 1604681595
transform 1 0 23368 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_247
timestamp 1604681595
transform 1 0 23828 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_258
timestamp 1604681595
transform 1 0 24840 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_262
timestamp 1604681595
transform 1 0 25208 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_270
timestamp 1604681595
transform 1 0 25944 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_274
timestamp 1604681595
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_280
timestamp 1604681595
transform 1 0 26864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_292
timestamp 1604681595
transform 1 0 27968 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp 1604681595
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604681595
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1604681595
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4416 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_32
timestamp 1604681595
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_45
timestamp 1604681595
transform 1 0 5244 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_66
timestamp 1604681595
transform 1 0 7176 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_74
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_78
timestamp 1604681595
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_82
timestamp 1604681595
transform 1 0 8648 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9752 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_90
timestamp 1604681595
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1604681595
transform 1 0 11500 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1604681595
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14444 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_143
timestamp 1604681595
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_11_166
timestamp 1604681595
transform 1 0 16376 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1604681595
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_176
timestamp 1604681595
transform 1 0 17296 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1604681595
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20056 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 18768 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_195
timestamp 1604681595
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_199
timestamp 1604681595
transform 1 0 19412 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_203
timestamp 1604681595
transform 1 0 19780 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 21988 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1604681595
transform 1 0 21804 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_229
timestamp 1604681595
transform 1 0 22172 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_235
timestamp 1604681595
transform 1 0 22724 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_238
timestamp 1604681595
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_242
timestamp 1604681595
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_254
timestamp 1604681595
transform 1 0 24472 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_258
timestamp 1604681595
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_262
timestamp 1604681595
transform 1 0 25208 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 26496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_274
timestamp 1604681595
transform 1 0 26312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_278
timestamp 1604681595
transform 1 0 26680 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_290
timestamp 1604681595
transform 1 0 27784 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_298
timestamp 1604681595
transform 1 0 28520 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 1932 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2300 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1604681595
transform 1 0 2116 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_38
timestamp 1604681595
transform 1 0 4600 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_50
timestamp 1604681595
transform 1 0 5704 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_62
timestamp 1604681595
transform 1 0 6808 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7728 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 6900 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_66
timestamp 1604681595
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_70
timestamp 1604681595
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_81
timestamp 1604681595
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 10396 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 9292 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1604681595
transform 1 0 8924 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1604681595
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_104
timestamp 1604681595
transform 1 0 10672 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_116
timestamp 1604681595
transform 1 0 11776 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 13156 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13524 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_128
timestamp 1604681595
transform 1 0 12880 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1604681595
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_137
timestamp 1604681595
transform 1 0 13708 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_145
timestamp 1604681595
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1604681595
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_166
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16744 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 18768 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19136 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19504 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_189
timestamp 1604681595
transform 1 0 18492 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1604681595
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_198
timestamp 1604681595
transform 1 0 19320 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1604681595
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 22080 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_226
timestamp 1604681595
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23184 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 22448 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_230
timestamp 1604681595
transform 1 0 22264 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_234
timestamp 1604681595
transform 1 0 22632 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_249
timestamp 1604681595
transform 1 0 24012 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25576 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1604681595
transform 1 0 24380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_265
timestamp 1604681595
transform 1 0 25484 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_268
timestamp 1604681595
transform 1 0 25760 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_274
timestamp 1604681595
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_280
timestamp 1604681595
transform 1 0 26864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_292
timestamp 1604681595
transform 1 0 27968 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_298
timestamp 1604681595
transform 1 0 28520 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604681595
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1564 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_18
timestamp 1604681595
transform 1 0 2760 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_14
timestamp 1604681595
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_19
timestamp 1604681595
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_11
timestamp 1604681595
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 2576 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604681595
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_23
timestamp 1604681595
transform 1 0 3220 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1604681595
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4140 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_52
timestamp 1604681595
transform 1 0 5888 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_58
timestamp 1604681595
transform 1 0 6440 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_61
timestamp 1604681595
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_65
timestamp 1604681595
transform 1 0 7084 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_68
timestamp 1604681595
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7176 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7728 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1604681595
transform 1 0 8372 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_75
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1604681595
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 8740 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1604681595
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_86
timestamp 1604681595
transform 1 0 9016 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_85
timestamp 1604681595
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9292 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9292 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_99
timestamp 1604681595
transform 1 0 10212 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_104
timestamp 1604681595
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_98
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10488 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_108
timestamp 1604681595
transform 1 0 11040 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_121
timestamp 1604681595
transform 1 0 12236 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 13156 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13432 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_127
timestamp 1604681595
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_129
timestamp 1604681595
transform 1 0 12972 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_133
timestamp 1604681595
transform 1 0 13340 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_143
timestamp 1604681595
transform 1 0 14260 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1604681595
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1604681595
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_150
timestamp 1604681595
transform 1 0 14904 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_163
timestamp 1604681595
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_160
timestamp 1604681595
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_164
timestamp 1604681595
transform 1 0 16192 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_172
timestamp 1604681595
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_167
timestamp 1604681595
transform 1 0 16468 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_184
timestamp 1604681595
transform 1 0 18032 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_176
timestamp 1604681595
transform 1 0 17296 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1604681595
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_176
timestamp 1604681595
transform 1 0 17296 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18308 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18768 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18768 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18584 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_188
timestamp 1604681595
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_201
timestamp 1604681595
transform 1 0 19596 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_205
timestamp 1604681595
transform 1 0 19964 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_189
timestamp 1604681595
transform 1 0 18492 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_201
timestamp 1604681595
transform 1 0 19596 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1604681595
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_218
timestamp 1604681595
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_215
timestamp 1604681595
transform 1 0 20884 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_211
timestamp 1604681595
transform 1 0 20516 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 20332 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 20332 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1604681595
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_222
timestamp 1604681595
transform 1 0 21528 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1604681595
transform 1 0 21988 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 21344 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1604681595
transform 1 0 23828 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 23644 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_236
timestamp 1604681595
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_240
timestamp 1604681595
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 25576 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 25392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_254
timestamp 1604681595
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_258
timestamp 1604681595
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_262
timestamp 1604681595
transform 1 0 25208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_256
timestamp 1604681595
transform 1 0 24656 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_268
timestamp 1604681595
transform 1 0 25760 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 27508 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_285
timestamp 1604681595
transform 1 0 27324 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_289
timestamp 1604681595
transform 1 0 27692 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_274
timestamp 1604681595
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_280
timestamp 1604681595
transform 1 0 26864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_297
timestamp 1604681595
transform 1 0 28428 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_292
timestamp 1604681595
transform 1 0 27968 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_298
timestamp 1604681595
transform 1 0 28520 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_7
timestamp 1604681595
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_11
timestamp 1604681595
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1604681595
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 3036 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_15_40
timestamp 1604681595
transform 1 0 4784 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_48
timestamp 1604681595
transform 1 0 5520 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7084 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_82
timestamp 1604681595
transform 1 0 8648 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10028 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_85
timestamp 1604681595
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1604681595
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1604681595
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 12604 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_106
timestamp 1604681595
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 14260 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 12972 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_127
timestamp 1604681595
transform 1 0 12788 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_131
timestamp 1604681595
transform 1 0 13156 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_139
timestamp 1604681595
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15824 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_152
timestamp 1604681595
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_156
timestamp 1604681595
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 18308 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1604681595
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_173
timestamp 1604681595
transform 1 0 17020 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18860 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_189
timestamp 1604681595
transform 1 0 18492 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_202
timestamp 1604681595
transform 1 0 19688 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 21988 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_214
timestamp 1604681595
transform 1 0 20792 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_222
timestamp 1604681595
transform 1 0 21528 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1604681595
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_229
timestamp 1604681595
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_233
timestamp 1604681595
transform 1 0 22540 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_241
timestamp 1604681595
transform 1 0 23276 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_248
timestamp 1604681595
transform 1 0 23920 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 25300 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_260
timestamp 1604681595
transform 1 0 25024 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_265
timestamp 1604681595
transform 1 0 25484 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 26404 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 27508 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 26956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 27324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_273
timestamp 1604681595
transform 1 0 26220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_279
timestamp 1604681595
transform 1 0 26772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_283
timestamp 1604681595
transform 1 0 27140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_291
timestamp 1604681595
transform 1 0 27876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 28060 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_295
timestamp 1604681595
transform 1 0 28244 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 1932 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604681595
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1604681595
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_18
timestamp 1604681595
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_22
timestamp 1604681595
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_26
timestamp 1604681595
transform 1 0 3496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1604681595
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6532 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_56
timestamp 1604681595
transform 1 0 6256 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_68
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_72
timestamp 1604681595
transform 1 0 7728 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_82
timestamp 1604681595
transform 1 0 8648 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_102
timestamp 1604681595
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12420 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_16_106
timestamp 1604681595
transform 1 0 10856 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_118
timestamp 1604681595
transform 1 0 11960 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_122
timestamp 1604681595
transform 1 0 12328 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_142
timestamp 1604681595
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 15732 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_146
timestamp 1604681595
transform 1 0 14536 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1604681595
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_157
timestamp 1604681595
transform 1 0 15548 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_161
timestamp 1604681595
transform 1 0 15916 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_165
timestamp 1604681595
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18308 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16744 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 17756 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_169
timestamp 1604681595
transform 1 0 16652 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_179
timestamp 1604681595
transform 1 0 17572 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_183
timestamp 1604681595
transform 1 0 17940 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19320 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_196
timestamp 1604681595
transform 1 0 19136 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_200
timestamp 1604681595
transform 1 0 19504 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1604681595
transform 1 0 21620 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 21436 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1604681595
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_219
timestamp 1604681595
transform 1 0 21252 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_232
timestamp 1604681595
transform 1 0 22448 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_244
timestamp 1604681595
transform 1 0 23552 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_250
timestamp 1604681595
transform 1 0 24104 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 25300 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 24840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_253
timestamp 1604681595
transform 1 0 24380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_257
timestamp 1604681595
transform 1 0 24748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_260
timestamp 1604681595
transform 1 0 25024 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_267
timestamp 1604681595
transform 1 0 25668 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 27600 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 27048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 27416 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_280
timestamp 1604681595
transform 1 0 26864 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_284
timestamp 1604681595
transform 1 0 27232 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_291
timestamp 1604681595
transform 1 0 27876 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 28888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_16
timestamp 1604681595
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_20
timestamp 1604681595
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1604681595
transform 1 0 4416 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604681595
transform 1 0 3312 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604681595
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_28
timestamp 1604681595
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_32
timestamp 1604681595
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_39
timestamp 1604681595
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_43
timestamp 1604681595
transform 1 0 5060 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604681595
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8464 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_71
timestamp 1604681595
transform 1 0 7636 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_77
timestamp 1604681595
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_99
timestamp 1604681595
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_103
timestamp 1604681595
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 10948 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13800 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_135
timestamp 1604681595
transform 1 0 13524 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15640 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_167
timestamp 1604681595
transform 1 0 16468 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 16652 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_171
timestamp 1604681595
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604681595
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604681595
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18400 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_197
timestamp 1604681595
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_201
timestamp 1604681595
transform 1 0 19596 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1604681595
transform 1 0 21436 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_209
timestamp 1604681595
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_213
timestamp 1604681595
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1604681595
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 24012 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_230
timestamp 1604681595
transform 1 0 22264 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_242
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 24196 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_17_270
timestamp 1604681595
transform 1 0 25944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1604681595
transform 1 0 26680 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 26496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 26128 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 27692 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_274
timestamp 1604681595
transform 1 0 26312 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_287
timestamp 1604681595
transform 1 0 27508 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_291
timestamp 1604681595
transform 1 0 27876 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 28888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1932 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_18
timestamp 1604681595
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4232 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_22
timestamp 1604681595
transform 1 0 3128 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_26
timestamp 1604681595
transform 1 0 3496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_53
timestamp 1604681595
transform 1 0 5980 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_61
timestamp 1604681595
transform 1 0 6716 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_64
timestamp 1604681595
transform 1 0 6992 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_76
timestamp 1604681595
transform 1 0 8096 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10212 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1604681595
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_108
timestamp 1604681595
transform 1 0 11040 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_120
timestamp 1604681595
transform 1 0 12144 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14260 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_132
timestamp 1604681595
transform 1 0 13248 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_138
timestamp 1604681595
transform 1 0 13800 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_142
timestamp 1604681595
transform 1 0 14168 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_145
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 17756 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_18_167
timestamp 1604681595
transform 1 0 16468 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_179
timestamp 1604681595
transform 1 0 17572 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_200
timestamp 1604681595
transform 1 0 19504 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_208
timestamp 1604681595
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1604681595
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_224
timestamp 1604681595
transform 1 0 21712 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 22448 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_235
timestamp 1604681595
transform 1 0 22724 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_247
timestamp 1604681595
transform 1 0 23828 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1604681595
transform 1 0 24840 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 24656 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 25852 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 24196 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_253
timestamp 1604681595
transform 1 0 24380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_267
timestamp 1604681595
transform 1 0 25668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 27508 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_271
timestamp 1604681595
transform 1 0 26036 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_285
timestamp 1604681595
transform 1 0 27324 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_289
timestamp 1604681595
transform 1 0 27692 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 28888 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp 1604681595
transform 1 0 28428 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_9
timestamp 1604681595
transform 1 0 1932 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1748 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_16
timestamp 1604681595
transform 1 0 2576 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_19
timestamp 1604681595
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2024 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_20
timestamp 1604681595
transform 1 0 2944 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_24
timestamp 1604681595
transform 1 0 3312 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_23
timestamp 1604681595
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3128 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_40
timestamp 1604681595
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1604681595
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4232 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_19_48
timestamp 1604681595
transform 1 0 5520 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_44
timestamp 1604681595
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_61
timestamp 1604681595
transform 1 0 6716 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_55
timestamp 1604681595
transform 1 0 6164 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_56
timestamp 1604681595
transform 1 0 6256 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_43
timestamp 1604681595
transform 1 0 5060 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 8188 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_81
timestamp 1604681595
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_64
timestamp 1604681595
transform 1 0 6992 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_72
timestamp 1604681595
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_76
timestamp 1604681595
transform 1 0 8096 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_80
timestamp 1604681595
transform 1 0 8464 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_89
timestamp 1604681595
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_86
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_85
timestamp 1604681595
transform 1 0 8924 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_102
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_103
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_99
timestamp 1604681595
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_95
timestamp 1604681595
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_112
timestamp 1604681595
transform 1 0 11408 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_108
timestamp 1604681595
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1604681595
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11224 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1604681595
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_117
timestamp 1604681595
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12052 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1604681595
transform 1 0 11684 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_20_124
timestamp 1604681595
transform 1 0 12512 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 14260 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_131
timestamp 1604681595
transform 1 0 13156 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_134
timestamp 1604681595
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_138
timestamp 1604681595
transform 1 0 13800 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_156
timestamp 1604681595
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_152
timestamp 1604681595
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1604681595
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_163
timestamp 1604681595
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_164
timestamp 1604681595
transform 1 0 16192 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18308 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_176
timestamp 1604681595
transform 1 0 17296 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_175
timestamp 1604681595
transform 1 0 17204 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_193
timestamp 1604681595
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_189
timestamp 1604681595
transform 1 0 18492 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_197
timestamp 1604681595
transform 1 0 19228 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_193
timestamp 1604681595
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18676 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_205
timestamp 1604681595
transform 1 0 19964 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1604681595
transform 1 0 19228 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 20424 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_229
timestamp 1604681595
transform 1 0 22172 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_209
timestamp 1604681595
transform 1 0 20332 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1604681595
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_229
timestamp 1604681595
transform 1 0 22172 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23644 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24012 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22448 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_241
timestamp 1604681595
transform 1 0 23276 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_234
timestamp 1604681595
transform 1 0 22632 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_242
timestamp 1604681595
transform 1 0 23368 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_247
timestamp 1604681595
transform 1 0 23828 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_257
timestamp 1604681595
transform 1 0 24748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_251
timestamp 1604681595
transform 1 0 24196 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_257
timestamp 1604681595
transform 1 0 24748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_253
timestamp 1604681595
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24196 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 24564 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1604681595
transform 1 0 24840 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_267
timestamp 1604681595
transform 1 0 25668 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_261
timestamp 1604681595
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 25300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1604681595
transform 1 0 25484 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_274
timestamp 1604681595
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_271
timestamp 1604681595
transform 1 0 26036 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_274
timestamp 1604681595
transform 1 0 26312 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 26496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_288
timestamp 1604681595
transform 1 0 27600 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_290
timestamp 1604681595
transform 1 0 27784 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_278
timestamp 1604681595
transform 1 0 26680 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_298
timestamp 1604681595
transform 1 0 28520 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_296
timestamp 1604681595
transform 1 0 28336 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 1748 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_16
timestamp 1604681595
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_20
timestamp 1604681595
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4232 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_24
timestamp 1604681595
transform 1 0 3312 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_30
timestamp 1604681595
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 5244 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_43
timestamp 1604681595
transform 1 0 5060 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_47
timestamp 1604681595
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7544 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7360 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_66
timestamp 1604681595
transform 1 0 7176 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_79
timestamp 1604681595
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1604681595
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9108 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_96
timestamp 1604681595
transform 1 0 9936 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1604681595
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14260 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13708 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_136
timestamp 1604681595
transform 1 0 13616 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_139
timestamp 1604681595
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_152
timestamp 1604681595
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_156
timestamp 1604681595
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_160
timestamp 1604681595
transform 1 0 15824 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18216 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_172
timestamp 1604681595
transform 1 0 16928 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_176
timestamp 1604681595
transform 1 0 17296 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1604681595
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 20148 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_205
timestamp 1604681595
transform 1 0 19964 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_209
timestamp 1604681595
transform 1 0 20332 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_221
timestamp 1604681595
transform 1 0 21436 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_236
timestamp 1604681595
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 25944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_254
timestamp 1604681595
transform 1 0 24472 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_266
timestamp 1604681595
transform 1 0 25576 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 26128 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_21_291
timestamp 1604681595
transform 1 0 27876 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 28888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1472 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_36
timestamp 1604681595
transform 1 0 4416 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7636 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_63
timestamp 1604681595
transform 1 0 6900 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_80
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9108 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_86
timestamp 1604681595
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_89
timestamp 1604681595
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_101
timestamp 1604681595
transform 1 0 10396 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1604681595
transform 1 0 11224 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_106
timestamp 1604681595
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_119
timestamp 1604681595
transform 1 0 12052 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_125
timestamp 1604681595
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1604681595
transform 1 0 12788 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14260 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_130
timestamp 1604681595
transform 1 0 13064 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_142
timestamp 1604681595
transform 1 0 14168 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18308 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_173
timestamp 1604681595
transform 1 0 17020 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_181
timestamp 1604681595
transform 1 0 17756 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_186
timestamp 1604681595
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 19872 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19320 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_196
timestamp 1604681595
transform 1 0 19136 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_200
timestamp 1604681595
transform 1 0 19504 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_207
timestamp 1604681595
transform 1 0 20148 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_213
timestamp 1604681595
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_229
timestamp 1604681595
transform 1 0 22172 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 22448 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 24564 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_251
timestamp 1604681595
transform 1 0 24196 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_257
timestamp 1604681595
transform 1 0 24748 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_269
timestamp 1604681595
transform 1 0 25852 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_288
timestamp 1604681595
transform 1 0 27600 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 28888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_296
timestamp 1604681595
transform 1 0 28336 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_7
timestamp 1604681595
transform 1 0 1748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_19
timestamp 1604681595
transform 1 0 2852 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_31
timestamp 1604681595
transform 1 0 3956 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_34
timestamp 1604681595
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_38
timestamp 1604681595
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_42
timestamp 1604681595
transform 1 0 4968 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_54
timestamp 1604681595
transform 1 0 6072 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7636 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7452 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 6992 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_66
timestamp 1604681595
transform 1 0 7176 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_90
timestamp 1604681595
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_94
timestamp 1604681595
transform 1 0 9752 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_106
timestamp 1604681595
transform 1 0 10856 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_110
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1604681595
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_117
timestamp 1604681595
transform 1 0 11868 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1604681595
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_147
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_153
timestamp 1604681595
transform 1 0 15180 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_156
timestamp 1604681595
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_160
timestamp 1604681595
transform 1 0 15824 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18216 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_172
timestamp 1604681595
transform 1 0 16928 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_176
timestamp 1604681595
transform 1 0 17296 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604681595
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18952 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18768 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_188
timestamp 1604681595
transform 1 0 18400 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 21436 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_213
timestamp 1604681595
transform 1 0 20700 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_224
timestamp 1604681595
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_228
timestamp 1604681595
transform 1 0 22080 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 24012 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 22264 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1604681595
transform 1 0 24564 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 24380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_251
timestamp 1604681595
transform 1 0 24196 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_264
timestamp 1604681595
transform 1 0 25392 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 26496 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_278
timestamp 1604681595
transform 1 0 26680 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_290
timestamp 1604681595
transform 1 0 27784 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_298
timestamp 1604681595
transform 1 0 28520 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1604681595
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_16
timestamp 1604681595
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_11
timestamp 1604681595
transform 1 0 2116 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2392 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1604681595
transform 1 0 2944 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_28
timestamp 1604681595
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1604681595
transform 1 0 4876 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1604681595
transform 1 0 5980 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_65
timestamp 1604681595
transform 1 0 7084 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_73
timestamp 1604681595
transform 1 0 7820 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1604681595
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 9200 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10304 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_86
timestamp 1604681595
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1604681595
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_99
timestamp 1604681595
transform 1 0 10212 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_102
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 11316 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_24_110
timestamp 1604681595
transform 1 0 11224 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_130
timestamp 1604681595
transform 1 0 13064 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_142
timestamp 1604681595
transform 1 0 14168 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1604681595
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 17756 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_173
timestamp 1604681595
transform 1 0 17020 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 19136 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1604681595
transform 1 0 18860 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_198
timestamp 1604681595
transform 1 0 19320 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 21712 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_210
timestamp 1604681595
transform 1 0 20424 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_223
timestamp 1604681595
transform 1 0 21620 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 24012 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_243
timestamp 1604681595
transform 1 0 23460 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 24380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 24748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_251
timestamp 1604681595
transform 1 0 24196 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_255
timestamp 1604681595
transform 1 0 24564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_259
timestamp 1604681595
transform 1 0 24932 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_267
timestamp 1604681595
transform 1 0 25668 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_271
timestamp 1604681595
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_280
timestamp 1604681595
transform 1 0 26864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_292
timestamp 1604681595
transform 1 0 27968 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_298
timestamp 1604681595
transform 1 0 28520 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3864 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3312 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_22
timestamp 1604681595
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_26
timestamp 1604681595
transform 1 0 3496 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 5244 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_43
timestamp 1604681595
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_47
timestamp 1604681595
transform 1 0 5428 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_55
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7360 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_66
timestamp 1604681595
transform 1 0 7176 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_70
timestamp 1604681595
transform 1 0 7544 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8832 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_25_103
timestamp 1604681595
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_107
timestamp 1604681595
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_111
timestamp 1604681595
transform 1 0 11316 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_119
timestamp 1604681595
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_127
timestamp 1604681595
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_131
timestamp 1604681595
transform 1 0 13156 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_143
timestamp 1604681595
transform 1 0 14260 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_151
timestamp 1604681595
transform 1 0 14996 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_156
timestamp 1604681595
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_160
timestamp 1604681595
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_164
timestamp 1604681595
transform 1 0 16192 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 18216 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_176
timestamp 1604681595
transform 1 0 17296 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_180
timestamp 1604681595
transform 1 0 17664 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1604681595
transform 1 0 19136 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 18952 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 18584 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_188
timestamp 1604681595
transform 1 0 18400 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_192
timestamp 1604681595
transform 1 0 18768 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_205
timestamp 1604681595
transform 1 0 19964 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_213
timestamp 1604681595
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_217
timestamp 1604681595
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_221
timestamp 1604681595
transform 1 0 21436 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1604681595
transform 1 0 23920 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_233
timestamp 1604681595
transform 1 0 22540 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_237
timestamp 1604681595
transform 1 0 22908 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604681595
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 25668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 24932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_257
timestamp 1604681595
transform 1 0 24748 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_261
timestamp 1604681595
transform 1 0 25116 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_288
timestamp 1604681595
transform 1 0 27600 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_296
timestamp 1604681595
transform 1 0 28336 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1604681595
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_7
timestamp 1604681595
transform 1 0 1748 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604681595
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_11
timestamp 1604681595
transform 1 0 2116 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_13
timestamp 1604681595
transform 1 0 2300 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2760 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4232 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_36
timestamp 1604681595
transform 1 0 4416 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_39
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_47
timestamp 1604681595
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_44
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 5244 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_54
timestamp 1604681595
transform 1 0 6072 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_81
timestamp 1604681595
transform 1 0 8556 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_77
timestamp 1604681595
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_81
timestamp 1604681595
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_92
timestamp 1604681595
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_89
timestamp 1604681595
transform 1 0 9292 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_85
timestamp 1604681595
transform 1 0 8924 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_89
timestamp 1604681595
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_98
timestamp 1604681595
transform 1 0 10120 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 9936 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9936 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10304 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1604681595
transform 1 0 11500 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_109
timestamp 1604681595
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_105
timestamp 1604681595
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10948 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1604681595
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_121
timestamp 1604681595
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1604681595
transform 1 0 11132 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_133
timestamp 1604681595
transform 1 0 13340 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_129
timestamp 1604681595
transform 1 0 12972 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12788 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13156 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1604681595
transform 1 0 14076 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_137
timestamp 1604681595
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_142
timestamp 1604681595
transform 1 0 14168 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 14260 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 14444 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_154
timestamp 1604681595
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_147
timestamp 1604681595
transform 1 0 14628 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_158
timestamp 1604681595
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_163
timestamp 1604681595
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16008 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1604681595
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_171
timestamp 1604681595
transform 1 0 16836 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1604681595
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_185
timestamp 1604681595
transform 1 0 18124 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_179
timestamp 1604681595
transform 1 0 17572 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18216 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18124 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_26_167
timestamp 1604681595
transform 1 0 16468 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_194
timestamp 1604681595
transform 1 0 18952 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_195
timestamp 1604681595
transform 1 0 19044 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 19228 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_203
timestamp 1604681595
transform 1 0 19780 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_199
timestamp 1604681595
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 19964 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_207
timestamp 1604681595
transform 1 0 20148 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_199
timestamp 1604681595
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_211
timestamp 1604681595
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_219
timestamp 1604681595
transform 1 0 21252 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_236
timestamp 1604681595
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_231
timestamp 1604681595
transform 1 0 22356 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_234
timestamp 1604681595
transform 1 0 22632 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22632 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_240
timestamp 1604681595
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_248
timestamp 1604681595
transform 1 0 23920 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_244
timestamp 1604681595
transform 1 0 23552 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23828 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24012 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24012 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_26_258
timestamp 1604681595
transform 1 0 24840 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_270
timestamp 1604681595
transform 1 0 25944 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_258
timestamp 1604681595
transform 1 0 24840 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_270
timestamp 1604681595
transform 1 0 25944 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 26404 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 26956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_274
timestamp 1604681595
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_288
timestamp 1604681595
transform 1 0 27600 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_274
timestamp 1604681595
transform 1 0 26312 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_279
timestamp 1604681595
transform 1 0 26772 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_283
timestamp 1604681595
transform 1 0 27140 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 28888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_296
timestamp 1604681595
transform 1 0 28336 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_295
timestamp 1604681595
transform 1 0 28244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2760 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_7
timestamp 1604681595
transform 1 0 1748 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_20
timestamp 1604681595
transform 1 0 2944 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3128 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_24
timestamp 1604681595
transform 1 0 3312 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1604681595
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 5244 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_28_44
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 7176 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7544 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_64
timestamp 1604681595
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_72
timestamp 1604681595
transform 1 0 7728 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10304 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9936 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_98
timestamp 1604681595
transform 1 0 10120 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1604681595
transform 1 0 11132 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1604681595
transform 1 0 12236 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_133
timestamp 1604681595
transform 1 0 13340 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_145
timestamp 1604681595
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16192 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16008 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18124 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_183
timestamp 1604681595
transform 1 0 17940 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_187
timestamp 1604681595
transform 1 0 18308 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_195
timestamp 1604681595
transform 1 0 19044 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_206
timestamp 1604681595
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 21344 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1604681595
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_222
timestamp 1604681595
transform 1 0 21528 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23368 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22632 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_236
timestamp 1604681595
transform 1 0 22816 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_240
timestamp 1604681595
transform 1 0 23184 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 24748 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_251
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_255
timestamp 1604681595
transform 1 0 24564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_259
timestamp 1604681595
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_271
timestamp 1604681595
transform 1 0 26036 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_274
timestamp 1604681595
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_288
timestamp 1604681595
transform 1 0 27600 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 28888 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_296
timestamp 1604681595
transform 1 0 28336 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_7
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_11
timestamp 1604681595
transform 1 0 2116 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_17
timestamp 1604681595
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 3036 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_30
timestamp 1604681595
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_34
timestamp 1604681595
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_38
timestamp 1604681595
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_42
timestamp 1604681595
transform 1 0 4968 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_54
timestamp 1604681595
transform 1 0 6072 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_71
timestamp 1604681595
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_75
timestamp 1604681595
transform 1 0 8004 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9752 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9568 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_87
timestamp 1604681595
transform 1 0 9108 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_90
timestamp 1604681595
transform 1 0 9384 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_103
timestamp 1604681595
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_107
timestamp 1604681595
transform 1 0 10948 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_111
timestamp 1604681595
transform 1 0 11316 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_119
timestamp 1604681595
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 14076 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13156 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12788 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_129
timestamp 1604681595
transform 1 0 12972 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_133
timestamp 1604681595
transform 1 0 13340 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_137
timestamp 1604681595
transform 1 0 13708 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 15088 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_150
timestamp 1604681595
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_154
timestamp 1604681595
transform 1 0 15272 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1604681595
transform 1 0 16376 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_170
timestamp 1604681595
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_174
timestamp 1604681595
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_178
timestamp 1604681595
transform 1 0 17480 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 17296 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1604681595
transform 1 0 19780 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_189
timestamp 1604681595
transform 1 0 18492 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_195
timestamp 1604681595
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_199
timestamp 1604681595
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 21160 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_212
timestamp 1604681595
transform 1 0 20608 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_229
timestamp 1604681595
transform 1 0 22172 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 22632 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_233
timestamp 1604681595
transform 1 0 22540 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_236
timestamp 1604681595
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_240
timestamp 1604681595
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 25944 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_254
timestamp 1604681595
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_258
timestamp 1604681595
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_262
timestamp 1604681595
transform 1 0 25208 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 26128 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_29_291
timestamp 1604681595
transform 1 0 27876 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1472 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_23
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1604681595
transform 1 0 4876 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1604681595
transform 1 0 6164 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_53
timestamp 1604681595
transform 1 0 5980 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_58
timestamp 1604681595
transform 1 0 6440 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7176 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_64
timestamp 1604681595
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_75
timestamp 1604681595
transform 1 0 8004 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1604681595
transform 1 0 8372 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1604681595
transform 1 0 8740 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10580 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_86
timestamp 1604681595
transform 1 0 9016 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_97
timestamp 1604681595
transform 1 0 10028 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_122
timestamp 1604681595
transform 1 0 12328 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_134
timestamp 1604681595
transform 1 0 13432 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_145
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 15732 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_158
timestamp 1604681595
transform 1 0 15640 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_161
timestamp 1604681595
transform 1 0 15916 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_165
timestamp 1604681595
transform 1 0 16284 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18308 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1604681595
transform 1 0 16560 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_177
timestamp 1604681595
transform 1 0 17388 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_185
timestamp 1604681595
transform 1 0 18124 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_206
timestamp 1604681595
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 21344 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_218
timestamp 1604681595
transform 1 0 21160 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_222
timestamp 1604681595
transform 1 0 21528 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_226
timestamp 1604681595
transform 1 0 21896 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_229
timestamp 1604681595
transform 1 0 22172 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1604681595
transform 1 0 22632 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23644 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 22356 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_233
timestamp 1604681595
transform 1 0 22540 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_243
timestamp 1604681595
transform 1 0 23460 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_247
timestamp 1604681595
transform 1 0 23828 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1604681595
transform 1 0 24380 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_30_262
timestamp 1604681595
transform 1 0 25208 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_274
timestamp 1604681595
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_288
timestamp 1604681595
transform 1 0 27600 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 28888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_296
timestamp 1604681595
transform 1 0 28336 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_17
timestamp 1604681595
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 4600 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 3036 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_31_30
timestamp 1604681595
transform 1 0 3864 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1604681595
transform 1 0 4876 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 5244 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_47
timestamp 1604681595
transform 1 0 5428 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604681595
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7084 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 8096 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_78
timestamp 1604681595
transform 1 0 8280 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8832 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1604681595
transform 1 0 9660 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10764 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_107
timestamp 1604681595
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_111
timestamp 1604681595
transform 1 0 11316 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1604681595
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 14352 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 13340 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 14168 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13708 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 12972 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_131
timestamp 1604681595
transform 1 0 13156 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_135
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_139
timestamp 1604681595
transform 1 0 13892 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 16284 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_163
timestamp 1604681595
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_174
timestamp 1604681595
transform 1 0 17112 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_171
timestamp 1604681595
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_167
timestamp 1604681595
transform 1 0 16468 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 17296 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1604681595
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_178
timestamp 1604681595
transform 1 0 17480 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 17664 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 21804 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 21436 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 21068 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_216
timestamp 1604681595
transform 1 0 20976 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_219
timestamp 1604681595
transform 1 0 21252 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_223
timestamp 1604681595
transform 1 0 21620 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_236
timestamp 1604681595
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_240
timestamp 1604681595
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1604681595
transform 1 0 25208 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 24656 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_254
timestamp 1604681595
transform 1 0 24472 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_258
timestamp 1604681595
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604681595
transform 1 0 26772 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1604681595
transform 1 0 26496 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_271
timestamp 1604681595
transform 1 0 26036 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_275
timestamp 1604681595
transform 1 0 26404 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_278
timestamp 1604681595
transform 1 0 26680 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_282
timestamp 1604681595
transform 1 0 27048 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 28888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_294
timestamp 1604681595
transform 1 0 28152 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_298
timestamp 1604681595
transform 1 0 28520 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 3036 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3496 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_23
timestamp 1604681595
transform 1 0 3220 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_28
timestamp 1604681595
transform 1 0 3680 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 5244 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7728 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 7544 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_64
timestamp 1604681595
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1604681595
transform 1 0 8556 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_86
timestamp 1604681595
transform 1 0 9016 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_32_124
timestamp 1604681595
transform 1 0 12512 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13340 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_132
timestamp 1604681595
transform 1 0 13248 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_142
timestamp 1604681595
transform 1 0 14168 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1604681595
transform 1 0 15732 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_146
timestamp 1604681595
transform 1 0 14536 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_152
timestamp 1604681595
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_158
timestamp 1604681595
transform 1 0 15640 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1604681595
transform 1 0 17296 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_168
timestamp 1604681595
transform 1 0 16560 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_185
timestamp 1604681595
transform 1 0 18124 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__0.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19228 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_199
timestamp 1604681595
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 21528 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_211
timestamp 1604681595
transform 1 0 20516 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_221
timestamp 1604681595
transform 1 0 21436 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 23644 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_241
timestamp 1604681595
transform 1 0 23276 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_247
timestamp 1604681595
transform 1 0 23828 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 25208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_259
timestamp 1604681595
transform 1 0 24932 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_264
timestamp 1604681595
transform 1 0 25392 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_272
timestamp 1604681595
transform 1 0 26128 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_280
timestamp 1604681595
transform 1 0 26864 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 28888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_292
timestamp 1604681595
transform 1 0 27968 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_298
timestamp 1604681595
transform 1 0 28520 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3496 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3312 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_23
timestamp 1604681595
transform 1 0 3220 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_45
timestamp 1604681595
transform 1 0 5244 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1604681595
transform 1 0 6348 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604681595
transform 1 0 6900 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8280 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 8096 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8280 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_67
timestamp 1604681595
transform 1 0 7268 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_75
timestamp 1604681595
transform 1 0 8004 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_76
timestamp 1604681595
transform 1 0 8096 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_97
timestamp 1604681595
transform 1 0 10028 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_109
timestamp 1604681595
transform 1 0 11132 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1604681595
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 13524 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 13340 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 13524 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_131
timestamp 1604681595
transform 1 0 13156 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_129
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_137
timestamp 1604681595
transform 1 0 13708 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_154
timestamp 1604681595
transform 1 0 15272 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_166
timestamp 1604681595
transform 1 0 16376 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_149
timestamp 1604681595
transform 1 0 14812 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_166
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1604681595
transform 1 0 17020 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_175
timestamp 1604681595
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_179
timestamp 1604681595
transform 1 0 17572 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_172
timestamp 1604681595
transform 1 0 16928 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_176
timestamp 1604681595
transform 1 0 17296 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_mode_io__0.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 19228 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__0.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_192
timestamp 1604681595
transform 1 0 18768 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_188
timestamp 1604681595
transform 1 0 18400 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_200
timestamp 1604681595
transform 1 0 19504 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 21712 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1604681595
transform 1 0 20976 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_228
timestamp 1604681595
transform 1 0 22080 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1604681595
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1604681595
transform 1 0 22264 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_240
timestamp 1604681595
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_247
timestamp 1604681595
transform 1 0 23828 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_264
timestamp 1604681595
transform 1 0 25392 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_259
timestamp 1604681595
transform 1 0 24932 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604681595
transform 1 0 26128 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604681595
transform 1 0 26680 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_276
timestamp 1604681595
transform 1 0 26496 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_280
timestamp 1604681595
transform 1 0 26864 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_271
timestamp 1604681595
transform 1 0 26036 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_288
timestamp 1604681595
transform 1 0 27600 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 28888 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_292
timestamp 1604681595
transform 1 0 27968 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_298
timestamp 1604681595
transform 1 0 28520 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_296
timestamp 1604681595
transform 1 0 28336 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1604681595
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1604681595
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_56
timestamp 1604681595
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_63
timestamp 1604681595
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_75
timestamp 1604681595
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_87
timestamp 1604681595
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1604681595
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_106
timestamp 1604681595
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1604681595
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1604681595
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_149
timestamp 1604681595
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1604681595
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_168
timestamp 1604681595
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_180
timestamp 1604681595
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_187
timestamp 1604681595
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_199
timestamp 1604681595
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_211
timestamp 1604681595
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_218
timestamp 1604681595
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23920 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_230
timestamp 1604681595
transform 1 0 22264 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_242
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1604681595
transform 1 0 24012 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1604681595
transform 1 0 25116 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 26772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1604681595
transform 1 0 26220 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_280
timestamp 1604681595
transform 1 0 26864 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 28888 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_292
timestamp 1604681595
transform 1 0 27968 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1604681595
transform 1 0 28520 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 27710 0 27766 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 4986 23520 5042 24000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 29182 0 29238 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 8298 23520 8354 24000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 2042 0 2098 480 6 bottom_grid_pin_0_
port 4 nsew default tristate
rlabel metal2 s 16302 0 16358 480 6 bottom_grid_pin_10_
port 5 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 bottom_grid_pin_11_
port 6 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 bottom_grid_pin_12_
port 7 nsew default tristate
rlabel metal2 s 20626 0 20682 480 6 bottom_grid_pin_13_
port 8 nsew default tristate
rlabel metal2 s 22006 0 22062 480 6 bottom_grid_pin_14_
port 9 nsew default tristate
rlabel metal2 s 23478 0 23534 480 6 bottom_grid_pin_15_
port 10 nsew default tristate
rlabel metal2 s 3514 0 3570 480 6 bottom_grid_pin_1_
port 11 nsew default tristate
rlabel metal2 s 4894 0 4950 480 6 bottom_grid_pin_2_
port 12 nsew default tristate
rlabel metal2 s 6366 0 6422 480 6 bottom_grid_pin_3_
port 13 nsew default tristate
rlabel metal2 s 7746 0 7802 480 6 bottom_grid_pin_4_
port 14 nsew default tristate
rlabel metal2 s 9218 0 9274 480 6 bottom_grid_pin_5_
port 15 nsew default tristate
rlabel metal2 s 10598 0 10654 480 6 bottom_grid_pin_6_
port 16 nsew default tristate
rlabel metal2 s 12070 0 12126 480 6 bottom_grid_pin_7_
port 17 nsew default tristate
rlabel metal2 s 13450 0 13506 480 6 bottom_grid_pin_8_
port 18 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 bottom_grid_pin_9_
port 19 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 bottom_width_0_height_0__pin_0_
port 20 nsew default input
rlabel metal2 s 26330 0 26386 480 6 bottom_width_0_height_0__pin_1_lower
port 21 nsew default tristate
rlabel metal2 s 662 0 718 480 6 bottom_width_0_height_0__pin_1_upper
port 22 nsew default tristate
rlabel metal2 s 11610 23520 11666 24000 6 ccff_head
port 23 nsew default input
rlabel metal2 s 14922 23520 14978 24000 6 ccff_tail
port 24 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[0]
port 25 nsew default input
rlabel metal3 s 0 18232 480 18352 6 chanx_left_in[10]
port 26 nsew default input
rlabel metal3 s 0 18776 480 18896 6 chanx_left_in[11]
port 27 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chanx_left_in[12]
port 28 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[13]
port 29 nsew default input
rlabel metal3 s 0 20544 480 20664 6 chanx_left_in[14]
port 30 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chanx_left_in[15]
port 31 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chanx_left_in[16]
port 32 nsew default input
rlabel metal3 s 0 22312 480 22432 6 chanx_left_in[17]
port 33 nsew default input
rlabel metal3 s 0 22992 480 23112 6 chanx_left_in[18]
port 34 nsew default input
rlabel metal3 s 0 23536 480 23656 6 chanx_left_in[19]
port 35 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[1]
port 36 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[2]
port 37 nsew default input
rlabel metal3 s 0 14016 480 14136 6 chanx_left_in[3]
port 38 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[4]
port 39 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chanx_left_in[5]
port 40 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[6]
port 41 nsew default input
rlabel metal3 s 0 16328 480 16448 6 chanx_left_in[7]
port 42 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chanx_left_in[8]
port 43 nsew default input
rlabel metal3 s 0 17552 480 17672 6 chanx_left_in[9]
port 44 nsew default input
rlabel metal3 s 0 280 480 400 6 chanx_left_out[0]
port 45 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[10]
port 46 nsew default tristate
rlabel metal3 s 0 6808 480 6928 6 chanx_left_out[11]
port 47 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[12]
port 48 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 chanx_left_out[13]
port 49 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_left_out[14]
port 50 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[15]
port 51 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[16]
port 52 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 chanx_left_out[17]
port 53 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[18]
port 54 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[19]
port 55 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[1]
port 56 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 57 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[3]
port 58 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[4]
port 59 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_out[5]
port 60 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[6]
port 61 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[7]
port 62 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[8]
port 63 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[9]
port 64 nsew default tristate
rlabel metal3 s 29520 12248 30000 12368 6 chanx_right_in[0]
port 65 nsew default input
rlabel metal3 s 29520 18232 30000 18352 6 chanx_right_in[10]
port 66 nsew default input
rlabel metal3 s 29520 18776 30000 18896 6 chanx_right_in[11]
port 67 nsew default input
rlabel metal3 s 29520 19320 30000 19440 6 chanx_right_in[12]
port 68 nsew default input
rlabel metal3 s 29520 20000 30000 20120 6 chanx_right_in[13]
port 69 nsew default input
rlabel metal3 s 29520 20544 30000 20664 6 chanx_right_in[14]
port 70 nsew default input
rlabel metal3 s 29520 21224 30000 21344 6 chanx_right_in[15]
port 71 nsew default input
rlabel metal3 s 29520 21768 30000 21888 6 chanx_right_in[16]
port 72 nsew default input
rlabel metal3 s 29520 22312 30000 22432 6 chanx_right_in[17]
port 73 nsew default input
rlabel metal3 s 29520 22992 30000 23112 6 chanx_right_in[18]
port 74 nsew default input
rlabel metal3 s 29520 23536 30000 23656 6 chanx_right_in[19]
port 75 nsew default input
rlabel metal3 s 29520 12792 30000 12912 6 chanx_right_in[1]
port 76 nsew default input
rlabel metal3 s 29520 13336 30000 13456 6 chanx_right_in[2]
port 77 nsew default input
rlabel metal3 s 29520 14016 30000 14136 6 chanx_right_in[3]
port 78 nsew default input
rlabel metal3 s 29520 14560 30000 14680 6 chanx_right_in[4]
port 79 nsew default input
rlabel metal3 s 29520 15240 30000 15360 6 chanx_right_in[5]
port 80 nsew default input
rlabel metal3 s 29520 15784 30000 15904 6 chanx_right_in[6]
port 81 nsew default input
rlabel metal3 s 29520 16328 30000 16448 6 chanx_right_in[7]
port 82 nsew default input
rlabel metal3 s 29520 17008 30000 17128 6 chanx_right_in[8]
port 83 nsew default input
rlabel metal3 s 29520 17552 30000 17672 6 chanx_right_in[9]
port 84 nsew default input
rlabel metal3 s 29520 280 30000 400 6 chanx_right_out[0]
port 85 nsew default tristate
rlabel metal3 s 29520 6264 30000 6384 6 chanx_right_out[10]
port 86 nsew default tristate
rlabel metal3 s 29520 6808 30000 6928 6 chanx_right_out[11]
port 87 nsew default tristate
rlabel metal3 s 29520 7352 30000 7472 6 chanx_right_out[12]
port 88 nsew default tristate
rlabel metal3 s 29520 8032 30000 8152 6 chanx_right_out[13]
port 89 nsew default tristate
rlabel metal3 s 29520 8576 30000 8696 6 chanx_right_out[14]
port 90 nsew default tristate
rlabel metal3 s 29520 9256 30000 9376 6 chanx_right_out[15]
port 91 nsew default tristate
rlabel metal3 s 29520 9800 30000 9920 6 chanx_right_out[16]
port 92 nsew default tristate
rlabel metal3 s 29520 10344 30000 10464 6 chanx_right_out[17]
port 93 nsew default tristate
rlabel metal3 s 29520 11024 30000 11144 6 chanx_right_out[18]
port 94 nsew default tristate
rlabel metal3 s 29520 11568 30000 11688 6 chanx_right_out[19]
port 95 nsew default tristate
rlabel metal3 s 29520 824 30000 944 6 chanx_right_out[1]
port 96 nsew default tristate
rlabel metal3 s 29520 1368 30000 1488 6 chanx_right_out[2]
port 97 nsew default tristate
rlabel metal3 s 29520 2048 30000 2168 6 chanx_right_out[3]
port 98 nsew default tristate
rlabel metal3 s 29520 2592 30000 2712 6 chanx_right_out[4]
port 99 nsew default tristate
rlabel metal3 s 29520 3272 30000 3392 6 chanx_right_out[5]
port 100 nsew default tristate
rlabel metal3 s 29520 3816 30000 3936 6 chanx_right_out[6]
port 101 nsew default tristate
rlabel metal3 s 29520 4360 30000 4480 6 chanx_right_out[7]
port 102 nsew default tristate
rlabel metal3 s 29520 5040 30000 5160 6 chanx_right_out[8]
port 103 nsew default tristate
rlabel metal3 s 29520 5584 30000 5704 6 chanx_right_out[9]
port 104 nsew default tristate
rlabel metal2 s 21638 23520 21694 24000 6 gfpga_pad_EMBEDDED_IO_SOC_DIR
port 105 nsew default tristate
rlabel metal2 s 24950 23520 25006 24000 6 gfpga_pad_EMBEDDED_IO_SOC_IN
port 106 nsew default input
rlabel metal2 s 28262 23520 28318 24000 6 gfpga_pad_EMBEDDED_IO_SOC_OUT
port 107 nsew default tristate
rlabel metal2 s 1674 23520 1730 24000 6 prog_clk
port 108 nsew default input
rlabel metal2 s 18326 23520 18382 24000 6 top_grid_pin_0_
port 109 nsew default tristate
rlabel metal4 s 5944 2128 6264 21808 6 VPWR
port 110 nsew default input
rlabel metal4 s 10944 2128 11264 21808 6 VGND
port 111 nsew default input
<< properties >>
string FIXED_BBOX 0 0 30000 24000
<< end >>
