* NGSPICE file created from cbx_1__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

.subckt cbx_1__1_ SC_IN_BOT SC_IN_TOP SC_OUT_BOT SC_OUT_TOP bottom_grid_pin_0_ bottom_grid_pin_10_
+ bottom_grid_pin_11_ bottom_grid_pin_12_ bottom_grid_pin_13_ bottom_grid_pin_14_
+ bottom_grid_pin_15_ bottom_grid_pin_1_ bottom_grid_pin_2_ bottom_grid_pin_3_ bottom_grid_pin_4_
+ bottom_grid_pin_5_ bottom_grid_pin_6_ bottom_grid_pin_7_ bottom_grid_pin_8_ bottom_grid_pin_9_
+ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12]
+ chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17]
+ chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11] chanx_right_out[12]
+ chanx_right_out[13] chanx_right_out[14] chanx_right_out[15] chanx_right_out[16]
+ chanx_right_out[17] chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chanx_right_out[9] prog_clk VPWR VGND
XANTENNA_mux_top_ipin_7.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_1__S mux_top_ipin_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_7.mux_l4_in_0_/S mux_top_ipin_8.mux_l1_in_1_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_26_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_12.mux_l2_in_0__A1 mux_top_ipin_12.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_13.mux_l3_in_0_ mux_top_ipin_13.mux_l2_in_1_/X mux_top_ipin_13.mux_l2_in_0_/X
+ mux_top_ipin_13.mux_l3_in_1_/S mux_top_ipin_13.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_66_ chanx_left_in[8] chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l2_in_2__A1 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_6.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_6.mux_l1_in_0_/X mux_top_ipin_6.mux_l2_in_3_/S
+ mux_top_ipin_6.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_0.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_7.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_5.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_2__S mux_top_ipin_5.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_49_ chanx_right_in[5] chanx_left_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xclkbuf_3_4_0_prog_clk clkbuf_2_2_0_prog_clk/X clkbuf_3_4_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_ipin_12.mux_l1_in_0__S mux_top_ipin_12.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_13.mux_l2_in_1_ chanx_left_in[9] chanx_right_in[3] mux_top_ipin_13.mux_l2_in_3_/S
+ mux_top_ipin_13.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_9.mux_l3_in_0__S mux_top_ipin_9.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l3_in_1__A1 mux_top_ipin_10.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_3__A1 chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l3_in_0__A1 mux_top_ipin_5.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.mux_l2_in_0__S mux_top_ipin_11.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_10.mux_l4_in_0__A1 mux_top_ipin_10.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_8.mux_l4_in_0__S mux_top_ipin_8.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_0.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_1.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_1.mux_l1_in_0_/S
+ mux_top_ipin_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_3.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_10.mux_l3_in_0__S mux_top_ipin_10.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_0.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_65_ chanx_left_in[9] chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_48_ chanx_right_in[6] chanx_left_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_0.mux_l3_in_0__A0 mux_top_ipin_0.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_13.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_13.mux_l1_in_0_/X mux_top_ipin_13.mux_l2_in_3_/S
+ mux_top_ipin_13.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_11.mux_l2_in_3__S mux_top_ipin_11.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_6.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_6.mux_l1_in_0_/S
+ mux_top_ipin_6.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_15.mux_l3_in_1__S mux_top_ipin_15.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_2.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_6.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_14.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_9.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_0.mux_l1_in_2__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_12.mux_l2_in_3__A0 _23_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_14.mux_l3_in_0__A0 mux_top_ipin_14.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_7.mux_l2_in_2__A0 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_0__S mux_top_ipin_7.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_14.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_0.mux_l2_in_1__A1 mux_top_ipin_0.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_64_ chanx_left_in[10] chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_4.mux_l4_in_0_/X bottom_grid_pin_4_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_7.mux_l3_in_1__A0 mux_top_ipin_7.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_9.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0__S mux_top_ipin_6.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_47_ chanx_right_in[7] chanx_left_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_0.mux_l3_in_0__A1 mux_top_ipin_0.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_1.mux_l2_in_2__S mux_top_ipin_1.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_7.mux_l4_in_0__A0 mux_top_ipin_7.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_5.mux_l3_in_0__S mux_top_ipin_5.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_13.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_13.mux_l1_in_0_/S
+ mux_top_ipin_13.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_9.mux_l2_in_0__A1 mux_top_ipin_9.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_12.mux_l2_in_3__A1 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_11.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l3_in_0__A1 mux_top_ipin_14.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l2_in_2__A1 chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_3__S mux_top_ipin_6.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l4_in_0__S mux_top_ipin_4.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_63_ chanx_left_in[11] chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l3_in_1__A1 mux_top_ipin_7.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_46_ chanx_right_in[8] chanx_left_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_12.mux_l2_in_1__S mux_top_ipin_12.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_4.mux_l2_in_0__A0 mux_top_ipin_4.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_29_ _29_/HI _29_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_ipin_7.mux_l4_in_0__A1 mux_top_ipin_7.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_3_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_11.mux_l4_in_0_/X bottom_grid_pin_11_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xclkbuf_3_3_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_10.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_11.mux_l3_in_1__S mux_top_ipin_11.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.mux_l2_in_2__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_11.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_11.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_2.mux_l2_in_3_ _27_/HI chanx_right_in[14] mux_top_ipin_2.mux_l2_in_1_/S
+ mux_top_ipin_2.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_2.mux_l3_in_1__A0 mux_top_ipin_2.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_62_ chanx_left_in[12] chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_3.mux_l1_in_0__S mux_top_ipin_3.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_5.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_2.mux_l4_in_0__A0 mux_top_ipin_2.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_13.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_45_ chanx_right_in[9] chanx_left_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_2.mux_l4_in_0_ mux_top_ipin_2.mux_l3_in_1_/X mux_top_ipin_2.mux_l3_in_0_/X
+ mux_top_ipin_2.mux_l4_in_0_/S mux_top_ipin_2.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_28_ _28_/HI _28_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_ipin_4.mux_l2_in_0__A1 mux_top_ipin_4.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0__S mux_top_ipin_2.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_7.mux_l2_in_3_ _16_/HI chanx_right_in[17] mux_top_ipin_7.mux_l2_in_0_/S
+ mux_top_ipin_7.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_9.mux_l2_in_3__A0 _18_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_2.mux_l3_in_1_ mux_top_ipin_2.mux_l2_in_3_/X mux_top_ipin_2.mux_l2_in_2_/X
+ mux_top_ipin_2.mux_l3_in_0_/S mux_top_ipin_2.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_8.mux_l1_in_1__S mux_top_ipin_8.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.mux_l2_in_2__A1 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_1.mux_l3_in_0__S mux_top_ipin_1.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_6.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_2.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[6] mux_top_ipin_2.mux_l2_in_1_/S
+ mux_top_ipin_2.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_7.mux_l2_in_1__S mux_top_ipin_7.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_7.mux_l4_in_0_ mux_top_ipin_7.mux_l3_in_1_/X mux_top_ipin_7.mux_l3_in_0_/X
+ mux_top_ipin_7.mux_l4_in_0_/S mux_top_ipin_7.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_2.mux_l3_in_1__A1 mux_top_ipin_2.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_61_ chanx_left_in[13] chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_2.mux_l2_in_3__S mux_top_ipin_2.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l4_in_0__S mux_top_ipin_0.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_7.mux_l3_in_1_ mux_top_ipin_7.mux_l2_in_3_/X mux_top_ipin_7.mux_l2_in_2_/X
+ mux_top_ipin_7.mux_l3_in_0_/S mux_top_ipin_7.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_2.mux_l4_in_0__A1 mux_top_ipin_2.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_44_ chanx_right_in[10] chanx_left_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l3_in_1__S mux_top_ipin_6.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_3_0_prog_clk_A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_27_ _27_/HI _27_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_top_ipin_7.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[11] mux_top_ipin_7.mux_l2_in_0_/S
+ mux_top_ipin_7.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_9.mux_l2_in_3__A1 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_2.mux_l3_in_0_ mux_top_ipin_2.mux_l2_in_1_/X mux_top_ipin_2.mux_l2_in_0_/X
+ mux_top_ipin_2.mux_l3_in_0_/S mux_top_ipin_2.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_8.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_14.mux_l2_in_3_ _25_/HI chanx_right_in[18] mux_top_ipin_14.mux_l2_in_0_/S
+ mux_top_ipin_14.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_13.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_2.mux_l2_in_1_ chanx_left_in[6] chanx_right_in[2] mux_top_ipin_2.mux_l2_in_1_/S
+ mux_top_ipin_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_13.mux_l2_in_2__S mux_top_ipin_13.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_11.mux_l2_in_2__A0 chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__42__A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
X_60_ chanx_left_in[14] chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_14.mux_l4_in_0_ mux_top_ipin_14.mux_l3_in_1_/X mux_top_ipin_14.mux_l3_in_0_/X
+ mux_top_ipin_14.mux_l4_in_0_/S mux_top_ipin_14.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_6.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_3_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_7.mux_l3_in_0_ mux_top_ipin_7.mux_l2_in_1_/X mux_top_ipin_7.mux_l2_in_0_/X
+ mux_top_ipin_7.mux_l3_in_0_/S mux_top_ipin_7.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA__37__A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_43_ chanx_right_in[11] chanx_left_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_11.mux_l3_in_1__A0 mux_top_ipin_11.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_7.mux_l4_in_0_/X bottom_grid_pin_7_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_9_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_4.mux_l2_in_3__A0 _29_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_14.mux_l3_in_1_ mux_top_ipin_14.mux_l2_in_3_/X mux_top_ipin_14.mux_l2_in_2_/X
+ mux_top_ipin_14.mux_l3_in_0_/S mux_top_ipin_14.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_6.mux_l3_in_0__A0 mux_top_ipin_6.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_26_ _26_/HI _26_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_top_ipin_7.mux_l2_in_1_ chanx_left_in[11] mux_top_ipin_7.mux_l1_in_2_/X mux_top_ipin_7.mux_l2_in_0_/S
+ mux_top_ipin_7.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_11.mux_l4_in_0__A0 mux_top_ipin_11.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__50__A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_13.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_14.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[10] mux_top_ipin_14.mux_l2_in_0_/S
+ mux_top_ipin_14.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__45__A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_13.mux_l2_in_0__A1 mux_top_ipin_13.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_7.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_top_ipin_7.mux_l1_in_2_/S
+ mux_top_ipin_7.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1__S mux_top_ipin_4.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_2.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_2.mux_l1_in_0_/X mux_top_ipin_2.mux_l2_in_1_/S
+ mux_top_ipin_2.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_11.mux_l2_in_2__A1 chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_8.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_6.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_1__S mux_top_ipin_3.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_1.mux_l3_in_1_/S mux_top_ipin_1.mux_l4_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__53__A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_42_ chanx_right_in[12] chanx_left_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_11.mux_l3_in_1__A1 mux_top_ipin_11.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_4.mux_l2_in_3__A1 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_14.mux_l3_in_0_ mux_top_ipin_14.mux_l2_in_1_/X mux_top_ipin_14.mux_l2_in_0_/X
+ mux_top_ipin_14.mux_l3_in_0_/S mux_top_ipin_14.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_6.mux_l3_in_0__A1 mux_top_ipin_6.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__48__A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_11.mux_l3_in_1_/S mux_top_ipin_11.mux_l4_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25_ _25_/HI _25_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_top_ipin_7.mux_l2_in_0_ mux_top_ipin_7.mux_l1_in_1_/X mux_top_ipin_7.mux_l1_in_0_/X
+ mux_top_ipin_7.mux_l2_in_0_/S mux_top_ipin_7.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_2.mux_l3_in_1__S mux_top_ipin_2.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_11.mux_l4_in_0__A1 mux_top_ipin_11.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_2_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l2_in_2__S mux_top_ipin_8.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_15.mux_l1_in_0__S mux_top_ipin_15.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_14.mux_l2_in_1_ chanx_left_in[10] chanx_right_in[2] mux_top_ipin_14.mux_l2_in_0_/S
+ mux_top_ipin_14.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_14.mux_l4_in_0_/X bottom_grid_pin_14_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__61__A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_7.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_7.mux_l1_in_2_/S
+ mux_top_ipin_7.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_1.mux_l2_in_1__A0 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__56__A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_4.mux_l3_in_0_/S mux_top_ipin_4.mux_l4_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_14.mux_l2_in_0__S mux_top_ipin_14.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_14.mux_l3_in_0_/S mux_top_ipin_14.mux_l4_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_1.mux_l3_in_0__A0 mux_top_ipin_1.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_2.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_2.mux_l1_in_0_/S
+ mux_top_ipin_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_15.mux_l1_in_2__A0 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_1.mux_l2_in_3_/S mux_top_ipin_1.mux_l3_in_1_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_14_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_41_ chanx_right_in[13] chanx_left_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_13.mux_l3_in_0__S mux_top_ipin_13.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__64__A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_11.mux_l2_in_2_/S mux_top_ipin_11.mux_l3_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24_ _24_/HI _24_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_15.mux_l2_in_1__A0 chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__59__A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_7.mux_l3_in_0_/S mux_top_ipin_7.mux_l4_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_13.mux_l2_in_3__A0 _24_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_14.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_14.mux_l1_in_0_/X mux_top_ipin_14.mux_l2_in_0_/S
+ mux_top_ipin_14.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_14.mux_l2_in_3__S mux_top_ipin_14.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_12.mux_l4_in_0__S mux_top_ipin_12.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_0.mux_l4_in_0_/X bottom_grid_pin_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_15.mux_l3_in_0__A0 mux_top_ipin_15.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_7.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_7.mux_l1_in_2_/S
+ mux_top_ipin_7.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_8.mux_l2_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_3_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_14.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_4.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_1.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_4.mux_l2_in_0_/S mux_top_ipin_4.mux_l3_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__72__A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1__S mux_top_ipin_0.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__67__A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l3_in_1__A0 mux_top_ipin_8.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_14.mux_l2_in_0_/S mux_top_ipin_14.mux_l3_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_1.mux_l3_in_0__A1 mux_top_ipin_1.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_15.mux_l1_in_2__A1 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_1.mux_l1_in_0_/S mux_top_ipin_1.mux_l2_in_3_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_22_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_40_ chanx_right_in[14] chanx_left_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l4_in_0__A0 mux_top_ipin_8.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_11.mux_l1_in_2_/S mux_top_ipin_11.mux_l2_in_2_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_15.mux_l2_in_1__A1 mux_top_ipin_15.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_23_ _23_/HI _23_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_5.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_15.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_7.mux_l2_in_0_/S mux_top_ipin_7.mux_l3_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_9.mux_l2_in_0__S mux_top_ipin_9.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_13.mux_l2_in_3__A1 chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_12.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_15.mux_l3_in_0__A1 mux_top_ipin_15.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_8.mux_l2_in_2__A1 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_4.mux_l2_in_2__S mux_top_ipin_4.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_11.mux_l1_in_0__S mux_top_ipin_11.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_4.mux_l1_in_0_/S mux_top_ipin_4.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_14.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_14.mux_l1_in_0_/S
+ mux_top_ipin_14.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_8.mux_l3_in_0__S mux_top_ipin_8.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_8.mux_l3_in_1__A1 mux_top_ipin_8.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_14.mux_l1_in_0_/S mux_top_ipin_14.mux_l2_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0_prog_clk clkbuf_2_0_0_prog_clk/X clkbuf_3_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_23_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_0.mux_l4_in_0_/S mux_top_ipin_1.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_10.mux_l2_in_1__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l2_in_0__S mux_top_ipin_10.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_9.mux_l2_in_3__S mux_top_ipin_9.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_7.mux_l4_in_0__S mux_top_ipin_7.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l4_in_0__A1 mux_top_ipin_8.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_10.mux_l4_in_0_/S mux_top_ipin_11.mux_l1_in_2_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_10.mux_l3_in_0__A0 mux_top_ipin_10.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_22_ _22_/HI _22_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_ipin_3.mux_l2_in_2__A0 chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_7.mux_l1_in_2_/S mux_top_ipin_7.mux_l2_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_15.mux_l2_in_1__S mux_top_ipin_15.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_12.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l3_in_1__A0 mux_top_ipin_3.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_10.mux_l2_in_3__S mux_top_ipin_10.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_3.mux_l4_in_0_/S mux_top_ipin_4.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_16_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_14.mux_l3_in_1__S mux_top_ipin_14.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_3.mux_l4_in_0__A0 mux_top_ipin_3.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_13.mux_l4_in_0_/S mux_top_ipin_14.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_3.mux_l2_in_3_ _28_/HI chanx_right_in[19] mux_top_ipin_3.mux_l2_in_3_/S
+ mux_top_ipin_3.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_10.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_12.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_2.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_5.mux_l2_in_0__A1 mux_top_ipin_5.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_21_ _21_/HI _21_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_10.mux_l3_in_0__A1 mux_top_ipin_10.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0__S mux_top_ipin_6.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_3.mux_l2_in_2__A1 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_6.mux_l4_in_0_/S mux_top_ipin_7.mux_l1_in_2_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_3.mux_l4_in_0_ mux_top_ipin_3.mux_l3_in_1_/X mux_top_ipin_3.mux_l3_in_0_/X
+ mux_top_ipin_3.mux_l4_in_0_/S mux_top_ipin_3.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_3.mux_l3_in_1__A1 mux_top_ipin_3.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0__S mux_top_ipin_5.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_8.mux_l2_in_3_ _17_/HI chanx_right_in[18] mux_top_ipin_8.mux_l2_in_0_/S
+ mux_top_ipin_8.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_3.mux_l3_in_1_ mux_top_ipin_3.mux_l2_in_3_/X mux_top_ipin_3.mux_l2_in_2_/X
+ mux_top_ipin_3.mux_l3_in_1_/S mux_top_ipin_3.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_0.mux_l2_in_2__S mux_top_ipin_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l4_in_0__A1 mux_top_ipin_3.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0__A0 mux_top_ipin_0.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_4.mux_l3_in_0__S mux_top_ipin_4.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_3.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[13] mux_top_ipin_3.mux_l2_in_3_/S
+ mux_top_ipin_3.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_8.mux_l4_in_0_ mux_top_ipin_8.mux_l3_in_1_/X mux_top_ipin_8.mux_l3_in_0_/X
+ mux_top_ipin_8.mux_l4_in_0_/S mux_top_ipin_8.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_10.mux_l2_in_3_ _21_/HI chanx_right_in[14] mux_top_ipin_10.mux_l2_in_3_/S
+ mux_top_ipin_10.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20_ _20_/HI _20_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_5.mux_l2_in_3__S mux_top_ipin_5.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_9.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l4_in_0__S mux_top_ipin_3.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_12.mux_l1_in_1__S mux_top_ipin_12.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_8.mux_l3_in_1_ mux_top_ipin_8.mux_l2_in_3_/X mux_top_ipin_8.mux_l2_in_2_/X
+ mux_top_ipin_8.mux_l3_in_1_/S mux_top_ipin_8.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_9.mux_l3_in_1__S mux_top_ipin_9.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_2.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_7.mux_l1_in_2__A0 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_4_0_prog_clk_A clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_10.mux_l4_in_0_ mux_top_ipin_10.mux_l3_in_1_/X mux_top_ipin_10.mux_l3_in_0_/X
+ mux_top_ipin_10.mux_l4_in_0_/S mux_top_ipin_10.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_3.mux_l4_in_0_/X bottom_grid_pin_3_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_top_ipin_8.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[12] mux_top_ipin_8.mux_l2_in_0_/S
+ mux_top_ipin_8.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_12.mux_l2_in_2__A0 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_11.mux_l2_in_1__S mux_top_ipin_11.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_3.mux_l3_in_0_ mux_top_ipin_3.mux_l2_in_1_/X mux_top_ipin_3.mux_l2_in_0_/X
+ mux_top_ipin_3.mux_l3_in_1_/S mux_top_ipin_3.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_7.mux_l2_in_1__A0 chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_15.mux_l2_in_3_ _26_/HI chanx_right_in[19] mux_top_ipin_15.mux_l2_in_3_/S
+ mux_top_ipin_15.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_0.mux_l2_in_0__A1 mux_top_ipin_0.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_10.mux_l3_in_1_ mux_top_ipin_10.mux_l2_in_3_/X mux_top_ipin_10.mux_l2_in_2_/X
+ mux_top_ipin_10.mux_l3_in_1_/S mux_top_ipin_10.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_12.mux_l3_in_1__A0 mux_top_ipin_12.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_5.mux_l2_in_3__A0 _30_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_3.mux_l2_in_1_ chanx_left_in[13] mux_top_ipin_3.mux_l1_in_2_/X mux_top_ipin_3.mux_l2_in_3_/S
+ mux_top_ipin_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_10.mux_l3_in_1__S mux_top_ipin_10.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l3_in_0__A0 mux_top_ipin_7.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_5.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_10.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[6] mux_top_ipin_10.mux_l2_in_3_/S
+ mux_top_ipin_10.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_12.mux_l4_in_0__A0 mux_top_ipin_12.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_prog_clk clkbuf_2_0_0_prog_clk/X clkbuf_3_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_24_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_15.mux_l4_in_0_ mux_top_ipin_15.mux_l3_in_1_/X mux_top_ipin_15.mux_l3_in_0_/X
+ ccff_tail mux_top_ipin_15.mux_l4_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_3.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_top_ipin_3.mux_l1_in_2_/S
+ mux_top_ipin_3.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_3.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_13.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_9.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_8.mux_l3_in_0_ mux_top_ipin_8.mux_l2_in_1_/X mux_top_ipin_8.mux_l2_in_0_/X
+ mux_top_ipin_8.mux_l3_in_1_/S mux_top_ipin_8.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_14.mux_l2_in_0__A1 mux_top_ipin_14.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_7.mux_l1_in_2__A1 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_2.mux_l1_in_0__S mux_top_ipin_2.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_15.mux_l3_in_1_ mux_top_ipin_15.mux_l2_in_3_/X mux_top_ipin_15.mux_l2_in_2_/X
+ mux_top_ipin_15.mux_l3_in_1_/S mux_top_ipin_15.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_8.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_8.mux_l1_in_2_/X mux_top_ipin_8.mux_l2_in_0_/S
+ mux_top_ipin_8.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_12.mux_l2_in_2__A1 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_7.mux_l2_in_1__A1 mux_top_ipin_7.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_15.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[15] mux_top_ipin_15.mux_l2_in_3_/S
+ mux_top_ipin_15.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_8.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0__S mux_top_ipin_1.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_10.mux_l3_in_0_ mux_top_ipin_10.mux_l2_in_1_/X mux_top_ipin_10.mux_l2_in_0_/X
+ mux_top_ipin_10.mux_l3_in_1_/S mux_top_ipin_10.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_12.mux_l3_in_1__A1 mux_top_ipin_12.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_8.mux_l1_in_2_ chanx_right_in[8] chanx_left_in[8] mux_top_ipin_8.mux_l1_in_1_/S
+ mux_top_ipin_8.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_7.mux_l1_in_1__S mux_top_ipin_7.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_14.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_3__A1 chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_3.mux_l2_in_0_ mux_top_ipin_3.mux_l1_in_1_/X mux_top_ipin_3.mux_l1_in_0_/X
+ mux_top_ipin_3.mux_l2_in_3_/S mux_top_ipin_3.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_10.mux_l4_in_0_/X bottom_grid_pin_10_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_13_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_4.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_7.mux_l3_in_0__A1 mux_top_ipin_7.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_10.mux_l2_in_1_ chanx_left_in[6] chanx_right_in[2] mux_top_ipin_10.mux_l2_in_3_/S
+ mux_top_ipin_10.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_12.mux_l4_in_0__A1 mux_top_ipin_12.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_0.mux_l3_in_0__S mux_top_ipin_0.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_3.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_3.mux_l1_in_2_/S
+ mux_top_ipin_3.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_6.mux_l2_in_1__S mux_top_ipin_6.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_9.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_15.mux_l3_in_0_ mux_top_ipin_15.mux_l2_in_1_/X mux_top_ipin_15.mux_l2_in_0_/X
+ mux_top_ipin_15.mux_l3_in_1_/S mux_top_ipin_15.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_1.mux_l2_in_3__S mux_top_ipin_1.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.mux_l2_in_1__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_8.mux_l2_in_0_ mux_top_ipin_8.mux_l1_in_1_/X mux_top_ipin_8.mux_l1_in_0_/X
+ mux_top_ipin_8.mux_l2_in_0_/S mux_top_ipin_8.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_5.mux_l3_in_1__S mux_top_ipin_5.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_0.mux_l2_in_3__A0 _19_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_15.mux_l2_in_1_ chanx_left_in[15] mux_top_ipin_15.mux_l1_in_2_/X mux_top_ipin_15.mux_l2_in_3_/S
+ mux_top_ipin_15.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_2.mux_l3_in_0__A0 mux_top_ipin_2.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_8.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_8.mux_l1_in_1_/S
+ mux_top_ipin_8.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_15.mux_l1_in_2_ chanx_right_in[9] chanx_left_in[9] mux_top_ipin_15.mux_l1_in_1_/S
+ mux_top_ipin_15.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_10.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_10.mux_l1_in_0_/X mux_top_ipin_10.mux_l2_in_3_/S
+ mux_top_ipin_10.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_3.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_3.mux_l1_in_2_/S
+ mux_top_ipin_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_14.mux_l2_in_3__A0 _25_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_12.mux_l2_in_2__S mux_top_ipin_12.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_9.mux_l2_in_2__A0 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_2.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_9.mux_l3_in_1__A0 mux_top_ipin_9.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_3__A1 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_11.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_15.mux_l2_in_0_ mux_top_ipin_15.mux_l1_in_1_/X mux_top_ipin_15.mux_l1_in_0_/X
+ mux_top_ipin_15.mux_l2_in_3_/S mux_top_ipin_15.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_2.mux_l3_in_0__A1 mux_top_ipin_2.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_15.mux_l4_in_0__S ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_12.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_8.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_8.mux_l1_in_1_/S
+ mux_top_ipin_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_9.mux_l4_in_0__A0 mux_top_ipin_9.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_15.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_15.mux_l1_in_1_/S
+ mux_top_ipin_15.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_3.mux_l1_in_1__S mux_top_ipin_3.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_14.mux_l2_in_3__A1 chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_10.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_10.mux_l1_in_0_/S
+ mux_top_ipin_10.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_9.mux_l2_in_2__A1 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_59_ chanx_left_in[15] chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_2.mux_l2_in_1__S mux_top_ipin_2.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_15.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.mux_l1_in_2__A0 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l1_in_2__S mux_top_ipin_8.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_9.mux_l3_in_1__A1 mux_top_ipin_9.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_6.mux_l4_in_0_/X bottom_grid_pin_6_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_11_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_11.mux_l2_in_1__A0 chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l3_in_1__S mux_top_ipin_1.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_3_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__32__A SC_IN_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_2__S mux_top_ipin_7.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_9.mux_l4_in_0__A1 mux_top_ipin_9.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_14.mux_l1_in_0__S mux_top_ipin_14.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_15.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_15.mux_l1_in_1_/S
+ mux_top_ipin_15.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_11.mux_l3_in_0__A0 mux_top_ipin_11.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_4.mux_l2_in_2__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_3_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l2_in_0__S mux_top_ipin_13.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__40__A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_4.mux_l3_in_1__A0 mux_top_ipin_4.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_58_ chanx_left_in[16] chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_11.mux_l1_in_2__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__35__A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_12.mux_l3_in_0__S mux_top_ipin_12.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l4_in_0__A0 mux_top_ipin_4.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_11.mux_l2_in_1__A1 mux_top_ipin_11.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_12.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_2.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0__A1 mux_top_ipin_6.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l2_in_3__S mux_top_ipin_13.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_11.mux_l4_in_0__S mux_top_ipin_11.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__43__A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_13.mux_l4_in_0_/X bottom_grid_pin_13_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_ipin_11.mux_l3_in_0__A1 mux_top_ipin_11.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l2_in_2__A1 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__38__A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_74_ chanx_left_in[0] chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_3_ _29_/HI chanx_right_in[14] mux_top_ipin_4.mux_l2_in_0_/S
+ mux_top_ipin_4.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_4.mux_l3_in_1__A1 mux_top_ipin_4.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_57_ chanx_left_in[17] chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__51__A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_3.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_13.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_9.mux_l1_in_0__S mux_top_ipin_9.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_1.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l4_in_0__A1 mux_top_ipin_4.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__46__A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l4_in_0_ mux_top_ipin_4.mux_l3_in_1_/X mux_top_ipin_4.mux_l3_in_0_/X
+ mux_top_ipin_4.mux_l4_in_0_/S mux_top_ipin_4.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_0.mux_l3_in_1_/S mux_top_ipin_0.mux_l4_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_4.mux_l1_in_2__S mux_top_ipin_4.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_9.mux_l2_in_3_ _18_/HI chanx_right_in[13] mux_top_ipin_9.mux_l2_in_2_/S
+ mux_top_ipin_9.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_8.mux_l2_in_0__S mux_top_ipin_8.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_10.mux_l3_in_1_/S mux_top_ipin_10.mux_l4_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_15.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_4.mux_l3_in_1_ mux_top_ipin_4.mux_l2_in_3_/X mux_top_ipin_4.mux_l2_in_2_/X
+ mux_top_ipin_4.mux_l3_in_0_/S mux_top_ipin_4.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_3.mux_l2_in_2__S mux_top_ipin_3.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_prog_clk_A clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_10.mux_l1_in_0__S mux_top_ipin_10.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__54__A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_73_ chanx_left_in[1] chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_15.mux_l2_in_0__A0 mux_top_ipin_15.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_7.mux_l3_in_0__S mux_top_ipin_7.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[8] mux_top_ipin_4.mux_l2_in_0_/S
+ mux_top_ipin_4.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_8.mux_l1_in_2__A0 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_9.mux_l4_in_0_ mux_top_ipin_9.mux_l3_in_1_/X mux_top_ipin_9.mux_l3_in_0_/X
+ mux_top_ipin_9.mux_l4_in_0_/S mux_top_ipin_9.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__49__A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_3.mux_l3_in_1_/S mux_top_ipin_3.mux_l4_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_56_ chanx_left_in[18] chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_13.mux_l2_in_2__A0 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_11.mux_l2_in_3_ _22_/HI chanx_right_in[15] mux_top_ipin_11.mux_l2_in_2_/S
+ mux_top_ipin_11.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_8.mux_l2_in_1__A0 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_8.mux_l2_in_3__S mux_top_ipin_8.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l4_in_0__S mux_top_ipin_6.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_9.mux_l3_in_1_ mux_top_ipin_9.mux_l2_in_3_/X mux_top_ipin_9.mux_l2_in_2_/X
+ mux_top_ipin_9.mux_l3_in_1_/S mux_top_ipin_9.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_39_ chanx_right_in[15] chanx_left_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_15.mux_l1_in_1__S mux_top_ipin_15.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_13.mux_l3_in_1_/S mux_top_ipin_13.mux_l4_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_1.mux_l2_in_0__A1 mux_top_ipin_1.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_3_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_13.mux_l3_in_1__A0 mux_top_ipin_13.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_0.mux_l2_in_3_/S mux_top_ipin_0.mux_l3_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__62__A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_6.mux_l2_in_3__A0 _31_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_5_0_prog_clk_A clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_8.mux_l3_in_0__A0 mux_top_ipin_8.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_11.mux_l4_in_0_ mux_top_ipin_11.mux_l3_in_1_/X mux_top_ipin_11.mux_l3_in_0_/X
+ mux_top_ipin_11.mux_l4_in_0_/S mux_top_ipin_11.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA__57__A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_9.mux_l2_in_2_ chanx_left_in[13] chanx_right_in[5] mux_top_ipin_9.mux_l2_in_2_/S
+ mux_top_ipin_9.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_10.mux_l2_in_3_/S mux_top_ipin_10.mux_l3_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_15.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l2_in_1__S mux_top_ipin_14.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l3_in_0_ mux_top_ipin_4.mux_l2_in_1_/X mux_top_ipin_4.mux_l2_in_0_/X
+ mux_top_ipin_4.mux_l3_in_0_/S mux_top_ipin_4.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_13.mux_l4_in_0__A0 mux_top_ipin_13.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_6.mux_l3_in_1_/S mux_top_ipin_6.mux_l4_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_11.mux_l3_in_1_ mux_top_ipin_11.mux_l2_in_3_/X mux_top_ipin_11.mux_l2_in_2_/X
+ mux_top_ipin_11.mux_l3_in_1_/S mux_top_ipin_11.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA__70__A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_72_ chanx_left_in[2] chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_15.mux_l2_in_0__A1 mux_top_ipin_15.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l2_in_1_ chanx_left_in[8] mux_top_ipin_4.mux_l1_in_2_/X mux_top_ipin_4.mux_l2_in_0_/S
+ mux_top_ipin_4.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_13.mux_l3_in_1__S mux_top_ipin_13.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l1_in_2__A1 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__65__A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_3.mux_l2_in_3_/S mux_top_ipin_3.mux_l3_in_1_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_13.mux_l2_in_2__A1 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_11.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[11] mux_top_ipin_11.mux_l2_in_2_/S
+ mux_top_ipin_11.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_55_ chanx_left_in[19] chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_4.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_4.mux_l1_in_0_/S
+ mux_top_ipin_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_8.mux_l2_in_1__A1 mux_top_ipin_8.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_9.mux_l3_in_0_ mux_top_ipin_9.mux_l2_in_1_/X mux_top_ipin_9.mux_l2_in_0_/X
+ mux_top_ipin_9.mux_l3_in_1_/S mux_top_ipin_9.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_13.mux_l2_in_3_/S mux_top_ipin_13.mux_l3_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_38_ chanx_right_in[16] chanx_left_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_13.mux_l3_in_1__A1 mux_top_ipin_13.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_0.mux_l1_in_2_/S mux_top_ipin_0.mux_l2_in_3_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_6.mux_l2_in_3__A1 chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0__S mux_top_ipin_5.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_9.mux_l3_in_1_/S mux_top_ipin_9.mux_l4_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_9.mux_l4_in_0_/X bottom_grid_pin_9_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_15.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_5.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l3_in_0__A1 mux_top_ipin_8.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__73__A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_9.mux_l2_in_1_ chanx_left_in[5] chanx_right_in[3] mux_top_ipin_9.mux_l2_in_2_/S
+ mux_top_ipin_9.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_10.mux_l1_in_0_/S mux_top_ipin_10.mux_l2_in_3_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_10.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l4_in_0__A1 mux_top_ipin_13.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_2__S mux_top_ipin_0.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_2__A0 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__68__A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_6.mux_l2_in_3_/S mux_top_ipin_6.mux_l3_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l2_in_0__S mux_top_ipin_4.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_11.mux_l3_in_0_ mux_top_ipin_11.mux_l2_in_1_/X mux_top_ipin_11.mux_l2_in_0_/X
+ mux_top_ipin_11.mux_l3_in_1_/S mux_top_ipin_11.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_71_ chanx_left_in[3] chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_0_ mux_top_ipin_4.mux_l1_in_1_/X mux_top_ipin_4.mux_l1_in_0_/X
+ mux_top_ipin_4.mux_l2_in_0_/S mux_top_ipin_4.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_3.mux_l2_in_1__A0 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_3.mux_l1_in_2_/S mux_top_ipin_3.mux_l2_in_3_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_54_ chanx_right_in[0] chanx_left_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_11.mux_l2_in_1_ chanx_left_in[11] mux_top_ipin_11.mux_l1_in_2_/X mux_top_ipin_11.mux_l2_in_2_/S
+ mux_top_ipin_11.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l3_in_0__S mux_top_ipin_3.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_3__A0 _20_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_4.mux_l1_in_0_/S
+ mux_top_ipin_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_9.mux_l2_in_1__S mux_top_ipin_9.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_3.mux_l3_in_0__A0 mux_top_ipin_3.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_13.mux_l1_in_0_/S mux_top_ipin_13.mux_l2_in_3_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_37_ chanx_right_in[17] chanx_left_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_28_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ ccff_head mux_top_ipin_0.mux_l1_in_2_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_11.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_11.mux_l1_in_2_/S
+ mux_top_ipin_11.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_9.mux_l2_in_2_/S mux_top_ipin_9.mux_l3_in_1_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_4.mux_l2_in_3__S mux_top_ipin_4.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_2.mux_l4_in_0__S mux_top_ipin_2.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.mux_l1_in_1__S mux_top_ipin_11.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_9.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_9.mux_l1_in_0_/X mux_top_ipin_9.mux_l2_in_2_/S
+ mux_top_ipin_9.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_9.mux_l4_in_0_/S mux_top_ipin_10.mux_l1_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_8.mux_l3_in_1__S mux_top_ipin_8.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l2_in_0__A1 mux_top_ipin_10.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_3.mux_l1_in_2__A1 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_6.mux_l1_in_0_/S mux_top_ipin_6.mux_l2_in_3_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_15.mux_l2_in_3__A0 _26_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l2_in_1__S mux_top_ipin_10.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_70_ chanx_left_in[4] chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_3.mux_l2_in_1__A1 mux_top_ipin_3.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_2.mux_l4_in_0_/S mux_top_ipin_3.mux_l1_in_2_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_53_ chanx_right_in[1] chanx_left_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_11.mux_l2_in_0_ mux_top_ipin_11.mux_l1_in_1_/X mux_top_ipin_11.mux_l1_in_0_/X
+ mux_top_ipin_11.mux_l2_in_2_/S mux_top_ipin_11.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_1.mux_l2_in_3__A1 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_4.mux_l1_in_0_/S
+ mux_top_ipin_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_11.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_3_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l3_in_0__A1 mux_top_ipin_3.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_36_ chanx_right_in[18] chanx_left_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_12.mux_l4_in_0_/S mux_top_ipin_13.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_15.mux_l2_in_2__S mux_top_ipin_15.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_11.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_11.mux_l1_in_2_/S
+ mux_top_ipin_11.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_9.mux_l1_in_0_/S mux_top_ipin_9.mux_l2_in_2_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_19_ _19_/HI _19_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_1.mux_l1_in_0__S mux_top_ipin_1.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_5.mux_l4_in_0_/S mux_top_ipin_6.mux_l1_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_15.mux_l2_in_3__A1 chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_2.mux_l4_in_0_/X bottom_grid_pin_2_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_top_ipin_9.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_9.mux_l1_in_0_/S
+ mux_top_ipin_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_12.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_2.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_0.mux_l2_in_0__S mux_top_ipin_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_12.mux_l1_in_2__A0 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_52_ chanx_right_in[2] chanx_left_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_0.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35_ chanx_right_in[19] chanx_left_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_12.mux_l2_in_1__A0 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_7.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_11.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_11.mux_l1_in_2_/S
+ mux_top_ipin_11.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0__A0 mux_top_ipin_7.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_5.mux_l2_in_1__S mux_top_ipin_5.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_18_ _18_/HI _18_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_8.mux_l4_in_0_/S mux_top_ipin_9.mux_l1_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_10.mux_l2_in_3__A0 _21_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_12.mux_l3_in_0__A0 mux_top_ipin_12.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_5.mux_l2_in_2__A0 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_0.mux_l2_in_3__S mux_top_ipin_0.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_1.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l3_in_1__S mux_top_ipin_4.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_5.mux_l3_in_1__A0 mux_top_ipin_5.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_12.mux_l1_in_2__A1 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_51_ chanx_right_in[3] chanx_left_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_7.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_12.mux_l1_in_2__S mux_top_ipin_12.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_5.mux_l4_in_0__A0 mux_top_ipin_5.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_34_ _34_/A SC_OUT_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_12.mux_l2_in_1__A1 mux_top_ipin_12.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0__A1 mux_top_ipin_7.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17_ _17_/HI _17_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_18_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_4.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l2_in_3__A1 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.mux_l2_in_2__S mux_top_ipin_11.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_12.mux_l3_in_0__A1 mux_top_ipin_12.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_15.mux_l3_in_0__S mux_top_ipin_15.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l2_in_3_ _19_/HI chanx_right_in[16] mux_top_ipin_0.mux_l2_in_3_/S
+ mux_top_ipin_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_5.mux_l2_in_2__A1 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_5.mux_l3_in_1__A1 mux_top_ipin_5.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l4_in_0__S mux_top_ipin_14.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_0.mux_l4_in_0_ mux_top_ipin_0.mux_l3_in_1_/X mux_top_ipin_0.mux_l3_in_0_/X
+ mux_top_ipin_0.mux_l4_in_0_/S mux_top_ipin_0.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_50_ chanx_right_in[4] chanx_left_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l4_in_0__A1 mux_top_ipin_5.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_7.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_5.mux_l2_in_3_ _30_/HI chanx_right_in[17] mux_top_ipin_5.mux_l2_in_3_/S
+ mux_top_ipin_5.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_33_ _33_/A SC_OUT_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_0.mux_l3_in_1_ mux_top_ipin_0.mux_l2_in_3_/X mux_top_ipin_0.mux_l2_in_2_/X
+ mux_top_ipin_0.mux_l3_in_1_/S mux_top_ipin_0.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_0.mux_l2_in_2__A0 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16_ _16_/HI _16_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_18_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_8.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_top_ipin_0.mux_l2_in_3_/S
+ mux_top_ipin_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_0.mux_l3_in_1__A0 mux_top_ipin_0.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_5.mux_l4_in_0_ mux_top_ipin_5.mux_l3_in_1_/X mux_top_ipin_5.mux_l3_in_0_/X
+ mux_top_ipin_5.mux_l4_in_0_/S mux_top_ipin_5.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_1.mux_l2_in_1__S mux_top_ipin_1.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_7.mux_l1_in_2__S mux_top_ipin_7.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_7_0_prog_clk clkbuf_3_6_0_prog_clk/A clkbuf_3_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_0.mux_l4_in_0__A0 mux_top_ipin_0.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l2_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_5.mux_l3_in_1_ mux_top_ipin_5.mux_l2_in_3_/X mux_top_ipin_5.mux_l2_in_2_/X
+ mux_top_ipin_5.mux_l3_in_1_/S mux_top_ipin_5.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_0.mux_l3_in_1__S mux_top_ipin_0.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_9.mux_l2_in_1__A0 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_6.mux_l2_in_2__S mux_top_ipin_6.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_prog_clk_A clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l1_in_0__S mux_top_ipin_13.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0__A1 mux_top_ipin_2.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_14.mux_l3_in_1__A0 mux_top_ipin_14.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_32_ SC_IN_BOT SC_IN_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_5.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[9] mux_top_ipin_5.mux_l2_in_3_/S
+ mux_top_ipin_5.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_9.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_7.mux_l2_in_3__A0 _16_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l3_in_0_ mux_top_ipin_0.mux_l2_in_1_/X mux_top_ipin_0.mux_l2_in_0_/X
+ mux_top_ipin_0.mux_l3_in_1_/S mux_top_ipin_0.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_9.mux_l3_in_0__A0 mux_top_ipin_9.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_12.mux_l2_in_3_ _23_/HI chanx_right_in[16] mux_top_ipin_12.mux_l2_in_2_/S
+ mux_top_ipin_12.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_12.mux_l2_in_0__S mux_top_ipin_12.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l4_in_0__A0 mux_top_ipin_14.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_9.mux_l4_in_0__S mux_top_ipin_9.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_0.mux_l2_in_1_ chanx_left_in[10] mux_top_ipin_0.mux_l1_in_2_/X mux_top_ipin_0.mux_l2_in_3_/S
+ mux_top_ipin_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l3_in_1__A1 mux_top_ipin_0.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_6_0_prog_clk_A clkbuf_3_6_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_11.mux_l3_in_0__S mux_top_ipin_11.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_12.mux_l4_in_0_ mux_top_ipin_12.mux_l3_in_1_/X mux_top_ipin_12.mux_l3_in_0_/X
+ mux_top_ipin_12.mux_l4_in_0_/S mux_top_ipin_12.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_10.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_0.mux_l1_in_2_/S
+ mux_top_ipin_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_0.mux_l4_in_0__A1 mux_top_ipin_0.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_5.mux_l3_in_0_ mux_top_ipin_5.mux_l2_in_1_/X mux_top_ipin_5.mux_l2_in_0_/X
+ mux_top_ipin_5.mux_l3_in_1_/S mux_top_ipin_5.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_5.mux_l4_in_0_/X bottom_grid_pin_5_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_9.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_12.mux_l3_in_1_ mux_top_ipin_12.mux_l2_in_3_/X mux_top_ipin_12.mux_l2_in_2_/X
+ mux_top_ipin_12.mux_l3_in_0_/S mux_top_ipin_12.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_12.mux_l2_in_3__S mux_top_ipin_12.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_10.mux_l4_in_0__S mux_top_ipin_10.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_11.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l3_in_1__A1 mux_top_ipin_14.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_5.mux_l2_in_1_ chanx_left_in[9] chanx_right_in[3] mux_top_ipin_5.mux_l2_in_3_/S
+ mux_top_ipin_5.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_31_ _31_/HI _31_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_7.mux_l2_in_3__A1 chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_9.mux_l3_in_0__A1 mux_top_ipin_9.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_12.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[12] mux_top_ipin_12.mux_l2_in_2_/S
+ mux_top_ipin_12.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_11.mux_l2_in_0__A0 mux_top_ipin_11.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l4_in_0__A1 mux_top_ipin_14.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_1.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_11.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_0.mux_l2_in_0_ mux_top_ipin_0.mux_l1_in_1_/X mux_top_ipin_0.mux_l1_in_0_/X
+ mux_top_ipin_0.mux_l2_in_3_/S mux_top_ipin_0.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_8.mux_l1_in_0__S mux_top_ipin_8.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_1__A0 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_3_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0__A mux_top_ipin_14.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_0.mux_l1_in_2_/S
+ mux_top_ipin_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_3.mux_l1_in_2__S mux_top_ipin_3.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_2.mux_l2_in_3__A0 _27_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l3_in_0__A0 mux_top_ipin_4.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0__S mux_top_ipin_7.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_12.mux_l3_in_0_ mux_top_ipin_12.mux_l2_in_1_/X mux_top_ipin_12.mux_l2_in_0_/X
+ mux_top_ipin_12.mux_l3_in_0_/S mux_top_ipin_12.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_11.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_5.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_5.mux_l1_in_0_/X mux_top_ipin_5.mux_l2_in_3_/S
+ mux_top_ipin_5.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_30_ _30_/HI _30_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_28_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_12.mux_l4_in_0_/X bottom_grid_pin_12_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_ipin_6.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_0_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.mux_l2_in_2__S mux_top_ipin_2.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_12.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_12.mux_l1_in_2_/X mux_top_ipin_12.mux_l2_in_2_/S
+ mux_top_ipin_12.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_6.mux_l3_in_0__S mux_top_ipin_6.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.mux_l2_in_0__A1 mux_top_ipin_11.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_2__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_12.mux_l1_in_2_ chanx_right_in[6] chanx_left_in[6] mux_top_ipin_12.mux_l1_in_2_/S
+ mux_top_ipin_12.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l2_in_3__S mux_top_ipin_7.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l4_in_0__S mux_top_ipin_5.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_1__A1 mux_top_ipin_4.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_0.mux_l1_in_2_/S
+ mux_top_ipin_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_2.mux_l2_in_3__A1 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_1.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_4.mux_l3_in_0__A1 mux_top_ipin_4.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_prog_clk clkbuf_3_6_0_prog_clk/A clkbuf_3_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_31_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_13.mux_l2_in_1__S mux_top_ipin_13.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__41__A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__36__A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_12.mux_l2_in_0_ mux_top_ipin_12.mux_l1_in_1_/X mux_top_ipin_12.mux_l1_in_0_/X
+ mux_top_ipin_12.mux_l2_in_2_/S mux_top_ipin_12.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_12.mux_l3_in_1__S mux_top_ipin_12.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_5.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_5.mux_l1_in_0_/S
+ mux_top_ipin_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_15.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_12.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_12.mux_l1_in_2_/S
+ mux_top_ipin_12.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__44__A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_4.mux_l1_in_0__S mux_top_ipin_4.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__39__A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_1.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l2_in_1__A0 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_7.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_8.mux_l2_in_0__A0 mux_top_ipin_8.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_3.mux_l2_in_0__S mux_top_ipin_3.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_11.mux_l2_in_3__A0 _22_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__52__A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_13.mux_l3_in_0__A0 mux_top_ipin_13.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_3_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__47__A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_15.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_12.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_12.mux_l1_in_2_/S
+ mux_top_ipin_12.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_2.mux_l3_in_0__S mux_top_ipin_2.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l3_in_1__A0 mux_top_ipin_6.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_8.mux_l2_in_1__S mux_top_ipin_8.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_2.mux_l3_in_0_/S mux_top_ipin_2.mux_l4_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__60__A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_8.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_3.mux_l2_in_3__S mux_top_ipin_3.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_1.mux_l4_in_0__S mux_top_ipin_1.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_6.mux_l4_in_0__A0 mux_top_ipin_6.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_12.mux_l3_in_0_/S mux_top_ipin_12.mux_l4_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__55__A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_8.mux_l4_in_0_/X bottom_grid_pin_8_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l3_in_1__S mux_top_ipin_7.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_8.mux_l2_in_0__A1 mux_top_ipin_8.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_11.mux_l2_in_3__A1 chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_10.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_13.mux_l3_in_0__A1 mux_top_ipin_13.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_6.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_15.mux_l1_in_2__S mux_top_ipin_15.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_5.mux_l3_in_1_/S mux_top_ipin_5.mux_l4_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D ccff_head VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_9.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__63__A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_3_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_6_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__58__A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l3_in_1__A1 mux_top_ipin_6.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_15.mux_l3_in_1_/S ccff_tail
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_2.mux_l2_in_1_/S mux_top_ipin_2.mux_l3_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_14.mux_l2_in_2__S mux_top_ipin_14.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_1.mux_l2_in_3_ _20_/HI chanx_right_in[13] mux_top_ipin_1.mux_l2_in_3_/S
+ mux_top_ipin_1.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_3.mux_l2_in_0__A0 mux_top_ipin_3.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_6.mux_l4_in_0__A1 mux_top_ipin_6.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_12.mux_l2_in_2_/S mux_top_ipin_12.mux_l3_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__71__A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_10.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_0.mux_l1_in_0__S mux_top_ipin_0.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_2__A0 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_8.mux_l3_in_1_/S mux_top_ipin_8.mux_l4_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__66__A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_1.mux_l4_in_0_ mux_top_ipin_1.mux_l3_in_1_/X mux_top_ipin_1.mux_l3_in_0_/X
+ mux_top_ipin_1.mux_l4_in_0_/S mux_top_ipin_1.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_10.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_5_0_prog_clk clkbuf_2_2_0_prog_clk/X clkbuf_3_5_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_15.mux_l4_in_0_/X bottom_grid_pin_15_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_18_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l3_in_1__A0 mux_top_ipin_1.mux_l2_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_69_ chanx_left_in[5] chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_5.mux_l2_in_3_/S mux_top_ipin_5.mux_l3_in_1_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_30_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_6.mux_l2_in_3_ _31_/HI chanx_right_in[18] mux_top_ipin_6.mux_l2_in_3_/S
+ mux_top_ipin_6.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_1.mux_l3_in_1_ mux_top_ipin_1.mux_l2_in_3_/X mux_top_ipin_1.mux_l2_in_2_/X
+ mux_top_ipin_1.mux_l3_in_1_/S mux_top_ipin_1.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_15.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__74__A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_15.mux_l2_in_3_/S mux_top_ipin_15.mux_l3_in_1_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_1.mux_l4_in_0__A0 mux_top_ipin_1.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_15.mux_l2_in_2__A0 chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_2.mux_l1_in_0_/S mux_top_ipin_2.mux_l2_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__CLK clkbuf_3_2_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__69__A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_1.mux_l2_in_2_ chanx_left_in[13] chanx_right_in[5] mux_top_ipin_1.mux_l2_in_3_/S
+ mux_top_ipin_1.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_6.mux_l4_in_0_ mux_top_ipin_6.mux_l3_in_1_/X mux_top_ipin_6.mux_l3_in_0_/X
+ mux_top_ipin_6.mux_l4_in_0_/S mux_top_ipin_6.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_4.mux_l2_in_1__S mux_top_ipin_4.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0__A1 mux_top_ipin_3.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_12.mux_l1_in_2_/S mux_top_ipin_12.mux_l2_in_2_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_15.mux_l3_in_1__A0 mux_top_ipin_15.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_8.mux_l2_in_3__A0 _17_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_1.mux_l2_in_2__A1 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_8.mux_l2_in_0_/S mux_top_ipin_8.mux_l3_in_1_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_6.mux_l3_in_1_ mux_top_ipin_6.mux_l2_in_3_/X mux_top_ipin_6.mux_l2_in_2_/X
+ mux_top_ipin_6.mux_l3_in_1_/S mux_top_ipin_6.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_15.mux_l4_in_0__A0 mux_top_ipin_15.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_3_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l3_in_1__S mux_top_ipin_3.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_2_0_prog_clk_A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_1.mux_l4_in_0_/X bottom_grid_pin_1_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_ipin_9.mux_l2_in_2__S mux_top_ipin_9.mux_l2_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_68_ chanx_left_in[6] chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_1.mux_l3_in_1__A1 mux_top_ipin_1.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_5.mux_l1_in_0_/S mux_top_ipin_5.mux_l2_in_3_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_6.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[10] mux_top_ipin_6.mux_l2_in_3_/S
+ mux_top_ipin_6.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_1.mux_l3_in_0_ mux_top_ipin_1.mux_l2_in_1_/X mux_top_ipin_1.mux_l2_in_0_/X
+ mux_top_ipin_1.mux_l3_in_1_/S mux_top_ipin_1.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_11.mux_l1_in_2__S mux_top_ipin_11.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_13.mux_l2_in_3_ _24_/HI chanx_right_in[17] mux_top_ipin_13.mux_l2_in_3_/S
+ mux_top_ipin_13.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_15.mux_l1_in_1_/S mux_top_ipin_15.mux_l2_in_3_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_1.mux_l4_in_0__A1 mux_top_ipin_1.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_15.mux_l2_in_2__A1 chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_1.mux_l4_in_0_/S mux_top_ipin_2.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_15.mux_l2_in_0__S mux_top_ipin_15.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_1.mux_l2_in_1_ chanx_left_in[5] chanx_right_in[3] mux_top_ipin_1.mux_l2_in_3_/S
+ mux_top_ipin_1.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_11.mux_l4_in_0_/S mux_top_ipin_12.mux_l1_in_2_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_12.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l2_in_2__S mux_top_ipin_10.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_7_0_prog_clk_A clkbuf_3_6_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_15.mux_l3_in_1__A1 mux_top_ipin_15.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_8.mux_l2_in_3__A1 chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_13.mux_l4_in_0_ mux_top_ipin_13.mux_l3_in_1_/X mux_top_ipin_13.mux_l3_in_0_/X
+ mux_top_ipin_13.mux_l4_in_0_/S mux_top_ipin_13.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_14.mux_l3_in_0__S mux_top_ipin_14.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_7.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_8.mux_l1_in_1_/S mux_top_ipin_8.mux_l2_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_26_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_6.mux_l3_in_0_ mux_top_ipin_6.mux_l2_in_1_/X mux_top_ipin_6.mux_l2_in_0_/X
+ mux_top_ipin_6.mux_l3_in_1_/S mux_top_ipin_6.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_12.mux_l2_in_0__A0 mux_top_ipin_12.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_15.mux_l4_in_0__A1 mux_top_ipin_15.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_ipin_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_13.mux_l3_in_1_ mux_top_ipin_13.mux_l2_in_3_/X mux_top_ipin_13.mux_l2_in_2_/X
+ mux_top_ipin_13.mux_l3_in_1_/S mux_top_ipin_13.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_67_ chanx_left_in[7] chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_15.mux_l2_in_3__S mux_top_ipin_15.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l4_in_0__S mux_top_ipin_13.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_4.mux_l4_in_0_/S mux_top_ipin_5.mux_l1_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_10.mux_l2_in_2__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_6.mux_l2_in_1_ chanx_left_in[10] chanx_right_in[2] mux_top_ipin_6.mux_l2_in_3_/S
+ mux_top_ipin_6.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_ipin_5.mux_l2_in_1__A0 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_13.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[9] mux_top_ipin_13.mux_l2_in_3_/S
+ mux_top_ipin_13.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_14.mux_l4_in_0_/S mux_top_ipin_15.mux_l1_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_10.mux_l3_in_1__A0 mux_top_ipin_10.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_3__A0 _28_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_6.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_2_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_1.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_1.mux_l1_in_0_/X mux_top_ipin_1.mux_l2_in_3_/S
+ mux_top_ipin_1.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_5.mux_l3_in_0__A0 mux_top_ipin_5.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_12.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_3_7_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l4_in_0__A0 mux_top_ipin_10.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

