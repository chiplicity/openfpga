magic
tech sky130A
magscale 1 2
timestamp 1606477556
<< locali >>
rect 18153 19839 18187 20009
rect 16129 19159 16163 19261
rect 12909 18683 12943 18853
rect 15761 18615 15795 18853
rect 4905 18207 4939 18377
rect 15577 18071 15611 18241
rect 10333 16983 10367 17153
rect 15301 17051 15335 17289
rect 15025 16643 15059 16745
rect 6653 16031 6687 16201
rect 9045 15895 9079 16133
rect 12633 15419 12667 15589
rect 3249 14875 3283 15045
rect 10241 14875 10275 15045
rect 18797 14943 18831 15113
rect 13185 14263 13219 14569
rect 15025 13175 15059 13277
rect 17325 13175 17359 13413
rect 16405 12223 16439 12393
rect 19809 12155 19843 12325
rect 16313 11747 16347 11849
rect 19533 11543 19567 11781
rect 19073 11135 19107 11305
rect 7573 10455 7607 10761
rect 9505 9911 9539 10081
rect 12449 8823 12483 8925
rect 15117 8823 15151 8993
rect 16129 8891 16163 9061
rect 9413 8347 9447 8449
rect 12265 8415 12299 8585
rect 2145 7939 2179 8041
rect 4905 7871 4939 7973
rect 9413 7735 9447 8041
rect 12115 7905 12207 7939
rect 12173 7735 12207 7905
rect 16865 7803 16899 7905
rect 9689 7259 9723 7429
rect 9781 6783 9815 6953
rect 11805 6851 11839 6953
rect 19073 6783 19107 6885
rect 3341 6647 3375 6749
rect 4997 6171 5031 6341
rect 15669 5083 15703 5253
rect 17785 5219 17819 5321
rect 13369 4471 13403 4709
rect 17325 4607 17359 4709
rect 18245 4471 18279 4777
rect 12449 4063 12483 4165
rect 14657 4131 14691 4233
rect 13001 3927 13035 4097
rect 17049 3519 17083 3689
rect 14013 2907 14047 3145
rect 18153 3043 18187 3145
rect 10701 2295 10735 2533
rect 11161 1683 11195 1785
rect 8769 1411 8803 1581
<< viali >>
rect 4077 20009 4111 20043
rect 10241 20009 10275 20043
rect 15025 20009 15059 20043
rect 18153 20009 18187 20043
rect 3525 19941 3559 19975
rect 6377 19941 6411 19975
rect 8953 19941 8987 19975
rect 11069 19941 11103 19975
rect 11897 19941 11931 19975
rect 14105 19941 14139 19975
rect 17049 19941 17083 19975
rect 1685 19873 1719 19907
rect 2421 19873 2455 19907
rect 3249 19873 3283 19907
rect 4445 19873 4479 19907
rect 5457 19873 5491 19907
rect 6101 19873 6135 19907
rect 7196 19873 7230 19907
rect 10149 19873 10183 19907
rect 10793 19873 10827 19907
rect 12633 19873 12667 19907
rect 14841 19873 14875 19907
rect 15853 19873 15887 19907
rect 16773 19873 16807 19907
rect 17509 19873 17543 19907
rect 19901 19941 19935 19975
rect 20637 19941 20671 19975
rect 18337 19873 18371 19907
rect 18889 19873 18923 19907
rect 19625 19873 19659 19907
rect 20361 19873 20395 19907
rect 1869 19805 1903 19839
rect 2697 19805 2731 19839
rect 4537 19805 4571 19839
rect 4721 19805 4755 19839
rect 5549 19805 5583 19839
rect 5733 19805 5767 19839
rect 6929 19805 6963 19839
rect 9045 19805 9079 19839
rect 9137 19805 9171 19839
rect 10425 19805 10459 19839
rect 11989 19805 12023 19839
rect 12081 19805 12115 19839
rect 12909 19805 12943 19839
rect 14197 19805 14231 19839
rect 14381 19805 14415 19839
rect 15945 19805 15979 19839
rect 16129 19805 16163 19839
rect 17785 19805 17819 19839
rect 18153 19805 18187 19839
rect 19165 19805 19199 19839
rect 13737 19737 13771 19771
rect 5089 19669 5123 19703
rect 8309 19669 8343 19703
rect 8585 19669 8619 19703
rect 9781 19669 9815 19703
rect 11529 19669 11563 19703
rect 15485 19669 15519 19703
rect 18521 19669 18555 19703
rect 8401 19465 8435 19499
rect 12449 19465 12483 19499
rect 3341 19397 3375 19431
rect 3801 19397 3835 19431
rect 10241 19397 10275 19431
rect 4445 19329 4479 19363
rect 11989 19329 12023 19363
rect 13093 19329 13127 19363
rect 16865 19329 16899 19363
rect 20729 19329 20763 19363
rect 1685 19261 1719 19295
rect 1961 19261 1995 19295
rect 2421 19261 2455 19295
rect 2697 19261 2731 19295
rect 3157 19261 3191 19295
rect 4169 19261 4203 19295
rect 4813 19261 4847 19295
rect 5080 19261 5114 19295
rect 7021 19261 7055 19295
rect 8861 19261 8895 19295
rect 10517 19261 10551 19295
rect 11805 19261 11839 19295
rect 13461 19261 13495 19295
rect 14370 19261 14404 19295
rect 15117 19261 15151 19295
rect 15669 19261 15703 19295
rect 16129 19261 16163 19295
rect 17233 19261 17267 19295
rect 17509 19261 17543 19295
rect 18061 19261 18095 19295
rect 18797 19261 18831 19295
rect 7288 19193 7322 19227
rect 9128 19193 9162 19227
rect 10793 19193 10827 19227
rect 12817 19193 12851 19227
rect 14657 19193 14691 19227
rect 19441 19193 19475 19227
rect 20637 19193 20671 19227
rect 4261 19125 4295 19159
rect 6193 19125 6227 19159
rect 11345 19125 11379 19159
rect 11713 19125 11747 19159
rect 12909 19125 12943 19159
rect 13645 19125 13679 19159
rect 15301 19125 15335 19159
rect 15853 19125 15887 19159
rect 16129 19125 16163 19159
rect 16221 19125 16255 19159
rect 16589 19125 16623 19159
rect 16681 19125 16715 19159
rect 18245 19125 18279 19159
rect 20177 19125 20211 19159
rect 20545 19125 20579 19159
rect 2329 18921 2363 18955
rect 2973 18921 3007 18955
rect 3341 18921 3375 18955
rect 6193 18921 6227 18955
rect 6929 18921 6963 18955
rect 9689 18921 9723 18955
rect 10057 18921 10091 18955
rect 17693 18921 17727 18955
rect 19257 18921 19291 18955
rect 19809 18921 19843 18955
rect 12909 18853 12943 18887
rect 13338 18853 13372 18887
rect 15761 18853 15795 18887
rect 18337 18853 18371 18887
rect 20177 18853 20211 18887
rect 1409 18785 1443 18819
rect 4077 18785 4111 18819
rect 4344 18785 4378 18819
rect 6101 18785 6135 18819
rect 6745 18785 6779 18819
rect 7389 18785 7423 18819
rect 7656 18785 7690 18819
rect 9045 18785 9079 18819
rect 10149 18785 10183 18819
rect 10701 18785 10735 18819
rect 11704 18785 11738 18819
rect 2421 18717 2455 18751
rect 2605 18717 2639 18751
rect 3433 18717 3467 18751
rect 3617 18717 3651 18751
rect 6285 18717 6319 18751
rect 10241 18717 10275 18751
rect 10977 18717 11011 18751
rect 11437 18717 11471 18751
rect 15301 18785 15335 18819
rect 13093 18717 13127 18751
rect 12817 18649 12851 18683
rect 12909 18649 12943 18683
rect 16120 18785 16154 18819
rect 17509 18785 17543 18819
rect 18061 18785 18095 18819
rect 19165 18785 19199 18819
rect 15853 18717 15887 18751
rect 19349 18717 19383 18751
rect 20269 18717 20303 18751
rect 20453 18717 20487 18751
rect 1593 18581 1627 18615
rect 1961 18581 1995 18615
rect 5457 18581 5491 18615
rect 5733 18581 5767 18615
rect 8769 18581 8803 18615
rect 9229 18581 9263 18615
rect 14473 18581 14507 18615
rect 15485 18581 15519 18615
rect 15761 18581 15795 18615
rect 17233 18581 17267 18615
rect 18797 18581 18831 18615
rect 1961 18377 1995 18411
rect 4905 18377 4939 18411
rect 7481 18377 7515 18411
rect 8493 18377 8527 18411
rect 9505 18377 9539 18411
rect 12081 18377 12115 18411
rect 12449 18377 12483 18411
rect 15761 18377 15795 18411
rect 20269 18377 20303 18411
rect 4721 18241 4755 18275
rect 7113 18309 7147 18343
rect 13461 18309 13495 18343
rect 17049 18309 17083 18343
rect 7941 18241 7975 18275
rect 8125 18241 8159 18275
rect 9045 18241 9079 18275
rect 10057 18241 10091 18275
rect 12909 18241 12943 18275
rect 13093 18241 13127 18275
rect 14105 18241 14139 18275
rect 15209 18241 15243 18275
rect 15301 18241 15335 18275
rect 15577 18241 15611 18275
rect 16313 18241 16347 18275
rect 17509 18241 17543 18275
rect 19073 18241 19107 18275
rect 19717 18241 19751 18275
rect 20821 18241 20855 18275
rect 1777 18173 1811 18207
rect 2421 18173 2455 18207
rect 4445 18173 4479 18207
rect 4537 18173 4571 18207
rect 4905 18173 4939 18207
rect 5089 18173 5123 18207
rect 6929 18173 6963 18207
rect 7849 18173 7883 18207
rect 8953 18173 8987 18207
rect 9965 18173 9999 18207
rect 10701 18173 10735 18207
rect 13921 18173 13955 18207
rect 15117 18173 15151 18207
rect 2688 18105 2722 18139
rect 5356 18105 5390 18139
rect 10968 18105 11002 18139
rect 13829 18105 13863 18139
rect 16129 18173 16163 18207
rect 16865 18173 16899 18207
rect 17233 18173 17267 18207
rect 18061 18173 18095 18207
rect 19533 18173 19567 18207
rect 18889 18105 18923 18139
rect 20729 18105 20763 18139
rect 3801 18037 3835 18071
rect 4077 18037 4111 18071
rect 6469 18037 6503 18071
rect 8861 18037 8895 18071
rect 9873 18037 9907 18071
rect 12817 18037 12851 18071
rect 14749 18037 14783 18071
rect 15577 18037 15611 18071
rect 16221 18037 16255 18071
rect 18245 18037 18279 18071
rect 18429 18037 18463 18071
rect 18797 18037 18831 18071
rect 20637 18037 20671 18071
rect 1777 17833 1811 17867
rect 2421 17833 2455 17867
rect 2881 17833 2915 17867
rect 4077 17833 4111 17867
rect 4537 17833 4571 17867
rect 5089 17833 5123 17867
rect 7297 17833 7331 17867
rect 8585 17833 8619 17867
rect 11345 17833 11379 17867
rect 13001 17833 13035 17867
rect 14657 17833 14691 17867
rect 15301 17833 15335 17867
rect 15761 17833 15795 17867
rect 16313 17833 16347 17867
rect 17785 17833 17819 17867
rect 18521 17833 18555 17867
rect 1869 17765 1903 17799
rect 4445 17765 4479 17799
rect 7665 17765 7699 17799
rect 10425 17765 10459 17799
rect 12081 17765 12115 17799
rect 13737 17765 13771 17799
rect 17693 17765 17727 17799
rect 19901 17765 19935 17799
rect 2789 17697 2823 17731
rect 3433 17697 3467 17731
rect 5457 17697 5491 17731
rect 6653 17697 6687 17731
rect 6745 17697 6779 17731
rect 8953 17697 8987 17731
rect 9045 17697 9079 17731
rect 10333 17697 10367 17731
rect 11161 17697 11195 17731
rect 12817 17697 12851 17731
rect 13461 17697 13495 17731
rect 14565 17697 14599 17731
rect 15669 17697 15703 17731
rect 16681 17697 16715 17731
rect 16773 17697 16807 17731
rect 18889 17697 18923 17731
rect 19993 17697 20027 17731
rect 2053 17629 2087 17663
rect 2973 17629 3007 17663
rect 4721 17629 4755 17663
rect 5549 17629 5583 17663
rect 5641 17629 5675 17663
rect 6929 17629 6963 17663
rect 7757 17629 7791 17663
rect 7941 17629 7975 17663
rect 9137 17629 9171 17663
rect 10609 17629 10643 17663
rect 12173 17629 12207 17663
rect 12265 17629 12299 17663
rect 14841 17629 14875 17663
rect 15853 17629 15887 17663
rect 16865 17629 16899 17663
rect 17877 17629 17911 17663
rect 18981 17629 19015 17663
rect 19073 17629 19107 17663
rect 20177 17629 20211 17663
rect 1409 17561 1443 17595
rect 3617 17561 3651 17595
rect 6285 17493 6319 17527
rect 9965 17493 9999 17527
rect 11713 17493 11747 17527
rect 14197 17493 14231 17527
rect 17325 17493 17359 17527
rect 18337 17493 18371 17527
rect 19533 17493 19567 17527
rect 3525 17289 3559 17323
rect 5181 17289 5215 17323
rect 8401 17289 8435 17323
rect 12449 17289 12483 17323
rect 15117 17289 15151 17323
rect 15301 17289 15335 17323
rect 18061 17289 18095 17323
rect 4077 17221 4111 17255
rect 8033 17221 8067 17255
rect 11989 17221 12023 17255
rect 4721 17153 4755 17187
rect 5825 17153 5859 17187
rect 6285 17153 6319 17187
rect 7389 17153 7423 17187
rect 9045 17153 9079 17187
rect 9965 17153 9999 17187
rect 10333 17153 10367 17187
rect 10977 17153 11011 17187
rect 12909 17153 12943 17187
rect 13093 17153 13127 17187
rect 1409 17085 1443 17119
rect 2145 17085 2179 17119
rect 2412 17085 2446 17119
rect 7297 17085 7331 17119
rect 7849 17085 7883 17119
rect 1685 17017 1719 17051
rect 4445 17017 4479 17051
rect 4537 17017 4571 17051
rect 7205 17017 7239 17051
rect 8769 17017 8803 17051
rect 9873 17017 9907 17051
rect 11805 17085 11839 17119
rect 13737 17085 13771 17119
rect 17141 17221 17175 17255
rect 15393 17153 15427 17187
rect 17693 17153 17727 17187
rect 18705 17153 18739 17187
rect 19717 17153 19751 17187
rect 20729 17153 20763 17187
rect 19441 17085 19475 17119
rect 10885 17017 10919 17051
rect 14004 17017 14038 17051
rect 15301 17017 15335 17051
rect 15638 17017 15672 17051
rect 18521 17017 18555 17051
rect 19533 17017 19567 17051
rect 20453 17017 20487 17051
rect 5273 16949 5307 16983
rect 5641 16949 5675 16983
rect 5733 16949 5767 16983
rect 6837 16949 6871 16983
rect 8861 16949 8895 16983
rect 9413 16949 9447 16983
rect 9781 16949 9815 16983
rect 10333 16949 10367 16983
rect 10425 16949 10459 16983
rect 10793 16949 10827 16983
rect 12817 16949 12851 16983
rect 16773 16949 16807 16983
rect 17509 16949 17543 16983
rect 17601 16949 17635 16983
rect 18429 16949 18463 16983
rect 19073 16949 19107 16983
rect 20085 16949 20119 16983
rect 20545 16949 20579 16983
rect 1961 16745 1995 16779
rect 2973 16745 3007 16779
rect 4537 16745 4571 16779
rect 7389 16745 7423 16779
rect 9321 16745 9355 16779
rect 10149 16745 10183 16779
rect 11897 16745 11931 16779
rect 14381 16745 14415 16779
rect 14841 16745 14875 16779
rect 15025 16745 15059 16779
rect 15577 16745 15611 16779
rect 15945 16745 15979 16779
rect 16037 16745 16071 16779
rect 16589 16745 16623 16779
rect 16957 16745 16991 16779
rect 17601 16745 17635 16779
rect 18981 16745 19015 16779
rect 19993 16745 20027 16779
rect 1869 16677 1903 16711
rect 2329 16677 2363 16711
rect 2421 16677 2455 16711
rect 8208 16677 8242 16711
rect 13268 16677 13302 16711
rect 18061 16677 18095 16711
rect 20085 16677 20119 16711
rect 3341 16609 3375 16643
rect 3433 16609 3467 16643
rect 4445 16609 4479 16643
rect 5540 16609 5574 16643
rect 7297 16609 7331 16643
rect 9965 16609 9999 16643
rect 10784 16609 10818 16643
rect 12265 16609 12299 16643
rect 12541 16609 12575 16643
rect 14657 16609 14691 16643
rect 15025 16609 15059 16643
rect 17969 16609 18003 16643
rect 19073 16609 19107 16643
rect 20913 16609 20947 16643
rect 2605 16541 2639 16575
rect 3525 16541 3559 16575
rect 4629 16541 4663 16575
rect 5273 16541 5307 16575
rect 7481 16541 7515 16575
rect 7941 16541 7975 16575
rect 10517 16541 10551 16575
rect 13001 16541 13035 16575
rect 16221 16541 16255 16575
rect 17049 16541 17083 16575
rect 17233 16541 17267 16575
rect 18245 16541 18279 16575
rect 19165 16541 19199 16575
rect 20177 16541 20211 16575
rect 6929 16473 6963 16507
rect 18613 16473 18647 16507
rect 4077 16405 4111 16439
rect 4905 16405 4939 16439
rect 6653 16405 6687 16439
rect 19625 16405 19659 16439
rect 1593 16201 1627 16235
rect 2605 16201 2639 16235
rect 3801 16201 3835 16235
rect 6653 16201 6687 16235
rect 12449 16201 12483 16235
rect 13461 16201 13495 16235
rect 15853 16201 15887 16235
rect 18245 16201 18279 16235
rect 3157 16065 3191 16099
rect 4261 16065 4295 16099
rect 4445 16065 4479 16099
rect 4813 16065 4847 16099
rect 5825 16065 5859 16099
rect 9045 16133 9079 16167
rect 9413 16133 9447 16167
rect 14841 16133 14875 16167
rect 16865 16133 16899 16167
rect 1409 15997 1443 16031
rect 1869 15997 1903 16031
rect 2145 15997 2179 16031
rect 3065 15997 3099 16031
rect 4169 15997 4203 16031
rect 6653 15997 6687 16031
rect 6837 15997 6871 16031
rect 8677 15997 8711 16031
rect 5733 15929 5767 15963
rect 7104 15929 7138 15963
rect 9965 16065 9999 16099
rect 13093 16065 13127 16099
rect 14013 16065 14047 16099
rect 15301 16065 15335 16099
rect 15485 16065 15519 16099
rect 16405 16065 16439 16099
rect 17417 16065 17451 16099
rect 18705 16065 18739 16099
rect 18797 16065 18831 16099
rect 19717 16065 19751 16099
rect 20637 16065 20671 16099
rect 10425 15997 10459 16031
rect 13921 15997 13955 16031
rect 15209 15997 15243 16031
rect 16313 15997 16347 16031
rect 9321 15929 9355 15963
rect 9873 15929 9907 15963
rect 10692 15929 10726 15963
rect 12817 15929 12851 15963
rect 17233 15929 17267 15963
rect 20453 15929 20487 15963
rect 2973 15861 3007 15895
rect 5273 15861 5307 15895
rect 5641 15861 5675 15895
rect 6285 15861 6319 15895
rect 8217 15861 8251 15895
rect 8861 15861 8895 15895
rect 9045 15861 9079 15895
rect 9781 15861 9815 15895
rect 11805 15861 11839 15895
rect 12909 15861 12943 15895
rect 13829 15861 13863 15895
rect 16221 15861 16255 15895
rect 17325 15861 17359 15895
rect 18613 15861 18647 15895
rect 19073 15861 19107 15895
rect 19441 15861 19475 15895
rect 19533 15861 19567 15895
rect 20085 15861 20119 15895
rect 20545 15861 20579 15895
rect 2329 15657 2363 15691
rect 8953 15657 8987 15691
rect 9689 15657 9723 15691
rect 10701 15657 10735 15691
rect 16405 15657 16439 15691
rect 18705 15657 18739 15691
rect 19441 15657 19475 15691
rect 19901 15657 19935 15691
rect 3433 15589 3467 15623
rect 4905 15589 4939 15623
rect 12633 15589 12667 15623
rect 13084 15589 13118 15623
rect 17785 15589 17819 15623
rect 1409 15521 1443 15555
rect 3341 15521 3375 15555
rect 4997 15521 5031 15555
rect 5917 15521 5951 15555
rect 6745 15521 6779 15555
rect 7196 15521 7230 15555
rect 9045 15521 9079 15555
rect 10057 15521 10091 15555
rect 11161 15521 11195 15555
rect 11428 15521 11462 15555
rect 2421 15453 2455 15487
rect 2513 15453 2547 15487
rect 3525 15453 3559 15487
rect 4077 15453 4111 15487
rect 5181 15453 5215 15487
rect 6009 15453 6043 15487
rect 6193 15453 6227 15487
rect 6929 15453 6963 15487
rect 9137 15453 9171 15487
rect 10149 15453 10183 15487
rect 10241 15453 10275 15487
rect 12817 15521 12851 15555
rect 14473 15521 14507 15555
rect 15669 15521 15703 15555
rect 16129 15521 16163 15555
rect 16773 15521 16807 15555
rect 17877 15521 17911 15555
rect 18613 15521 18647 15555
rect 19809 15521 19843 15555
rect 14657 15453 14691 15487
rect 15761 15453 15795 15487
rect 15853 15453 15887 15487
rect 16865 15453 16899 15487
rect 17049 15453 17083 15487
rect 17969 15453 18003 15487
rect 18889 15453 18923 15487
rect 19993 15453 20027 15487
rect 8309 15385 8343 15419
rect 8585 15385 8619 15419
rect 12541 15385 12575 15419
rect 12633 15385 12667 15419
rect 15301 15385 15335 15419
rect 1593 15317 1627 15351
rect 1961 15317 1995 15351
rect 2973 15317 3007 15351
rect 4537 15317 4571 15351
rect 5549 15317 5583 15351
rect 6561 15317 6595 15351
rect 14197 15317 14231 15351
rect 17417 15317 17451 15351
rect 18245 15317 18279 15351
rect 6837 15113 6871 15147
rect 11713 15113 11747 15147
rect 12449 15113 12483 15147
rect 18797 15113 18831 15147
rect 3065 15045 3099 15079
rect 3249 15045 3283 15079
rect 8033 15045 8067 15079
rect 8401 15045 8435 15079
rect 10057 15045 10091 15079
rect 10241 15045 10275 15079
rect 1685 14909 1719 14943
rect 7481 14977 7515 15011
rect 8677 14977 8711 15011
rect 3341 14909 3375 14943
rect 4997 14909 5031 14943
rect 7849 14909 7883 14943
rect 8585 14909 8619 14943
rect 13001 14977 13035 15011
rect 14105 14977 14139 15011
rect 16221 14977 16255 15011
rect 20085 15045 20119 15079
rect 19533 14977 19567 15011
rect 19717 14977 19751 15011
rect 20545 14977 20579 15011
rect 20729 14977 20763 15011
rect 10333 14909 10367 14943
rect 12265 14909 12299 14943
rect 12817 14909 12851 14943
rect 13553 14909 13587 14943
rect 18797 14909 18831 14943
rect 18889 14909 18923 14943
rect 19441 14909 19475 14943
rect 1952 14841 1986 14875
rect 3249 14841 3283 14875
rect 3586 14841 3620 14875
rect 5264 14841 5298 14875
rect 8944 14841 8978 14875
rect 10241 14841 10275 14875
rect 10578 14841 10612 14875
rect 14372 14841 14406 14875
rect 16488 14841 16522 14875
rect 4721 14773 4755 14807
rect 6377 14773 6411 14807
rect 7205 14773 7239 14807
rect 7297 14773 7331 14807
rect 12081 14773 12115 14807
rect 12909 14773 12943 14807
rect 13737 14773 13771 14807
rect 15485 14773 15519 14807
rect 15761 14773 15795 14807
rect 17601 14773 17635 14807
rect 19073 14773 19107 14807
rect 20453 14773 20487 14807
rect 3341 14569 3375 14603
rect 4261 14569 4295 14603
rect 4629 14569 4663 14603
rect 7573 14569 7607 14603
rect 8585 14569 8619 14603
rect 9873 14569 9907 14603
rect 10333 14569 10367 14603
rect 12817 14569 12851 14603
rect 13185 14569 13219 14603
rect 13737 14569 13771 14603
rect 16037 14569 16071 14603
rect 18981 14569 19015 14603
rect 19625 14569 19659 14603
rect 20085 14569 20119 14603
rect 20913 14569 20947 14603
rect 6162 14501 6196 14535
rect 8953 14501 8987 14535
rect 11713 14501 11747 14535
rect 12725 14501 12759 14535
rect 1409 14433 1443 14467
rect 2237 14433 2271 14467
rect 3249 14433 3283 14467
rect 4721 14433 4755 14467
rect 5273 14433 5307 14467
rect 5917 14433 5951 14467
rect 7941 14433 7975 14467
rect 9689 14433 9723 14467
rect 10701 14433 10735 14467
rect 2329 14365 2363 14399
rect 2513 14365 2547 14399
rect 3525 14365 3559 14399
rect 4813 14365 4847 14399
rect 8033 14365 8067 14399
rect 8125 14365 8159 14399
rect 9045 14365 9079 14399
rect 9137 14365 9171 14399
rect 10793 14365 10827 14399
rect 10885 14365 10919 14399
rect 11805 14365 11839 14399
rect 11897 14365 11931 14399
rect 13001 14365 13035 14399
rect 12357 14297 12391 14331
rect 20177 14501 20211 14535
rect 13829 14433 13863 14467
rect 14473 14433 14507 14467
rect 15301 14433 15335 14467
rect 16405 14433 16439 14467
rect 17049 14433 17083 14467
rect 17316 14433 17350 14467
rect 18889 14433 18923 14467
rect 13921 14365 13955 14399
rect 14749 14365 14783 14399
rect 15577 14365 15611 14399
rect 16497 14365 16531 14399
rect 16681 14365 16715 14399
rect 19073 14365 19107 14399
rect 20361 14365 20395 14399
rect 13369 14297 13403 14331
rect 18429 14297 18463 14331
rect 1869 14229 1903 14263
rect 2881 14229 2915 14263
rect 5457 14229 5491 14263
rect 7297 14229 7331 14263
rect 11345 14229 11379 14263
rect 13185 14229 13219 14263
rect 18521 14229 18555 14263
rect 19717 14229 19751 14263
rect 1869 14025 1903 14059
rect 5733 14025 5767 14059
rect 9137 14025 9171 14059
rect 9965 14025 9999 14059
rect 14749 14025 14783 14059
rect 16773 14025 16807 14059
rect 20913 14025 20947 14059
rect 2881 13957 2915 13991
rect 9597 13957 9631 13991
rect 14197 13957 14231 13991
rect 16497 13957 16531 13991
rect 19717 13957 19751 13991
rect 2513 13889 2547 13923
rect 3525 13889 3559 13923
rect 6285 13889 6319 13923
rect 7021 13889 7055 13923
rect 10517 13889 10551 13923
rect 11529 13889 11563 13923
rect 17417 13889 17451 13923
rect 20269 13889 20303 13923
rect 3893 13821 3927 13855
rect 4149 13821 4183 13855
rect 6193 13821 6227 13855
rect 6837 13821 6871 13855
rect 7757 13821 7791 13855
rect 8024 13821 8058 13855
rect 9413 13821 9447 13855
rect 12817 13821 12851 13855
rect 13084 13821 13118 13855
rect 14565 13821 14599 13855
rect 15117 13821 15151 13855
rect 18061 13821 18095 13855
rect 18317 13821 18351 13855
rect 20177 13821 20211 13855
rect 20729 13821 20763 13855
rect 3341 13753 3375 13787
rect 11345 13753 11379 13787
rect 15362 13753 15396 13787
rect 17233 13753 17267 13787
rect 1409 13685 1443 13719
rect 2237 13685 2271 13719
rect 2329 13685 2363 13719
rect 3249 13685 3283 13719
rect 5273 13685 5307 13719
rect 6101 13685 6135 13719
rect 10333 13685 10367 13719
rect 10425 13685 10459 13719
rect 10977 13685 11011 13719
rect 11437 13685 11471 13719
rect 17141 13685 17175 13719
rect 19441 13685 19475 13719
rect 20085 13685 20119 13719
rect 4537 13481 4571 13515
rect 5181 13481 5215 13515
rect 6837 13481 6871 13515
rect 11253 13481 11287 13515
rect 11621 13481 11655 13515
rect 12541 13481 12575 13515
rect 15301 13481 15335 13515
rect 15761 13481 15795 13515
rect 16405 13481 16439 13515
rect 17785 13481 17819 13515
rect 19441 13481 19475 13515
rect 19809 13481 19843 13515
rect 1869 13413 1903 13447
rect 5549 13413 5583 13447
rect 8309 13413 8343 13447
rect 10149 13413 10183 13447
rect 12909 13413 12943 13447
rect 17325 13413 17359 13447
rect 19901 13413 19935 13447
rect 1593 13345 1627 13379
rect 2329 13345 2363 13379
rect 2596 13345 2630 13379
rect 4629 13345 4663 13379
rect 6193 13345 6227 13379
rect 7205 13345 7239 13379
rect 8217 13345 8251 13379
rect 8861 13345 8895 13379
rect 10057 13345 10091 13379
rect 10701 13345 10735 13379
rect 13820 13345 13854 13379
rect 15669 13345 15703 13379
rect 16773 13345 16807 13379
rect 4721 13277 4755 13311
rect 5641 13277 5675 13311
rect 5733 13277 5767 13311
rect 7297 13277 7331 13311
rect 7481 13277 7515 13311
rect 8493 13277 8527 13311
rect 10241 13277 10275 13311
rect 11713 13277 11747 13311
rect 11897 13277 11931 13311
rect 13001 13277 13035 13311
rect 13185 13277 13219 13311
rect 13553 13277 13587 13311
rect 15025 13277 15059 13311
rect 15945 13277 15979 13311
rect 16865 13277 16899 13311
rect 16957 13277 16991 13311
rect 10885 13209 10919 13243
rect 3709 13141 3743 13175
rect 4169 13141 4203 13175
rect 6377 13141 6411 13175
rect 7849 13141 7883 13175
rect 9045 13141 9079 13175
rect 9689 13141 9723 13175
rect 14933 13141 14967 13175
rect 15025 13141 15059 13175
rect 17877 13345 17911 13379
rect 18797 13345 18831 13379
rect 17969 13277 18003 13311
rect 18889 13277 18923 13311
rect 19073 13277 19107 13311
rect 19993 13277 20027 13311
rect 17325 13141 17359 13175
rect 17417 13141 17451 13175
rect 18429 13141 18463 13175
rect 1593 12937 1627 12971
rect 5457 12937 5491 12971
rect 6469 12937 6503 12971
rect 7205 12937 7239 12971
rect 9965 12937 9999 12971
rect 10977 12937 11011 12971
rect 15761 12937 15795 12971
rect 16313 12937 16347 12971
rect 3985 12869 4019 12903
rect 8677 12869 8711 12903
rect 14105 12869 14139 12903
rect 14381 12869 14415 12903
rect 15301 12869 15335 12903
rect 2053 12801 2087 12835
rect 2237 12801 2271 12835
rect 4813 12801 4847 12835
rect 6009 12801 6043 12835
rect 9505 12801 9539 12835
rect 10517 12801 10551 12835
rect 11437 12801 11471 12835
rect 11621 12801 11655 12835
rect 11897 12801 11931 12835
rect 14979 12801 15013 12835
rect 16129 12801 16163 12835
rect 16957 12801 16991 12835
rect 19441 12801 19475 12835
rect 20453 12801 20487 12835
rect 2605 12733 2639 12767
rect 4721 12733 4755 12767
rect 6653 12733 6687 12767
rect 7297 12733 7331 12767
rect 9321 12733 9355 12767
rect 10333 12733 10367 12767
rect 10425 12733 10459 12767
rect 11345 12733 11379 12767
rect 12725 12733 12759 12767
rect 15485 12733 15519 12767
rect 15577 12733 15611 12767
rect 16681 12733 16715 12767
rect 17417 12733 17451 12767
rect 18153 12733 18187 12767
rect 19257 12733 19291 12767
rect 20361 12733 20395 12767
rect 2872 12665 2906 12699
rect 5825 12665 5859 12699
rect 6837 12665 6871 12699
rect 7542 12665 7576 12699
rect 12992 12665 13026 12699
rect 18429 12665 18463 12699
rect 20269 12665 20303 12699
rect 1961 12597 1995 12631
rect 4261 12597 4295 12631
rect 4629 12597 4663 12631
rect 5917 12597 5951 12631
rect 8953 12597 8987 12631
rect 9413 12597 9447 12631
rect 14749 12597 14783 12631
rect 14841 12597 14875 12631
rect 16773 12597 16807 12631
rect 17601 12597 17635 12631
rect 18889 12597 18923 12631
rect 19349 12597 19383 12631
rect 19901 12597 19935 12631
rect 1593 12393 1627 12427
rect 1961 12393 1995 12427
rect 2329 12393 2363 12427
rect 2973 12393 3007 12427
rect 4261 12393 4295 12427
rect 6101 12393 6135 12427
rect 6745 12393 6779 12427
rect 7389 12393 7423 12427
rect 8861 12393 8895 12427
rect 13093 12393 13127 12427
rect 14105 12393 14139 12427
rect 14473 12393 14507 12427
rect 16405 12393 16439 12427
rect 17877 12393 17911 12427
rect 2421 12325 2455 12359
rect 15853 12325 15887 12359
rect 1409 12257 1443 12291
rect 3341 12257 3375 12291
rect 4077 12257 4111 12291
rect 4977 12257 5011 12291
rect 6837 12257 6871 12291
rect 7757 12257 7791 12291
rect 8769 12257 8803 12291
rect 9781 12257 9815 12291
rect 10048 12257 10082 12291
rect 11704 12257 11738 12291
rect 13461 12257 13495 12291
rect 19809 12325 19843 12359
rect 20177 12325 20211 12359
rect 16764 12257 16798 12291
rect 18245 12257 18279 12291
rect 18512 12257 18546 12291
rect 2605 12189 2639 12223
rect 3433 12189 3467 12223
rect 3617 12189 3651 12223
rect 4721 12189 4755 12223
rect 6929 12189 6963 12223
rect 7849 12189 7883 12223
rect 7941 12189 7975 12223
rect 9045 12189 9079 12223
rect 11437 12189 11471 12223
rect 13553 12189 13587 12223
rect 13737 12189 13771 12223
rect 14565 12189 14599 12223
rect 14657 12189 14691 12223
rect 15945 12189 15979 12223
rect 16129 12189 16163 12223
rect 16405 12189 16439 12223
rect 16497 12189 16531 12223
rect 19901 12257 19935 12291
rect 20913 12189 20947 12223
rect 6377 12121 6411 12155
rect 11161 12121 11195 12155
rect 19809 12121 19843 12155
rect 8401 12053 8435 12087
rect 12817 12053 12851 12087
rect 15485 12053 15519 12087
rect 19625 12053 19659 12087
rect 5089 11849 5123 11883
rect 5549 11849 5583 11883
rect 6837 11849 6871 11883
rect 7849 11849 7883 11883
rect 9045 11849 9079 11883
rect 9873 11849 9907 11883
rect 15761 11849 15795 11883
rect 16037 11849 16071 11883
rect 16313 11849 16347 11883
rect 16589 11849 16623 11883
rect 19441 11849 19475 11883
rect 20913 11849 20947 11883
rect 2145 11781 2179 11815
rect 4629 11781 4663 11815
rect 11529 11781 11563 11815
rect 13829 11781 13863 11815
rect 14105 11781 14139 11815
rect 19533 11781 19567 11815
rect 19717 11781 19751 11815
rect 2789 11713 2823 11747
rect 6101 11713 6135 11747
rect 7389 11713 7423 11747
rect 8309 11713 8343 11747
rect 8401 11713 8435 11747
rect 9597 11713 9631 11747
rect 10517 11713 10551 11747
rect 11253 11713 11287 11747
rect 12173 11713 12207 11747
rect 12449 11713 12483 11747
rect 16313 11713 16347 11747
rect 17417 11713 17451 11747
rect 17601 11713 17635 11747
rect 1409 11645 1443 11679
rect 3249 11645 3283 11679
rect 3505 11645 3539 11679
rect 4905 11645 4939 11679
rect 5917 11645 5951 11679
rect 7205 11645 7239 11679
rect 8217 11645 8251 11679
rect 10333 11645 10367 11679
rect 11069 11645 11103 11679
rect 12716 11645 12750 11679
rect 14289 11645 14323 11679
rect 14381 11645 14415 11679
rect 16221 11645 16255 11679
rect 16405 11645 16439 11679
rect 18061 11645 18095 11679
rect 18328 11645 18362 11679
rect 1685 11577 1719 11611
rect 9413 11577 9447 11611
rect 9505 11577 9539 11611
rect 14637 11577 14671 11611
rect 20269 11713 20303 11747
rect 20085 11645 20119 11679
rect 20729 11645 20763 11679
rect 20177 11577 20211 11611
rect 2513 11509 2547 11543
rect 2605 11509 2639 11543
rect 6009 11509 6043 11543
rect 7297 11509 7331 11543
rect 10241 11509 10275 11543
rect 10701 11509 10735 11543
rect 11161 11509 11195 11543
rect 11897 11509 11931 11543
rect 11989 11509 12023 11543
rect 16957 11509 16991 11543
rect 17325 11509 17359 11543
rect 19533 11509 19567 11543
rect 3249 11305 3283 11339
rect 3525 11305 3559 11339
rect 4077 11305 4111 11339
rect 5273 11305 5307 11339
rect 8769 11305 8803 11339
rect 9413 11305 9447 11339
rect 9873 11305 9907 11339
rect 15669 11305 15703 11339
rect 16589 11305 16623 11339
rect 17969 11305 18003 11339
rect 18797 11305 18831 11339
rect 19073 11305 19107 11339
rect 20545 11305 20579 11339
rect 6000 11237 6034 11271
rect 10425 11237 10459 11271
rect 12173 11237 12207 11271
rect 14473 11237 14507 11271
rect 15761 11237 15795 11271
rect 18061 11237 18095 11271
rect 1869 11169 1903 11203
rect 2136 11169 2170 11203
rect 4445 11169 4479 11203
rect 5089 11169 5123 11203
rect 5733 11169 5767 11203
rect 7389 11169 7423 11203
rect 7645 11169 7679 11203
rect 9229 11169 9263 11203
rect 9689 11169 9723 11203
rect 12449 11169 12483 11203
rect 12716 11169 12750 11203
rect 14565 11169 14599 11203
rect 16957 11169 16991 11203
rect 18613 11169 18647 11203
rect 19165 11169 19199 11203
rect 19432 11169 19466 11203
rect 1409 11101 1443 11135
rect 4537 11101 4571 11135
rect 4629 11101 4663 11135
rect 14657 11101 14691 11135
rect 15853 11101 15887 11135
rect 17049 11101 17083 11135
rect 17233 11101 17267 11135
rect 18245 11101 18279 11135
rect 19073 11101 19107 11135
rect 7113 11033 7147 11067
rect 13829 11033 13863 11067
rect 14105 11033 14139 11067
rect 17601 11033 17635 11067
rect 15301 10965 15335 10999
rect 3249 10761 3283 10795
rect 3709 10761 3743 10795
rect 3985 10761 4019 10795
rect 6377 10761 6411 10795
rect 7573 10761 7607 10795
rect 7665 10761 7699 10795
rect 8861 10761 8895 10795
rect 11161 10761 11195 10795
rect 11713 10761 11747 10795
rect 12081 10761 12115 10795
rect 14841 10761 14875 10795
rect 16957 10761 16991 10795
rect 19717 10761 19751 10795
rect 1869 10625 1903 10659
rect 4537 10625 4571 10659
rect 5733 10625 5767 10659
rect 3525 10557 3559 10591
rect 5089 10557 5123 10591
rect 5549 10557 5583 10591
rect 6193 10557 6227 10591
rect 2136 10489 2170 10523
rect 4445 10489 4479 10523
rect 7849 10693 7883 10727
rect 8493 10625 8527 10659
rect 9321 10625 9355 10659
rect 9505 10625 9539 10659
rect 13093 10625 13127 10659
rect 14013 10625 14047 10659
rect 15301 10625 15335 10659
rect 15485 10625 15519 10659
rect 16405 10625 16439 10659
rect 17509 10625 17543 10659
rect 20545 10625 20579 10659
rect 9781 10557 9815 10591
rect 11529 10557 11563 10591
rect 11897 10557 11931 10591
rect 18061 10557 18095 10591
rect 18328 10557 18362 10591
rect 20269 10557 20303 10591
rect 20361 10557 20395 10591
rect 10048 10489 10082 10523
rect 16313 10489 16347 10523
rect 17325 10489 17359 10523
rect 1409 10421 1443 10455
rect 4353 10421 4387 10455
rect 5181 10421 5215 10455
rect 5641 10421 5675 10455
rect 7573 10421 7607 10455
rect 8217 10421 8251 10455
rect 8309 10421 8343 10455
rect 9229 10421 9263 10455
rect 12449 10421 12483 10455
rect 12817 10421 12851 10455
rect 12909 10421 12943 10455
rect 13461 10421 13495 10455
rect 13829 10421 13863 10455
rect 13921 10421 13955 10455
rect 15209 10421 15243 10455
rect 15853 10421 15887 10455
rect 16221 10421 16255 10455
rect 17417 10421 17451 10455
rect 19441 10421 19475 10455
rect 19901 10421 19935 10455
rect 1685 10217 1719 10251
rect 3249 10217 3283 10251
rect 5457 10217 5491 10251
rect 7757 10217 7791 10251
rect 8217 10217 8251 10251
rect 10701 10217 10735 10251
rect 12817 10217 12851 10251
rect 14841 10217 14875 10251
rect 16773 10217 16807 10251
rect 17417 10217 17451 10251
rect 17785 10217 17819 10251
rect 20453 10217 20487 10251
rect 2421 10149 2455 10183
rect 6469 10149 6503 10183
rect 12909 10149 12943 10183
rect 19340 10149 19374 10183
rect 1501 10081 1535 10115
rect 2513 10081 2547 10115
rect 3065 10081 3099 10115
rect 4077 10081 4111 10115
rect 4333 10081 4367 10115
rect 6377 10081 6411 10115
rect 7205 10081 7239 10115
rect 7297 10081 7331 10115
rect 7941 10081 7975 10115
rect 8033 10081 8067 10115
rect 8953 10081 8987 10115
rect 9505 10081 9539 10115
rect 10057 10081 10091 10115
rect 11069 10081 11103 10115
rect 11897 10081 11931 10115
rect 13829 10081 13863 10115
rect 14657 10081 14691 10115
rect 15568 10081 15602 10115
rect 17877 10081 17911 10115
rect 18521 10081 18555 10115
rect 19073 10081 19107 10115
rect 2605 10013 2639 10047
rect 6561 10013 6595 10047
rect 7389 10013 7423 10047
rect 9045 10013 9079 10047
rect 9137 10013 9171 10047
rect 8585 9945 8619 9979
rect 10149 10013 10183 10047
rect 10333 10013 10367 10047
rect 11161 10013 11195 10047
rect 11345 10013 11379 10047
rect 13001 10013 13035 10047
rect 13921 10013 13955 10047
rect 14105 10013 14139 10047
rect 15301 10013 15335 10047
rect 17233 10013 17267 10047
rect 17969 10013 18003 10047
rect 10517 9945 10551 9979
rect 18705 9945 18739 9979
rect 2053 9877 2087 9911
rect 6009 9877 6043 9911
rect 6837 9877 6871 9911
rect 9505 9877 9539 9911
rect 9689 9877 9723 9911
rect 12081 9877 12115 9911
rect 12449 9877 12483 9911
rect 13461 9877 13495 9911
rect 16681 9877 16715 9911
rect 3157 9673 3191 9707
rect 10149 9673 10183 9707
rect 13829 9673 13863 9707
rect 1777 9605 1811 9639
rect 4077 9605 4111 9639
rect 5733 9605 5767 9639
rect 11989 9605 12023 9639
rect 14381 9605 14415 9639
rect 17233 9605 17267 9639
rect 18061 9605 18095 9639
rect 19073 9605 19107 9639
rect 20085 9605 20119 9639
rect 2697 9537 2731 9571
rect 3801 9537 3835 9571
rect 4629 9537 4663 9571
rect 5457 9537 5491 9571
rect 6193 9537 6227 9571
rect 6285 9537 6319 9571
rect 7113 9537 7147 9571
rect 11069 9537 11103 9571
rect 12449 9537 12483 9571
rect 14933 9537 14967 9571
rect 15393 9537 15427 9571
rect 15853 9537 15887 9571
rect 18705 9537 18739 9571
rect 19533 9537 19567 9571
rect 19625 9537 19659 9571
rect 20637 9537 20671 9571
rect 1593 9469 1627 9503
rect 3525 9469 3559 9503
rect 4445 9469 4479 9503
rect 7021 9469 7055 9503
rect 7380 9469 7414 9503
rect 8769 9469 8803 9503
rect 10885 9469 10919 9503
rect 11805 9469 11839 9503
rect 12716 9469 12750 9503
rect 14289 9469 14323 9503
rect 14749 9469 14783 9503
rect 18521 9469 18555 9503
rect 6101 9401 6135 9435
rect 9036 9401 9070 9435
rect 10793 9401 10827 9435
rect 16120 9401 16154 9435
rect 17509 9401 17543 9435
rect 18429 9401 18463 9435
rect 2145 9333 2179 9367
rect 2513 9333 2547 9367
rect 2605 9333 2639 9367
rect 3617 9333 3651 9367
rect 4537 9333 4571 9367
rect 4905 9333 4939 9367
rect 5273 9333 5307 9367
rect 5365 9333 5399 9367
rect 6837 9333 6871 9367
rect 8493 9333 8527 9367
rect 10425 9333 10459 9367
rect 14105 9333 14139 9367
rect 14841 9333 14875 9367
rect 19441 9333 19475 9367
rect 20453 9333 20487 9367
rect 20545 9333 20579 9367
rect 1961 9129 1995 9163
rect 2421 9129 2455 9163
rect 2973 9129 3007 9163
rect 4077 9129 4111 9163
rect 6469 9129 6503 9163
rect 7205 9129 7239 9163
rect 9229 9129 9263 9163
rect 10057 9129 10091 9163
rect 13001 9129 13035 9163
rect 14841 9129 14875 9163
rect 16313 9129 16347 9163
rect 19625 9129 19659 9163
rect 2329 9061 2363 9095
rect 3341 9061 3375 9095
rect 4445 9061 4479 9095
rect 5356 9061 5390 9095
rect 8116 9061 8150 9095
rect 10149 9061 10183 9095
rect 12909 9061 12943 9095
rect 14013 9061 14047 9095
rect 15761 9061 15795 9095
rect 16129 9061 16163 9095
rect 18512 9061 18546 9095
rect 1409 8993 1443 9027
rect 4537 8993 4571 9027
rect 5089 8993 5123 9027
rect 7113 8993 7147 9027
rect 7849 8993 7883 9027
rect 10885 8993 10919 9027
rect 11152 8993 11186 9027
rect 13921 8993 13955 9027
rect 14657 8993 14691 9027
rect 15117 8993 15151 9027
rect 15669 8993 15703 9027
rect 2605 8925 2639 8959
rect 3433 8925 3467 8959
rect 3525 8925 3559 8959
rect 4629 8925 4663 8959
rect 7297 8925 7331 8959
rect 10241 8925 10275 8959
rect 12449 8925 12483 8959
rect 13093 8925 13127 8959
rect 14105 8925 14139 8959
rect 1593 8857 1627 8891
rect 15853 8925 15887 8959
rect 16681 8993 16715 9027
rect 16773 8993 16807 9027
rect 17509 8993 17543 9027
rect 18245 8993 18279 9027
rect 19901 8993 19935 9027
rect 16865 8925 16899 8959
rect 17693 8925 17727 8959
rect 20085 8925 20119 8959
rect 15301 8857 15335 8891
rect 16129 8857 16163 8891
rect 6745 8789 6779 8823
rect 9689 8789 9723 8823
rect 12265 8789 12299 8823
rect 12449 8789 12483 8823
rect 12541 8789 12575 8823
rect 13553 8789 13587 8823
rect 15117 8789 15151 8823
rect 2421 8585 2455 8619
rect 3617 8585 3651 8619
rect 5733 8585 5767 8619
rect 12265 8585 12299 8619
rect 12449 8585 12483 8619
rect 19073 8585 19107 8619
rect 20085 8585 20119 8619
rect 5457 8517 5491 8551
rect 11989 8517 12023 8551
rect 1869 8449 1903 8483
rect 2053 8449 2087 8483
rect 2973 8449 3007 8483
rect 6193 8449 6227 8483
rect 6285 8449 6319 8483
rect 6837 8449 6871 8483
rect 9045 8449 9079 8483
rect 9413 8449 9447 8483
rect 10149 8449 10183 8483
rect 11069 8449 11103 8483
rect 1777 8381 1811 8415
rect 2789 8381 2823 8415
rect 3433 8381 3467 8415
rect 4077 8381 4111 8415
rect 8861 8381 8895 8415
rect 13461 8517 13495 8551
rect 14473 8517 14507 8551
rect 17509 8517 17543 8551
rect 18061 8517 18095 8551
rect 12909 8449 12943 8483
rect 13093 8449 13127 8483
rect 14105 8449 14139 8483
rect 14933 8449 14967 8483
rect 15025 8449 15059 8483
rect 18613 8449 18647 8483
rect 19533 8449 19567 8483
rect 19717 8449 19751 8483
rect 20637 8449 20671 8483
rect 11805 8381 11839 8415
rect 12265 8381 12299 8415
rect 12817 8381 12851 8415
rect 13921 8381 13955 8415
rect 15577 8381 15611 8415
rect 16129 8381 16163 8415
rect 16396 8381 16430 8415
rect 18521 8381 18555 8415
rect 20453 8381 20487 8415
rect 20545 8381 20579 8415
rect 2881 8313 2915 8347
rect 4344 8313 4378 8347
rect 7104 8313 7138 8347
rect 9413 8313 9447 8347
rect 9873 8313 9907 8347
rect 10885 8313 10919 8347
rect 14841 8313 14875 8347
rect 19441 8313 19475 8347
rect 1409 8245 1443 8279
rect 6101 8245 6135 8279
rect 8217 8245 8251 8279
rect 8493 8245 8527 8279
rect 8953 8245 8987 8279
rect 9505 8245 9539 8279
rect 9965 8245 9999 8279
rect 10517 8245 10551 8279
rect 10977 8245 11011 8279
rect 13829 8245 13863 8279
rect 15761 8245 15795 8279
rect 18429 8245 18463 8279
rect 2145 8041 2179 8075
rect 4077 8041 4111 8075
rect 4537 8041 4571 8075
rect 5089 8041 5123 8075
rect 5549 8041 5583 8075
rect 6101 8041 6135 8075
rect 6561 8041 6595 8075
rect 6929 8041 6963 8075
rect 9321 8041 9355 8075
rect 9413 8041 9447 8075
rect 12725 8041 12759 8075
rect 15301 8041 15335 8075
rect 15761 8041 15795 8075
rect 16681 8041 16715 8075
rect 18705 8041 18739 8075
rect 19717 8041 19751 8075
rect 4905 7973 4939 8007
rect 7297 7973 7331 8007
rect 1593 7905 1627 7939
rect 1869 7905 1903 7939
rect 2145 7905 2179 7939
rect 2596 7905 2630 7939
rect 4445 7905 4479 7939
rect 5457 7905 5491 7939
rect 6285 7905 6319 7939
rect 6377 7905 6411 7939
rect 8208 7905 8242 7939
rect 2329 7837 2363 7871
rect 4629 7837 4663 7871
rect 4905 7837 4939 7871
rect 5641 7837 5675 7871
rect 7389 7837 7423 7871
rect 7573 7837 7607 7871
rect 7941 7837 7975 7871
rect 3709 7769 3743 7803
rect 10876 7973 10910 8007
rect 12633 7973 12667 8007
rect 19073 7973 19107 8007
rect 9965 7905 9999 7939
rect 10609 7905 10643 7939
rect 12081 7905 12115 7939
rect 13461 7905 13495 7939
rect 13820 7905 13854 7939
rect 15669 7905 15703 7939
rect 16497 7905 16531 7939
rect 16865 7905 16899 7939
rect 17316 7905 17350 7939
rect 19165 7905 19199 7939
rect 20085 7905 20119 7939
rect 12817 7837 12851 7871
rect 13553 7837 13587 7871
rect 15853 7837 15887 7871
rect 17049 7837 17083 7871
rect 19349 7837 19383 7871
rect 20177 7837 20211 7871
rect 20269 7837 20303 7871
rect 13277 7769 13311 7803
rect 16865 7769 16899 7803
rect 9413 7701 9447 7735
rect 10149 7701 10183 7735
rect 11989 7701 12023 7735
rect 12173 7701 12207 7735
rect 12265 7701 12299 7735
rect 14933 7701 14967 7735
rect 18429 7701 18463 7735
rect 3157 7497 3191 7531
rect 5457 7497 5491 7531
rect 8493 7497 8527 7531
rect 8861 7497 8895 7531
rect 15117 7497 15151 7531
rect 16405 7497 16439 7531
rect 17601 7497 17635 7531
rect 18061 7497 18095 7531
rect 20085 7497 20119 7531
rect 5181 7429 5215 7463
rect 9689 7429 9723 7463
rect 13829 7429 13863 7463
rect 14105 7429 14139 7463
rect 19073 7429 19107 7463
rect 1777 7361 1811 7395
rect 3801 7361 3835 7395
rect 6101 7361 6135 7395
rect 9413 7361 9447 7395
rect 5825 7293 5859 7327
rect 7113 7293 7147 7327
rect 10333 7361 10367 7395
rect 10517 7361 10551 7395
rect 11437 7361 11471 7395
rect 11897 7361 11931 7395
rect 12449 7361 12483 7395
rect 14749 7361 14783 7395
rect 16037 7361 16071 7395
rect 16865 7361 16899 7395
rect 16957 7361 16991 7395
rect 18521 7361 18555 7395
rect 18613 7361 18647 7395
rect 19717 7361 19751 7395
rect 20637 7361 20671 7395
rect 10241 7293 10275 7327
rect 11253 7293 11287 7327
rect 14473 7293 14507 7327
rect 15301 7293 15335 7327
rect 17417 7293 17451 7327
rect 19441 7293 19475 7327
rect 2044 7225 2078 7259
rect 4068 7225 4102 7259
rect 5917 7225 5951 7259
rect 7380 7225 7414 7259
rect 9321 7225 9355 7259
rect 9689 7225 9723 7259
rect 11345 7225 11379 7259
rect 12716 7225 12750 7259
rect 14565 7225 14599 7259
rect 15853 7225 15887 7259
rect 18429 7225 18463 7259
rect 19533 7225 19567 7259
rect 20545 7225 20579 7259
rect 9229 7157 9263 7191
rect 9873 7157 9907 7191
rect 10885 7157 10919 7191
rect 15393 7157 15427 7191
rect 15761 7157 15795 7191
rect 16773 7157 16807 7191
rect 20453 7157 20487 7191
rect 2513 6953 2547 6987
rect 2605 6953 2639 6987
rect 4077 6953 4111 6987
rect 6653 6953 6687 6987
rect 7297 6953 7331 6987
rect 7573 6953 7607 6987
rect 7941 6953 7975 6987
rect 8585 6953 8619 6987
rect 9045 6953 9079 6987
rect 9781 6953 9815 6987
rect 10241 6953 10275 6987
rect 10333 6953 10367 6987
rect 11253 6953 11287 6987
rect 11805 6953 11839 6987
rect 11897 6953 11931 6987
rect 12357 6953 12391 6987
rect 15669 6953 15703 6987
rect 17877 6953 17911 6987
rect 18245 6953 18279 6987
rect 18337 6953 18371 6987
rect 4445 6885 4479 6919
rect 5457 6885 5491 6919
rect 8953 6885 8987 6919
rect 1593 6817 1627 6851
rect 3433 6817 3467 6851
rect 4537 6817 4571 6851
rect 6745 6817 6779 6851
rect 7481 6817 7515 6851
rect 12265 6885 12299 6919
rect 13277 6885 13311 6919
rect 14565 6885 14599 6919
rect 17233 6885 17267 6919
rect 19073 6885 19107 6919
rect 11805 6817 11839 6851
rect 14657 6817 14691 6851
rect 16313 6817 16347 6851
rect 19421 6817 19455 6851
rect 20913 6817 20947 6851
rect 2697 6749 2731 6783
rect 3341 6749 3375 6783
rect 4721 6749 4755 6783
rect 5549 6749 5583 6783
rect 5733 6749 5767 6783
rect 6193 6749 6227 6783
rect 6837 6749 6871 6783
rect 8033 6749 8067 6783
rect 8217 6749 8251 6783
rect 9229 6749 9263 6783
rect 9781 6749 9815 6783
rect 10425 6749 10459 6783
rect 11345 6749 11379 6783
rect 11529 6749 11563 6783
rect 12449 6749 12483 6783
rect 13369 6749 13403 6783
rect 13553 6749 13587 6783
rect 14105 6749 14139 6783
rect 14841 6749 14875 6783
rect 15761 6749 15795 6783
rect 15945 6749 15979 6783
rect 17325 6749 17359 6783
rect 17509 6749 17543 6783
rect 18429 6749 18463 6783
rect 19073 6749 19107 6783
rect 19165 6749 19199 6783
rect 1777 6681 1811 6715
rect 10885 6681 10919 6715
rect 14197 6681 14231 6715
rect 2145 6613 2179 6647
rect 3341 6613 3375 6647
rect 3617 6613 3651 6647
rect 5089 6613 5123 6647
rect 6285 6613 6319 6647
rect 9873 6613 9907 6647
rect 12909 6613 12943 6647
rect 15301 6613 15335 6647
rect 16497 6613 16531 6647
rect 16865 6613 16899 6647
rect 20545 6613 20579 6647
rect 1593 6409 1627 6443
rect 2881 6409 2915 6443
rect 14013 6409 14047 6443
rect 16957 6409 16991 6443
rect 20729 6409 20763 6443
rect 4997 6341 5031 6375
rect 5089 6341 5123 6375
rect 7665 6341 7699 6375
rect 16405 6341 16439 6375
rect 2513 6273 2547 6307
rect 3525 6273 3559 6307
rect 4537 6273 4571 6307
rect 4721 6273 4755 6307
rect 1409 6205 1443 6239
rect 3985 6205 4019 6239
rect 4445 6205 4479 6239
rect 5549 6273 5583 6307
rect 5733 6273 5767 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 8493 6273 8527 6307
rect 9781 6273 9815 6307
rect 15025 6273 15059 6307
rect 17417 6273 17451 6307
rect 17509 6273 17543 6307
rect 18521 6273 18555 6307
rect 18613 6273 18647 6307
rect 8217 6205 8251 6239
rect 9229 6205 9263 6239
rect 11805 6205 11839 6239
rect 12633 6205 12667 6239
rect 12900 6205 12934 6239
rect 14473 6205 14507 6239
rect 19349 6205 19383 6239
rect 3341 6137 3375 6171
rect 4997 6137 5031 6171
rect 8309 6137 8343 6171
rect 10026 6137 10060 6171
rect 15292 6137 15326 6171
rect 18429 6137 18463 6171
rect 19616 6137 19650 6171
rect 1961 6069 1995 6103
rect 2329 6069 2363 6103
rect 2421 6069 2455 6103
rect 3249 6069 3283 6103
rect 4077 6069 4111 6103
rect 5457 6069 5491 6103
rect 5917 6069 5951 6103
rect 6285 6069 6319 6103
rect 6837 6069 6871 6103
rect 7849 6069 7883 6103
rect 9413 6069 9447 6103
rect 11161 6069 11195 6103
rect 11989 6069 12023 6103
rect 14657 6069 14691 6103
rect 17325 6069 17359 6103
rect 18061 6069 18095 6103
rect 5733 5865 5767 5899
rect 7205 5865 7239 5899
rect 7665 5865 7699 5899
rect 8217 5865 8251 5899
rect 8585 5865 8619 5899
rect 11805 5865 11839 5899
rect 15485 5865 15519 5899
rect 15853 5865 15887 5899
rect 18797 5865 18831 5899
rect 19809 5865 19843 5899
rect 1869 5797 1903 5831
rect 4344 5797 4378 5831
rect 9956 5797 9990 5831
rect 11713 5797 11747 5831
rect 13360 5797 13394 5831
rect 18889 5797 18923 5831
rect 19901 5797 19935 5831
rect 1593 5729 1627 5763
rect 2596 5729 2630 5763
rect 4077 5729 4111 5763
rect 6561 5729 6595 5763
rect 6653 5729 6687 5763
rect 7573 5729 7607 5763
rect 9689 5729 9723 5763
rect 12541 5729 12575 5763
rect 13093 5729 13127 5763
rect 16773 5729 16807 5763
rect 17040 5729 17074 5763
rect 2329 5661 2363 5695
rect 6745 5661 6779 5695
rect 7849 5661 7883 5695
rect 8677 5661 8711 5695
rect 8769 5661 8803 5695
rect 11989 5661 12023 5695
rect 14749 5661 14783 5695
rect 15945 5661 15979 5695
rect 16037 5661 16071 5695
rect 18981 5661 19015 5695
rect 19993 5661 20027 5695
rect 12725 5593 12759 5627
rect 14473 5593 14507 5627
rect 18429 5593 18463 5627
rect 3709 5525 3743 5559
rect 5457 5525 5491 5559
rect 6193 5525 6227 5559
rect 11069 5525 11103 5559
rect 11345 5525 11379 5559
rect 18153 5525 18187 5559
rect 19441 5525 19475 5559
rect 1593 5321 1627 5355
rect 3617 5321 3651 5355
rect 5733 5321 5767 5355
rect 8217 5321 8251 5355
rect 17233 5321 17267 5355
rect 17785 5321 17819 5355
rect 20269 5321 20303 5355
rect 15669 5253 15703 5287
rect 1961 5185 1995 5219
rect 4169 5185 4203 5219
rect 5181 5185 5215 5219
rect 6377 5185 6411 5219
rect 11621 5185 11655 5219
rect 12909 5185 12943 5219
rect 13093 5185 13127 5219
rect 14381 5185 14415 5219
rect 15301 5185 15335 5219
rect 15393 5185 15427 5219
rect 1409 5117 1443 5151
rect 3985 5117 4019 5151
rect 4997 5117 5031 5151
rect 6101 5117 6135 5151
rect 6193 5117 6227 5151
rect 6837 5117 6871 5151
rect 8769 5117 8803 5151
rect 9036 5117 9070 5151
rect 10425 5117 10459 5151
rect 15209 5117 15243 5151
rect 15853 5185 15887 5219
rect 17509 5185 17543 5219
rect 17785 5185 17819 5219
rect 20729 5185 20763 5219
rect 18061 5117 18095 5151
rect 18889 5117 18923 5151
rect 20545 5117 20579 5151
rect 2228 5049 2262 5083
rect 7104 5049 7138 5083
rect 11345 5049 11379 5083
rect 15669 5049 15703 5083
rect 16098 5049 16132 5083
rect 19156 5049 19190 5083
rect 3341 4981 3375 5015
rect 4077 4981 4111 5015
rect 4629 4981 4663 5015
rect 5089 4981 5123 5015
rect 10149 4981 10183 5015
rect 10609 4981 10643 5015
rect 10977 4981 11011 5015
rect 11437 4981 11471 5015
rect 12449 4981 12483 5015
rect 12817 4981 12851 5015
rect 13277 4981 13311 5015
rect 13737 4981 13771 5015
rect 14105 4981 14139 5015
rect 14197 4981 14231 5015
rect 14841 4981 14875 5015
rect 18245 4981 18279 5015
rect 2881 4777 2915 4811
rect 3341 4777 3375 4811
rect 5089 4777 5123 4811
rect 7113 4777 7147 4811
rect 7389 4777 7423 4811
rect 7757 4777 7791 4811
rect 7849 4777 7883 4811
rect 8401 4777 8435 4811
rect 8769 4777 8803 4811
rect 10149 4777 10183 4811
rect 10517 4777 10551 4811
rect 10885 4777 10919 4811
rect 10977 4777 11011 4811
rect 13001 4777 13035 4811
rect 13921 4777 13955 4811
rect 14013 4777 14047 4811
rect 17417 4777 17451 4811
rect 17785 4777 17819 4811
rect 18245 4777 18279 4811
rect 20361 4777 20395 4811
rect 5978 4709 6012 4743
rect 11897 4709 11931 4743
rect 12909 4709 12943 4743
rect 13369 4709 13403 4743
rect 1501 4641 1535 4675
rect 1768 4641 1802 4675
rect 3433 4641 3467 4675
rect 4077 4641 4111 4675
rect 4997 4641 5031 4675
rect 5733 4641 5767 4675
rect 8861 4641 8895 4675
rect 9965 4641 9999 4675
rect 3617 4573 3651 4607
rect 5273 4573 5307 4607
rect 7941 4573 7975 4607
rect 8953 4573 8987 4607
rect 11069 4573 11103 4607
rect 11989 4573 12023 4607
rect 12173 4573 12207 4607
rect 13093 4573 13127 4607
rect 4629 4505 4663 4539
rect 17325 4709 17359 4743
rect 17877 4709 17911 4743
rect 14657 4641 14691 4675
rect 15669 4641 15703 4675
rect 16773 4641 16807 4675
rect 14105 4573 14139 4607
rect 15761 4573 15795 4607
rect 15945 4573 15979 4607
rect 16865 4573 16899 4607
rect 17049 4573 17083 4607
rect 17325 4573 17359 4607
rect 17969 4573 18003 4607
rect 13553 4505 13587 4539
rect 15301 4505 15335 4539
rect 18429 4641 18463 4675
rect 19533 4641 19567 4675
rect 20177 4641 20211 4675
rect 18705 4573 18739 4607
rect 19625 4573 19659 4607
rect 19717 4573 19751 4607
rect 20913 4573 20947 4607
rect 2973 4437 3007 4471
rect 4261 4437 4295 4471
rect 11529 4437 11563 4471
rect 12541 4437 12575 4471
rect 13369 4437 13403 4471
rect 14841 4437 14875 4471
rect 16405 4437 16439 4471
rect 18245 4437 18279 4471
rect 19165 4437 19199 4471
rect 14657 4233 14691 4267
rect 14749 4233 14783 4267
rect 19717 4233 19751 4267
rect 4721 4165 4755 4199
rect 6837 4165 6871 4199
rect 8309 4165 8343 4199
rect 12449 4165 12483 4199
rect 14473 4165 14507 4199
rect 2237 4097 2271 4131
rect 3157 4097 3191 4131
rect 3341 4097 3375 4131
rect 4261 4097 4295 4131
rect 5641 4097 5675 4131
rect 7297 4097 7331 4131
rect 7481 4097 7515 4131
rect 11713 4097 11747 4131
rect 11805 4097 11839 4131
rect 20913 4165 20947 4199
rect 13001 4097 13035 4131
rect 14657 4097 14691 4131
rect 15301 4097 15335 4131
rect 16957 4097 16991 4131
rect 18061 4097 18095 4131
rect 20361 4097 20395 4131
rect 2145 4029 2179 4063
rect 4537 4029 4571 4063
rect 6193 4029 6227 4063
rect 7205 4029 7239 4063
rect 8125 4029 8159 4063
rect 8677 4029 8711 4063
rect 10333 4029 10367 4063
rect 12449 4029 12483 4063
rect 12541 4029 12575 4063
rect 2053 3961 2087 3995
rect 3065 3961 3099 3995
rect 5365 3961 5399 3995
rect 5457 3961 5491 3995
rect 8944 3961 8978 3995
rect 10609 3961 10643 3995
rect 13093 4029 13127 4063
rect 15761 4029 15795 4063
rect 17325 4029 17359 4063
rect 17509 4029 17543 4063
rect 20177 4029 20211 4063
rect 20729 4029 20763 4063
rect 13360 3961 13394 3995
rect 16037 3961 16071 3995
rect 18306 3961 18340 3995
rect 1685 3893 1719 3927
rect 2697 3893 2731 3927
rect 3709 3893 3743 3927
rect 4077 3893 4111 3927
rect 4169 3893 4203 3927
rect 4997 3893 5031 3927
rect 6377 3893 6411 3927
rect 10057 3893 10091 3927
rect 11253 3893 11287 3927
rect 11621 3893 11655 3927
rect 12725 3893 12759 3927
rect 13001 3893 13035 3927
rect 15117 3893 15151 3927
rect 15209 3893 15243 3927
rect 16313 3893 16347 3927
rect 16681 3893 16715 3927
rect 16773 3893 16807 3927
rect 19441 3893 19475 3927
rect 20085 3893 20119 3927
rect 2053 3689 2087 3723
rect 3525 3689 3559 3723
rect 4813 3689 4847 3723
rect 5825 3689 5859 3723
rect 7021 3689 7055 3723
rect 7665 3689 7699 3723
rect 9689 3689 9723 3723
rect 10149 3689 10183 3723
rect 12449 3689 12483 3723
rect 12817 3689 12851 3723
rect 13461 3689 13495 3723
rect 15301 3689 15335 3723
rect 17049 3689 17083 3723
rect 18521 3689 18555 3723
rect 1685 3621 1719 3655
rect 7113 3621 7147 3655
rect 8033 3621 8067 3655
rect 9137 3621 9171 3655
rect 10057 3621 10091 3655
rect 11060 3621 11094 3655
rect 12909 3621 12943 3655
rect 1409 3553 1443 3587
rect 2145 3553 2179 3587
rect 2412 3553 2446 3587
rect 3617 3553 3651 3587
rect 4905 3553 4939 3587
rect 8125 3553 8159 3587
rect 8861 3553 8895 3587
rect 13829 3553 13863 3587
rect 14841 3553 14875 3587
rect 15669 3553 15703 3587
rect 16405 3553 16439 3587
rect 16681 3553 16715 3587
rect 17408 3621 17442 3655
rect 20269 3621 20303 3655
rect 19165 3553 19199 3587
rect 20177 3553 20211 3587
rect 5089 3485 5123 3519
rect 5917 3485 5951 3519
rect 6009 3485 6043 3519
rect 7297 3485 7331 3519
rect 8309 3485 8343 3519
rect 10241 3485 10275 3519
rect 10793 3485 10827 3519
rect 13001 3485 13035 3519
rect 13921 3485 13955 3519
rect 14013 3485 14047 3519
rect 15761 3485 15795 3519
rect 15945 3485 15979 3519
rect 17049 3485 17083 3519
rect 17141 3485 17175 3519
rect 19257 3485 19291 3519
rect 19349 3485 19383 3519
rect 20361 3485 20395 3519
rect 3801 3417 3835 3451
rect 4261 3417 4295 3451
rect 4445 3417 4479 3451
rect 16129 3417 16163 3451
rect 19809 3417 19843 3451
rect 5273 3349 5307 3383
rect 5457 3349 5491 3383
rect 6653 3349 6687 3383
rect 12173 3349 12207 3383
rect 18797 3349 18831 3383
rect 5733 3145 5767 3179
rect 8217 3145 8251 3179
rect 14013 3145 14047 3179
rect 17233 3145 17267 3179
rect 18153 3145 18187 3179
rect 18245 3145 18279 3179
rect 19533 3145 19567 3179
rect 1685 3077 1719 3111
rect 5273 3077 5307 3111
rect 12081 3077 12115 3111
rect 12449 3077 12483 3111
rect 2237 3009 2271 3043
rect 3157 3009 3191 3043
rect 3341 3009 3375 3043
rect 3893 3009 3927 3043
rect 6285 3009 6319 3043
rect 8493 3009 8527 3043
rect 10701 3009 10735 3043
rect 12909 3009 12943 3043
rect 13093 3009 13127 3043
rect 13645 3009 13679 3043
rect 3525 2941 3559 2975
rect 5365 2941 5399 2975
rect 6101 2941 6135 2975
rect 6837 2941 6871 2975
rect 8760 2941 8794 2975
rect 10149 2941 10183 2975
rect 10968 2941 11002 2975
rect 12817 2941 12851 2975
rect 13461 2941 13495 2975
rect 14105 3009 14139 3043
rect 14933 3009 14967 3043
rect 18153 3009 18187 3043
rect 18797 3009 18831 3043
rect 19993 3009 20027 3043
rect 20085 3009 20119 3043
rect 15209 2941 15243 2975
rect 15853 2941 15887 2975
rect 19901 2941 19935 2975
rect 20545 2941 20579 2975
rect 4160 2873 4194 2907
rect 7104 2873 7138 2907
rect 14013 2873 14047 2907
rect 14749 2873 14783 2907
rect 15485 2873 15519 2907
rect 16098 2873 16132 2907
rect 20821 2873 20855 2907
rect 2053 2805 2087 2839
rect 2145 2805 2179 2839
rect 2697 2805 2731 2839
rect 3065 2805 3099 2839
rect 3709 2805 3743 2839
rect 5549 2805 5583 2839
rect 6193 2805 6227 2839
rect 9873 2805 9907 2839
rect 10333 2805 10367 2839
rect 14381 2805 14415 2839
rect 14841 2805 14875 2839
rect 18613 2805 18647 2839
rect 18705 2805 18739 2839
rect 1961 2601 1995 2635
rect 2329 2601 2363 2635
rect 5917 2601 5951 2635
rect 6929 2601 6963 2635
rect 8309 2601 8343 2635
rect 10241 2601 10275 2635
rect 11161 2601 11195 2635
rect 12633 2601 12667 2635
rect 13001 2601 13035 2635
rect 14841 2601 14875 2635
rect 16681 2601 16715 2635
rect 17233 2601 17267 2635
rect 18705 2601 18739 2635
rect 19349 2601 19383 2635
rect 19717 2601 19751 2635
rect 4690 2533 4724 2567
rect 6377 2533 6411 2567
rect 10701 2533 10735 2567
rect 13921 2533 13955 2567
rect 14749 2533 14783 2567
rect 16589 2533 16623 2567
rect 17601 2533 17635 2567
rect 18797 2533 18831 2567
rect 20637 2533 20671 2567
rect 2421 2465 2455 2499
rect 3525 2465 3559 2499
rect 4445 2465 4479 2499
rect 6285 2465 6319 2499
rect 7297 2465 7331 2499
rect 9137 2465 9171 2499
rect 10149 2465 10183 2499
rect 2605 2397 2639 2431
rect 3065 2397 3099 2431
rect 3617 2397 3651 2431
rect 3801 2397 3835 2431
rect 6469 2397 6503 2431
rect 7389 2397 7423 2431
rect 7573 2397 7607 2431
rect 8401 2397 8435 2431
rect 8585 2397 8619 2431
rect 10425 2397 10459 2431
rect 3157 2329 3191 2363
rect 4353 2329 4387 2363
rect 5825 2329 5859 2363
rect 7941 2329 7975 2363
rect 11805 2465 11839 2499
rect 13645 2465 13679 2499
rect 15669 2465 15703 2499
rect 17693 2465 17727 2499
rect 20361 2465 20395 2499
rect 11253 2397 11287 2431
rect 11345 2397 11379 2431
rect 11989 2397 12023 2431
rect 13093 2397 13127 2431
rect 13185 2397 13219 2431
rect 15025 2397 15059 2431
rect 16865 2397 16899 2431
rect 17785 2397 17819 2431
rect 18889 2397 18923 2431
rect 19809 2397 19843 2431
rect 19993 2397 20027 2431
rect 14381 2329 14415 2363
rect 15853 2329 15887 2363
rect 18337 2329 18371 2363
rect 9321 2261 9355 2295
rect 9781 2261 9815 2295
rect 10701 2261 10735 2295
rect 10793 2261 10827 2295
rect 16221 2261 16255 2295
rect 11161 1785 11195 1819
rect 11161 1649 11195 1683
rect 8769 1581 8803 1615
rect 8769 1377 8803 1411
<< metal1 >>
rect 4062 21360 4068 21412
rect 4120 21400 4126 21412
rect 10502 21400 10508 21412
rect 4120 21372 10508 21400
rect 4120 21360 4126 21372
rect 10502 21360 10508 21372
rect 10560 21360 10566 21412
rect 3694 21088 3700 21140
rect 3752 21128 3758 21140
rect 8754 21128 8760 21140
rect 3752 21100 8760 21128
rect 3752 21088 3758 21100
rect 8754 21088 8760 21100
rect 8812 21088 8818 21140
rect 14458 20680 14464 20732
rect 14516 20720 14522 20732
rect 18138 20720 18144 20732
rect 14516 20692 18144 20720
rect 14516 20680 14522 20692
rect 18138 20680 18144 20692
rect 18196 20680 18202 20732
rect 1670 20476 1676 20528
rect 1728 20516 1734 20528
rect 4246 20516 4252 20528
rect 1728 20488 4252 20516
rect 1728 20476 1734 20488
rect 4246 20476 4252 20488
rect 4304 20476 4310 20528
rect 2590 20408 2596 20460
rect 2648 20448 2654 20460
rect 8570 20448 8576 20460
rect 2648 20420 8576 20448
rect 2648 20408 2654 20420
rect 8570 20408 8576 20420
rect 8628 20408 8634 20460
rect 4706 20340 4712 20392
rect 4764 20380 4770 20392
rect 5166 20380 5172 20392
rect 4764 20352 5172 20380
rect 4764 20340 4770 20352
rect 5166 20340 5172 20352
rect 5224 20340 5230 20392
rect 9398 20340 9404 20392
rect 9456 20380 9462 20392
rect 10778 20380 10784 20392
rect 9456 20352 10784 20380
rect 9456 20340 9462 20352
rect 10778 20340 10784 20352
rect 10836 20340 10842 20392
rect 14366 20340 14372 20392
rect 14424 20380 14430 20392
rect 21450 20380 21456 20392
rect 14424 20352 21456 20380
rect 14424 20340 14430 20352
rect 21450 20340 21456 20352
rect 21508 20340 21514 20392
rect 3786 20272 3792 20324
rect 3844 20312 3850 20324
rect 10870 20312 10876 20324
rect 3844 20284 10876 20312
rect 3844 20272 3850 20284
rect 10870 20272 10876 20284
rect 10928 20272 10934 20324
rect 19610 20272 19616 20324
rect 19668 20312 19674 20324
rect 20346 20312 20352 20324
rect 19668 20284 20352 20312
rect 19668 20272 19674 20284
rect 20346 20272 20352 20284
rect 20404 20272 20410 20324
rect 4062 20204 4068 20256
rect 4120 20244 4126 20256
rect 13170 20244 13176 20256
rect 4120 20216 13176 20244
rect 4120 20204 4126 20216
rect 13170 20204 13176 20216
rect 13228 20204 13234 20256
rect 13722 20204 13728 20256
rect 13780 20244 13786 20256
rect 19058 20244 19064 20256
rect 13780 20216 19064 20244
rect 13780 20204 13786 20216
rect 19058 20204 19064 20216
rect 19116 20204 19122 20256
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 3786 20040 3792 20052
rect 1688 20012 3792 20040
rect 1688 19913 1716 20012
rect 3786 20000 3792 20012
rect 3844 20000 3850 20052
rect 4065 20043 4123 20049
rect 4065 20009 4077 20043
rect 4111 20040 4123 20043
rect 6638 20040 6644 20052
rect 4111 20012 6644 20040
rect 4111 20009 4123 20012
rect 4065 20003 4123 20009
rect 6638 20000 6644 20012
rect 6696 20000 6702 20052
rect 10226 20040 10232 20052
rect 10187 20012 10232 20040
rect 10226 20000 10232 20012
rect 10284 20000 10290 20052
rect 14366 20040 14372 20052
rect 11072 20012 14372 20040
rect 2498 19932 2504 19984
rect 2556 19972 2562 19984
rect 3513 19975 3571 19981
rect 2556 19944 3372 19972
rect 2556 19932 2562 19944
rect 1673 19907 1731 19913
rect 1673 19873 1685 19907
rect 1719 19873 1731 19907
rect 1673 19867 1731 19873
rect 2409 19907 2467 19913
rect 2409 19873 2421 19907
rect 2455 19904 2467 19907
rect 2590 19904 2596 19916
rect 2455 19876 2596 19904
rect 2455 19873 2467 19876
rect 2409 19867 2467 19873
rect 2590 19864 2596 19876
rect 2648 19864 2654 19916
rect 3234 19904 3240 19916
rect 3195 19876 3240 19904
rect 3234 19864 3240 19876
rect 3292 19864 3298 19916
rect 3344 19904 3372 19944
rect 3513 19941 3525 19975
rect 3559 19972 3571 19975
rect 6365 19975 6423 19981
rect 3559 19944 6316 19972
rect 3559 19941 3571 19944
rect 3513 19935 3571 19941
rect 4433 19907 4491 19913
rect 4433 19904 4445 19907
rect 3344 19876 4445 19904
rect 4433 19873 4445 19876
rect 4479 19904 4491 19907
rect 4982 19904 4988 19916
rect 4479 19876 4988 19904
rect 4479 19873 4491 19876
rect 4433 19867 4491 19873
rect 4982 19864 4988 19876
rect 5040 19864 5046 19916
rect 5442 19904 5448 19916
rect 5184 19876 5448 19904
rect 1854 19836 1860 19848
rect 1815 19808 1860 19836
rect 1854 19796 1860 19808
rect 1912 19796 1918 19848
rect 2685 19839 2743 19845
rect 2685 19805 2697 19839
rect 2731 19836 2743 19839
rect 2774 19836 2780 19848
rect 2731 19808 2780 19836
rect 2731 19805 2743 19808
rect 2685 19799 2743 19805
rect 2774 19796 2780 19808
rect 2832 19796 2838 19848
rect 4246 19796 4252 19848
rect 4304 19836 4310 19848
rect 4525 19839 4583 19845
rect 4525 19836 4537 19839
rect 4304 19808 4537 19836
rect 4304 19796 4310 19808
rect 4525 19805 4537 19808
rect 4571 19805 4583 19839
rect 4706 19836 4712 19848
rect 4667 19808 4712 19836
rect 4525 19799 4583 19805
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 4154 19728 4160 19780
rect 4212 19768 4218 19780
rect 5184 19768 5212 19876
rect 5442 19864 5448 19876
rect 5500 19864 5506 19916
rect 6086 19904 6092 19916
rect 6047 19876 6092 19904
rect 6086 19864 6092 19876
rect 6144 19864 6150 19916
rect 6288 19904 6316 19944
rect 6365 19941 6377 19975
rect 6411 19972 6423 19975
rect 6914 19972 6920 19984
rect 6411 19944 6920 19972
rect 6411 19941 6423 19944
rect 6365 19935 6423 19941
rect 6914 19932 6920 19944
rect 6972 19932 6978 19984
rect 7098 19932 7104 19984
rect 7156 19932 7162 19984
rect 7466 19932 7472 19984
rect 7524 19972 7530 19984
rect 8941 19975 8999 19981
rect 8941 19972 8953 19975
rect 7524 19944 8953 19972
rect 7524 19932 7530 19944
rect 8941 19941 8953 19944
rect 8987 19941 8999 19975
rect 8941 19935 8999 19941
rect 9674 19932 9680 19984
rect 9732 19972 9738 19984
rect 10962 19972 10968 19984
rect 9732 19944 10968 19972
rect 9732 19932 9738 19944
rect 10962 19932 10968 19944
rect 11020 19932 11026 19984
rect 11072 19981 11100 20012
rect 14366 20000 14372 20012
rect 14424 20000 14430 20052
rect 15013 20043 15071 20049
rect 15013 20009 15025 20043
rect 15059 20040 15071 20043
rect 18046 20040 18052 20052
rect 15059 20012 18052 20040
rect 15059 20009 15071 20012
rect 15013 20003 15071 20009
rect 18046 20000 18052 20012
rect 18104 20000 18110 20052
rect 18141 20043 18199 20049
rect 18141 20009 18153 20043
rect 18187 20040 18199 20043
rect 22554 20040 22560 20052
rect 18187 20012 22560 20040
rect 18187 20009 18199 20012
rect 18141 20003 18199 20009
rect 22554 20000 22560 20012
rect 22612 20000 22618 20052
rect 11057 19975 11115 19981
rect 11057 19941 11069 19975
rect 11103 19941 11115 19975
rect 11057 19935 11115 19941
rect 11885 19975 11943 19981
rect 11885 19941 11897 19975
rect 11931 19972 11943 19975
rect 12986 19972 12992 19984
rect 11931 19944 12992 19972
rect 11931 19941 11943 19944
rect 11885 19935 11943 19941
rect 12986 19932 12992 19944
rect 13044 19932 13050 19984
rect 14093 19975 14151 19981
rect 14093 19941 14105 19975
rect 14139 19972 14151 19975
rect 16942 19972 16948 19984
rect 14139 19944 16948 19972
rect 14139 19941 14151 19944
rect 14093 19935 14151 19941
rect 16942 19932 16948 19944
rect 17000 19932 17006 19984
rect 17037 19975 17095 19981
rect 17037 19941 17049 19975
rect 17083 19972 17095 19975
rect 17954 19972 17960 19984
rect 17083 19944 17960 19972
rect 17083 19941 17095 19944
rect 17037 19935 17095 19941
rect 17954 19932 17960 19944
rect 18012 19932 18018 19984
rect 19886 19972 19892 19984
rect 18064 19944 19748 19972
rect 19847 19944 19892 19972
rect 6730 19904 6736 19916
rect 6288 19876 6736 19904
rect 6730 19864 6736 19876
rect 6788 19864 6794 19916
rect 7116 19904 7144 19932
rect 6932 19876 7144 19904
rect 7184 19907 7242 19913
rect 5258 19796 5264 19848
rect 5316 19836 5322 19848
rect 6932 19845 6960 19876
rect 7184 19873 7196 19907
rect 7230 19904 7242 19907
rect 8386 19904 8392 19916
rect 7230 19876 8392 19904
rect 7230 19873 7242 19876
rect 7184 19867 7242 19873
rect 8386 19864 8392 19876
rect 8444 19864 8450 19916
rect 10134 19904 10140 19916
rect 10095 19876 10140 19904
rect 10134 19864 10140 19876
rect 10192 19864 10198 19916
rect 10318 19904 10324 19916
rect 10231 19876 10324 19904
rect 5537 19839 5595 19845
rect 5537 19836 5549 19839
rect 5316 19808 5549 19836
rect 5316 19796 5322 19808
rect 5537 19805 5549 19808
rect 5583 19805 5595 19839
rect 5537 19799 5595 19805
rect 5721 19839 5779 19845
rect 5721 19805 5733 19839
rect 5767 19836 5779 19839
rect 6917 19839 6975 19845
rect 5767 19808 6408 19836
rect 5767 19805 5779 19808
rect 5721 19799 5779 19805
rect 4212 19740 5212 19768
rect 4212 19728 4218 19740
rect 5350 19728 5356 19780
rect 5408 19768 5414 19780
rect 5736 19768 5764 19799
rect 5408 19740 5764 19768
rect 5408 19728 5414 19740
rect 5077 19703 5135 19709
rect 5077 19669 5089 19703
rect 5123 19700 5135 19703
rect 6178 19700 6184 19712
rect 5123 19672 6184 19700
rect 5123 19669 5135 19672
rect 5077 19663 5135 19669
rect 6178 19660 6184 19672
rect 6236 19660 6242 19712
rect 6380 19700 6408 19808
rect 6917 19805 6929 19839
rect 6963 19805 6975 19839
rect 9030 19836 9036 19848
rect 8991 19808 9036 19836
rect 6917 19799 6975 19805
rect 9030 19796 9036 19808
rect 9088 19796 9094 19848
rect 9125 19839 9183 19845
rect 9125 19805 9137 19839
rect 9171 19805 9183 19839
rect 9125 19799 9183 19805
rect 8386 19728 8392 19780
rect 8444 19768 8450 19780
rect 9140 19768 9168 19799
rect 8444 19740 9168 19768
rect 8444 19728 8450 19740
rect 9214 19728 9220 19780
rect 9272 19768 9278 19780
rect 10244 19768 10272 19876
rect 10318 19864 10324 19876
rect 10376 19904 10382 19916
rect 10781 19907 10839 19913
rect 10376 19876 10456 19904
rect 10376 19864 10382 19876
rect 10428 19845 10456 19876
rect 10781 19873 10793 19907
rect 10827 19904 10839 19907
rect 10870 19904 10876 19916
rect 10827 19876 10876 19904
rect 10827 19873 10839 19876
rect 10781 19867 10839 19873
rect 10870 19864 10876 19876
rect 10928 19864 10934 19916
rect 12618 19904 12624 19916
rect 12579 19876 12624 19904
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 14829 19907 14887 19913
rect 14829 19873 14841 19907
rect 14875 19904 14887 19907
rect 15841 19907 15899 19913
rect 14875 19876 15792 19904
rect 14875 19873 14887 19876
rect 14829 19867 14887 19873
rect 10413 19839 10471 19845
rect 10413 19805 10425 19839
rect 10459 19805 10471 19839
rect 10413 19799 10471 19805
rect 11977 19839 12035 19845
rect 11977 19805 11989 19839
rect 12023 19805 12035 19839
rect 11977 19799 12035 19805
rect 9272 19740 10272 19768
rect 11992 19768 12020 19799
rect 12066 19796 12072 19848
rect 12124 19836 12130 19848
rect 12897 19839 12955 19845
rect 12124 19808 12169 19836
rect 12124 19796 12130 19808
rect 12897 19805 12909 19839
rect 12943 19836 12955 19839
rect 13446 19836 13452 19848
rect 12943 19808 13452 19836
rect 12943 19805 12955 19808
rect 12897 19799 12955 19805
rect 13446 19796 13452 19808
rect 13504 19796 13510 19848
rect 14182 19836 14188 19848
rect 14143 19808 14188 19836
rect 14182 19796 14188 19808
rect 14240 19796 14246 19848
rect 14369 19839 14427 19845
rect 14369 19805 14381 19839
rect 14415 19836 14427 19839
rect 15102 19836 15108 19848
rect 14415 19808 15108 19836
rect 14415 19805 14427 19808
rect 14369 19799 14427 19805
rect 15102 19796 15108 19808
rect 15160 19796 15166 19848
rect 13722 19768 13728 19780
rect 11992 19740 12940 19768
rect 13683 19740 13728 19768
rect 9272 19728 9278 19740
rect 12912 19712 12940 19740
rect 13722 19728 13728 19740
rect 13780 19728 13786 19780
rect 8297 19703 8355 19709
rect 8297 19700 8309 19703
rect 6380 19672 8309 19700
rect 8297 19669 8309 19672
rect 8343 19669 8355 19703
rect 8297 19663 8355 19669
rect 8573 19703 8631 19709
rect 8573 19669 8585 19703
rect 8619 19700 8631 19703
rect 9674 19700 9680 19712
rect 8619 19672 9680 19700
rect 8619 19669 8631 19672
rect 8573 19663 8631 19669
rect 9674 19660 9680 19672
rect 9732 19660 9738 19712
rect 9766 19660 9772 19712
rect 9824 19700 9830 19712
rect 9824 19672 9869 19700
rect 9824 19660 9830 19672
rect 10042 19660 10048 19712
rect 10100 19700 10106 19712
rect 10594 19700 10600 19712
rect 10100 19672 10600 19700
rect 10100 19660 10106 19672
rect 10594 19660 10600 19672
rect 10652 19660 10658 19712
rect 11517 19703 11575 19709
rect 11517 19669 11529 19703
rect 11563 19700 11575 19703
rect 12802 19700 12808 19712
rect 11563 19672 12808 19700
rect 11563 19669 11575 19672
rect 11517 19663 11575 19669
rect 12802 19660 12808 19672
rect 12860 19660 12866 19712
rect 12894 19660 12900 19712
rect 12952 19660 12958 19712
rect 15194 19660 15200 19712
rect 15252 19700 15258 19712
rect 15473 19703 15531 19709
rect 15473 19700 15485 19703
rect 15252 19672 15485 19700
rect 15252 19660 15258 19672
rect 15473 19669 15485 19672
rect 15519 19669 15531 19703
rect 15764 19700 15792 19876
rect 15841 19873 15853 19907
rect 15887 19904 15899 19907
rect 16574 19904 16580 19916
rect 15887 19876 16580 19904
rect 15887 19873 15899 19876
rect 15841 19867 15899 19873
rect 16574 19864 16580 19876
rect 16632 19864 16638 19916
rect 16758 19904 16764 19916
rect 16719 19876 16764 19904
rect 16758 19864 16764 19876
rect 16816 19864 16822 19916
rect 17494 19904 17500 19916
rect 17455 19876 17500 19904
rect 17494 19864 17500 19876
rect 17552 19904 17558 19916
rect 18064 19904 18092 19944
rect 17552 19876 18092 19904
rect 18325 19907 18383 19913
rect 17552 19864 17558 19876
rect 18325 19873 18337 19907
rect 18371 19873 18383 19907
rect 18874 19904 18880 19916
rect 18835 19876 18880 19904
rect 18325 19867 18383 19873
rect 15930 19836 15936 19848
rect 15891 19808 15936 19836
rect 15930 19796 15936 19808
rect 15988 19796 15994 19848
rect 16114 19836 16120 19848
rect 16075 19808 16120 19836
rect 16114 19796 16120 19808
rect 16172 19796 16178 19848
rect 17773 19839 17831 19845
rect 17773 19805 17785 19839
rect 17819 19836 17831 19839
rect 18141 19839 18199 19845
rect 18141 19836 18153 19839
rect 17819 19808 18153 19836
rect 17819 19805 17831 19808
rect 17773 19799 17831 19805
rect 18141 19805 18153 19808
rect 18187 19805 18199 19839
rect 18141 19799 18199 19805
rect 16206 19728 16212 19780
rect 16264 19768 16270 19780
rect 18340 19768 18368 19867
rect 18874 19864 18880 19876
rect 18932 19864 18938 19916
rect 19610 19904 19616 19916
rect 19571 19876 19616 19904
rect 19610 19864 19616 19876
rect 19668 19864 19674 19916
rect 19720 19904 19748 19944
rect 19886 19932 19892 19944
rect 19944 19932 19950 19984
rect 20622 19972 20628 19984
rect 20583 19944 20628 19972
rect 20622 19932 20628 19944
rect 20680 19932 20686 19984
rect 20346 19904 20352 19916
rect 19720 19876 20352 19904
rect 20346 19864 20352 19876
rect 20404 19864 20410 19916
rect 19153 19839 19211 19845
rect 19153 19805 19165 19839
rect 19199 19836 19211 19839
rect 22186 19836 22192 19848
rect 19199 19808 22192 19836
rect 19199 19805 19211 19808
rect 19153 19799 19211 19805
rect 22186 19796 22192 19808
rect 22244 19796 22250 19848
rect 16264 19740 18368 19768
rect 16264 19728 16270 19740
rect 17126 19700 17132 19712
rect 15764 19672 17132 19700
rect 15473 19663 15531 19669
rect 17126 19660 17132 19672
rect 17184 19660 17190 19712
rect 18509 19703 18567 19709
rect 18509 19669 18521 19703
rect 18555 19700 18567 19703
rect 18598 19700 18604 19712
rect 18555 19672 18604 19700
rect 18555 19669 18567 19672
rect 18509 19663 18567 19669
rect 18598 19660 18604 19672
rect 18656 19660 18662 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 5810 19496 5816 19508
rect 4448 19468 5816 19496
rect 3326 19428 3332 19440
rect 3287 19400 3332 19428
rect 3326 19388 3332 19400
rect 3384 19388 3390 19440
rect 3786 19428 3792 19440
rect 3747 19400 3792 19428
rect 3786 19388 3792 19400
rect 3844 19388 3850 19440
rect 2608 19332 3740 19360
rect 1673 19295 1731 19301
rect 1673 19261 1685 19295
rect 1719 19261 1731 19295
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1673 19255 1731 19261
rect 934 19184 940 19236
rect 992 19224 998 19236
rect 1578 19224 1584 19236
rect 992 19196 1584 19224
rect 992 19184 998 19196
rect 1578 19184 1584 19196
rect 1636 19184 1642 19236
rect 1688 19224 1716 19255
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2406 19292 2412 19304
rect 2367 19264 2412 19292
rect 2406 19252 2412 19264
rect 2464 19252 2470 19304
rect 2498 19224 2504 19236
rect 1688 19196 2504 19224
rect 2498 19184 2504 19196
rect 2556 19184 2562 19236
rect 1302 19116 1308 19168
rect 1360 19156 1366 19168
rect 2608 19156 2636 19332
rect 2685 19295 2743 19301
rect 2685 19261 2697 19295
rect 2731 19292 2743 19295
rect 2866 19292 2872 19304
rect 2731 19264 2872 19292
rect 2731 19261 2743 19264
rect 2685 19255 2743 19261
rect 2866 19252 2872 19264
rect 2924 19252 2930 19304
rect 3050 19252 3056 19304
rect 3108 19292 3114 19304
rect 3145 19295 3203 19301
rect 3145 19292 3157 19295
rect 3108 19264 3157 19292
rect 3108 19252 3114 19264
rect 3145 19261 3157 19264
rect 3191 19261 3203 19295
rect 3145 19255 3203 19261
rect 3712 19224 3740 19332
rect 4062 19320 4068 19372
rect 4120 19360 4126 19372
rect 4338 19360 4344 19372
rect 4120 19332 4344 19360
rect 4120 19320 4126 19332
rect 4338 19320 4344 19332
rect 4396 19320 4402 19372
rect 4448 19369 4476 19468
rect 5810 19456 5816 19468
rect 5868 19456 5874 19508
rect 7190 19456 7196 19508
rect 7248 19496 7254 19508
rect 8386 19496 8392 19508
rect 7248 19468 8248 19496
rect 8347 19468 8392 19496
rect 7248 19456 7254 19468
rect 4433 19363 4491 19369
rect 4433 19329 4445 19363
rect 4479 19329 4491 19363
rect 8220 19360 8248 19468
rect 8386 19456 8392 19468
rect 8444 19456 8450 19508
rect 9490 19456 9496 19508
rect 9548 19496 9554 19508
rect 11606 19496 11612 19508
rect 9548 19468 11612 19496
rect 9548 19456 9554 19468
rect 11606 19456 11612 19468
rect 11664 19456 11670 19508
rect 12434 19496 12440 19508
rect 12395 19468 12440 19496
rect 12434 19456 12440 19468
rect 12492 19456 12498 19508
rect 14274 19456 14280 19508
rect 14332 19496 14338 19508
rect 14332 19468 14412 19496
rect 14332 19456 14338 19468
rect 10229 19431 10287 19437
rect 10229 19397 10241 19431
rect 10275 19428 10287 19431
rect 10318 19428 10324 19440
rect 10275 19400 10324 19428
rect 10275 19397 10287 19400
rect 10229 19391 10287 19397
rect 10318 19388 10324 19400
rect 10376 19388 10382 19440
rect 11977 19363 12035 19369
rect 8220 19332 8892 19360
rect 4433 19323 4491 19329
rect 4157 19295 4215 19301
rect 4157 19261 4169 19295
rect 4203 19292 4215 19295
rect 4246 19292 4252 19304
rect 4203 19264 4252 19292
rect 4203 19261 4215 19264
rect 4157 19255 4215 19261
rect 4246 19252 4252 19264
rect 4304 19292 4310 19304
rect 4798 19292 4804 19304
rect 4304 19264 4568 19292
rect 4759 19264 4804 19292
rect 4304 19252 4310 19264
rect 4540 19224 4568 19264
rect 4798 19252 4804 19264
rect 4856 19252 4862 19304
rect 5068 19295 5126 19301
rect 5068 19261 5080 19295
rect 5114 19292 5126 19295
rect 5350 19292 5356 19304
rect 5114 19264 5356 19292
rect 5114 19261 5126 19264
rect 5068 19255 5126 19261
rect 5350 19252 5356 19264
rect 5408 19252 5414 19304
rect 5626 19252 5632 19304
rect 5684 19292 5690 19304
rect 6546 19292 6552 19304
rect 5684 19264 6552 19292
rect 5684 19252 5690 19264
rect 6546 19252 6552 19264
rect 6604 19252 6610 19304
rect 7009 19295 7067 19301
rect 7009 19261 7021 19295
rect 7055 19292 7067 19295
rect 7098 19292 7104 19304
rect 7055 19264 7104 19292
rect 7055 19261 7067 19264
rect 7009 19255 7067 19261
rect 7098 19252 7104 19264
rect 7156 19252 7162 19304
rect 8662 19292 8668 19304
rect 7208 19264 8668 19292
rect 5442 19224 5448 19236
rect 3712 19196 4292 19224
rect 4540 19196 5448 19224
rect 1360 19128 2636 19156
rect 1360 19116 1366 19128
rect 2682 19116 2688 19168
rect 2740 19156 2746 19168
rect 4154 19156 4160 19168
rect 2740 19128 4160 19156
rect 2740 19116 2746 19128
rect 4154 19116 4160 19128
rect 4212 19116 4218 19168
rect 4264 19165 4292 19196
rect 5442 19184 5448 19196
rect 5500 19184 5506 19236
rect 5534 19184 5540 19236
rect 5592 19224 5598 19236
rect 7208 19224 7236 19264
rect 8662 19252 8668 19264
rect 8720 19252 8726 19304
rect 8864 19301 8892 19332
rect 11977 19329 11989 19363
rect 12023 19360 12035 19363
rect 12066 19360 12072 19372
rect 12023 19332 12072 19360
rect 12023 19329 12035 19332
rect 11977 19323 12035 19329
rect 12066 19320 12072 19332
rect 12124 19320 12130 19372
rect 13081 19363 13139 19369
rect 13081 19329 13093 19363
rect 13127 19360 13139 19363
rect 13722 19360 13728 19372
rect 13127 19332 13728 19360
rect 13127 19329 13139 19332
rect 13081 19323 13139 19329
rect 13722 19320 13728 19332
rect 13780 19320 13786 19372
rect 8849 19295 8907 19301
rect 8849 19261 8861 19295
rect 8895 19292 8907 19295
rect 8895 19264 8929 19292
rect 8895 19261 8907 19264
rect 8849 19255 8907 19261
rect 9674 19252 9680 19304
rect 9732 19292 9738 19304
rect 10505 19295 10563 19301
rect 10505 19292 10517 19295
rect 9732 19264 10517 19292
rect 9732 19252 9738 19264
rect 10505 19261 10517 19264
rect 10551 19261 10563 19295
rect 10505 19255 10563 19261
rect 11793 19295 11851 19301
rect 11793 19261 11805 19295
rect 11839 19292 11851 19295
rect 12434 19292 12440 19304
rect 11839 19264 12440 19292
rect 11839 19261 11851 19264
rect 11793 19255 11851 19261
rect 12434 19252 12440 19264
rect 12492 19252 12498 19304
rect 13446 19292 13452 19304
rect 13407 19264 13452 19292
rect 13446 19252 13452 19264
rect 13504 19252 13510 19304
rect 13998 19252 14004 19304
rect 14056 19292 14062 19304
rect 14384 19301 14412 19468
rect 17954 19456 17960 19508
rect 18012 19496 18018 19508
rect 18874 19496 18880 19508
rect 18012 19468 18880 19496
rect 18012 19456 18018 19468
rect 18874 19456 18880 19468
rect 18932 19456 18938 19508
rect 16868 19400 20484 19428
rect 16868 19369 16896 19400
rect 20456 19372 20484 19400
rect 16853 19363 16911 19369
rect 16853 19329 16865 19363
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 16942 19320 16948 19372
rect 17000 19360 17006 19372
rect 17402 19360 17408 19372
rect 17000 19332 17408 19360
rect 17000 19320 17006 19332
rect 17402 19320 17408 19332
rect 17460 19320 17466 19372
rect 20438 19320 20444 19372
rect 20496 19360 20502 19372
rect 20717 19363 20775 19369
rect 20717 19360 20729 19363
rect 20496 19332 20729 19360
rect 20496 19320 20502 19332
rect 20717 19329 20729 19332
rect 20763 19329 20775 19363
rect 20717 19323 20775 19329
rect 14358 19295 14416 19301
rect 14056 19264 14320 19292
rect 14056 19252 14062 19264
rect 5592 19196 7236 19224
rect 7276 19227 7334 19233
rect 5592 19184 5598 19196
rect 7276 19193 7288 19227
rect 7322 19224 7334 19227
rect 7742 19224 7748 19236
rect 7322 19196 7748 19224
rect 7322 19193 7334 19196
rect 7276 19187 7334 19193
rect 7742 19184 7748 19196
rect 7800 19184 7806 19236
rect 8294 19184 8300 19236
rect 8352 19184 8358 19236
rect 9116 19227 9174 19233
rect 9116 19193 9128 19227
rect 9162 19224 9174 19227
rect 9582 19224 9588 19236
rect 9162 19196 9588 19224
rect 9162 19193 9174 19196
rect 9116 19187 9174 19193
rect 9582 19184 9588 19196
rect 9640 19184 9646 19236
rect 9950 19184 9956 19236
rect 10008 19224 10014 19236
rect 10781 19227 10839 19233
rect 10781 19224 10793 19227
rect 10008 19196 10793 19224
rect 10008 19184 10014 19196
rect 10781 19193 10793 19196
rect 10827 19193 10839 19227
rect 11882 19224 11888 19236
rect 10781 19187 10839 19193
rect 11348 19196 11888 19224
rect 4249 19159 4307 19165
rect 4249 19125 4261 19159
rect 4295 19156 4307 19159
rect 4890 19156 4896 19168
rect 4295 19128 4896 19156
rect 4295 19125 4307 19128
rect 4249 19119 4307 19125
rect 4890 19116 4896 19128
rect 4948 19116 4954 19168
rect 5810 19116 5816 19168
rect 5868 19156 5874 19168
rect 6181 19159 6239 19165
rect 6181 19156 6193 19159
rect 5868 19128 6193 19156
rect 5868 19116 5874 19128
rect 6181 19125 6193 19128
rect 6227 19125 6239 19159
rect 6181 19119 6239 19125
rect 6362 19116 6368 19168
rect 6420 19156 6426 19168
rect 8312 19156 8340 19184
rect 6420 19128 8340 19156
rect 6420 19116 6426 19128
rect 8386 19116 8392 19168
rect 8444 19156 8450 19168
rect 10042 19156 10048 19168
rect 8444 19128 10048 19156
rect 8444 19116 8450 19128
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 10318 19116 10324 19168
rect 10376 19156 10382 19168
rect 10502 19156 10508 19168
rect 10376 19128 10508 19156
rect 10376 19116 10382 19128
rect 10502 19116 10508 19128
rect 10560 19116 10566 19168
rect 11348 19165 11376 19196
rect 11882 19184 11888 19196
rect 11940 19184 11946 19236
rect 12805 19227 12863 19233
rect 12805 19224 12817 19227
rect 11992 19196 12817 19224
rect 11333 19159 11391 19165
rect 11333 19125 11345 19159
rect 11379 19125 11391 19159
rect 11698 19156 11704 19168
rect 11659 19128 11704 19156
rect 11333 19119 11391 19125
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 11790 19116 11796 19168
rect 11848 19156 11854 19168
rect 11992 19156 12020 19196
rect 12805 19193 12817 19196
rect 12851 19193 12863 19227
rect 12805 19187 12863 19193
rect 13078 19184 13084 19236
rect 13136 19224 13142 19236
rect 14292 19224 14320 19264
rect 14358 19261 14370 19295
rect 14404 19261 14416 19295
rect 15105 19295 15163 19301
rect 15105 19292 15117 19295
rect 14358 19255 14416 19261
rect 14568 19264 15117 19292
rect 14568 19224 14596 19264
rect 15105 19261 15117 19264
rect 15151 19261 15163 19295
rect 15105 19255 15163 19261
rect 15657 19295 15715 19301
rect 15657 19261 15669 19295
rect 15703 19261 15715 19295
rect 15657 19255 15715 19261
rect 16117 19295 16175 19301
rect 16117 19261 16129 19295
rect 16163 19292 16175 19295
rect 16163 19264 16988 19292
rect 16163 19261 16175 19264
rect 16117 19255 16175 19261
rect 13136 19196 14228 19224
rect 14292 19196 14596 19224
rect 14645 19227 14703 19233
rect 13136 19184 13142 19196
rect 11848 19128 12020 19156
rect 11848 19116 11854 19128
rect 12158 19116 12164 19168
rect 12216 19156 12222 19168
rect 12897 19159 12955 19165
rect 12897 19156 12909 19159
rect 12216 19128 12909 19156
rect 12216 19116 12222 19128
rect 12897 19125 12909 19128
rect 12943 19125 12955 19159
rect 12897 19119 12955 19125
rect 13633 19159 13691 19165
rect 13633 19125 13645 19159
rect 13679 19156 13691 19159
rect 13814 19156 13820 19168
rect 13679 19128 13820 19156
rect 13679 19125 13691 19128
rect 13633 19119 13691 19125
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 14200 19156 14228 19196
rect 14645 19193 14657 19227
rect 14691 19224 14703 19227
rect 15672 19224 15700 19255
rect 16850 19224 16856 19236
rect 14691 19196 15700 19224
rect 15856 19196 16856 19224
rect 14691 19193 14703 19196
rect 14645 19187 14703 19193
rect 15856 19165 15884 19196
rect 16850 19184 16856 19196
rect 16908 19184 16914 19236
rect 16960 19224 16988 19264
rect 17034 19252 17040 19304
rect 17092 19292 17098 19304
rect 17221 19295 17279 19301
rect 17221 19292 17233 19295
rect 17092 19264 17233 19292
rect 17092 19252 17098 19264
rect 17221 19261 17233 19264
rect 17267 19261 17279 19295
rect 17494 19292 17500 19304
rect 17455 19264 17500 19292
rect 17221 19255 17279 19261
rect 17494 19252 17500 19264
rect 17552 19252 17558 19304
rect 18049 19295 18107 19301
rect 18049 19261 18061 19295
rect 18095 19292 18107 19295
rect 18690 19292 18696 19304
rect 18095 19264 18696 19292
rect 18095 19261 18107 19264
rect 18049 19255 18107 19261
rect 18690 19252 18696 19264
rect 18748 19252 18754 19304
rect 18785 19295 18843 19301
rect 18785 19261 18797 19295
rect 18831 19292 18843 19295
rect 19794 19292 19800 19304
rect 18831 19264 19800 19292
rect 18831 19261 18843 19264
rect 18785 19255 18843 19261
rect 19794 19252 19800 19264
rect 19852 19252 19858 19304
rect 17770 19224 17776 19236
rect 16960 19196 17776 19224
rect 17770 19184 17776 19196
rect 17828 19184 17834 19236
rect 18138 19184 18144 19236
rect 18196 19224 18202 19236
rect 19429 19227 19487 19233
rect 19429 19224 19441 19227
rect 18196 19196 19441 19224
rect 18196 19184 18202 19196
rect 19429 19193 19441 19196
rect 19475 19193 19487 19227
rect 19429 19187 19487 19193
rect 19610 19184 19616 19236
rect 19668 19224 19674 19236
rect 20625 19227 20683 19233
rect 20625 19224 20637 19227
rect 19668 19196 20637 19224
rect 19668 19184 19674 19196
rect 20625 19193 20637 19196
rect 20671 19193 20683 19227
rect 20625 19187 20683 19193
rect 15289 19159 15347 19165
rect 15289 19156 15301 19159
rect 14200 19128 15301 19156
rect 15289 19125 15301 19128
rect 15335 19125 15347 19159
rect 15289 19119 15347 19125
rect 15841 19159 15899 19165
rect 15841 19125 15853 19159
rect 15887 19125 15899 19159
rect 15841 19119 15899 19125
rect 16117 19159 16175 19165
rect 16117 19125 16129 19159
rect 16163 19156 16175 19159
rect 16209 19159 16267 19165
rect 16209 19156 16221 19159
rect 16163 19128 16221 19156
rect 16163 19125 16175 19128
rect 16117 19119 16175 19125
rect 16209 19125 16221 19128
rect 16255 19125 16267 19159
rect 16209 19119 16267 19125
rect 16390 19116 16396 19168
rect 16448 19156 16454 19168
rect 16577 19159 16635 19165
rect 16577 19156 16589 19159
rect 16448 19128 16589 19156
rect 16448 19116 16454 19128
rect 16577 19125 16589 19128
rect 16623 19125 16635 19159
rect 16577 19119 16635 19125
rect 16669 19159 16727 19165
rect 16669 19125 16681 19159
rect 16715 19156 16727 19159
rect 17862 19156 17868 19168
rect 16715 19128 17868 19156
rect 16715 19125 16727 19128
rect 16669 19119 16727 19125
rect 17862 19116 17868 19128
rect 17920 19116 17926 19168
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 18874 19156 18880 19168
rect 18279 19128 18880 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 18874 19116 18880 19128
rect 18932 19116 18938 19168
rect 20162 19156 20168 19168
rect 20123 19128 20168 19156
rect 20162 19116 20168 19128
rect 20220 19116 20226 19168
rect 20530 19156 20536 19168
rect 20491 19128 20536 19156
rect 20530 19116 20536 19128
rect 20588 19116 20594 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 2314 18952 2320 18964
rect 2275 18924 2320 18952
rect 2314 18912 2320 18924
rect 2372 18912 2378 18964
rect 2961 18955 3019 18961
rect 2961 18921 2973 18955
rect 3007 18952 3019 18955
rect 3234 18952 3240 18964
rect 3007 18924 3240 18952
rect 3007 18921 3019 18924
rect 2961 18915 3019 18921
rect 3234 18912 3240 18924
rect 3292 18912 3298 18964
rect 3329 18955 3387 18961
rect 3329 18921 3341 18955
rect 3375 18952 3387 18955
rect 5074 18952 5080 18964
rect 3375 18924 5080 18952
rect 3375 18921 3387 18924
rect 3329 18915 3387 18921
rect 5074 18912 5080 18924
rect 5132 18912 5138 18964
rect 6178 18952 6184 18964
rect 6139 18924 6184 18952
rect 6178 18912 6184 18924
rect 6236 18912 6242 18964
rect 6917 18955 6975 18961
rect 6917 18921 6929 18955
rect 6963 18952 6975 18955
rect 9490 18952 9496 18964
rect 6963 18924 9496 18952
rect 6963 18921 6975 18924
rect 6917 18915 6975 18921
rect 9490 18912 9496 18924
rect 9548 18912 9554 18964
rect 9677 18955 9735 18961
rect 9677 18921 9689 18955
rect 9723 18952 9735 18955
rect 9723 18924 9996 18952
rect 9723 18921 9735 18924
rect 9677 18915 9735 18921
rect 566 18844 572 18896
rect 624 18884 630 18896
rect 2682 18884 2688 18896
rect 624 18856 2688 18884
rect 624 18844 630 18856
rect 2682 18844 2688 18856
rect 2740 18844 2746 18896
rect 4798 18884 4804 18896
rect 4080 18856 4804 18884
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 2130 18816 2136 18828
rect 1443 18788 2136 18816
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 2130 18776 2136 18788
rect 2188 18776 2194 18828
rect 4080 18825 4108 18856
rect 4798 18844 4804 18856
rect 4856 18844 4862 18896
rect 4890 18844 4896 18896
rect 4948 18884 4954 18896
rect 8386 18884 8392 18896
rect 4948 18856 8392 18884
rect 4948 18844 4954 18856
rect 8386 18844 8392 18856
rect 8444 18844 8450 18896
rect 9582 18844 9588 18896
rect 9640 18884 9646 18896
rect 9968 18884 9996 18924
rect 10042 18912 10048 18964
rect 10100 18952 10106 18964
rect 12158 18952 12164 18964
rect 10100 18924 12164 18952
rect 10100 18912 10106 18924
rect 12158 18912 12164 18924
rect 12216 18912 12222 18964
rect 14366 18912 14372 18964
rect 14424 18952 14430 18964
rect 17218 18952 17224 18964
rect 14424 18924 17224 18952
rect 14424 18912 14430 18924
rect 17218 18912 17224 18924
rect 17276 18912 17282 18964
rect 17310 18912 17316 18964
rect 17368 18952 17374 18964
rect 17681 18955 17739 18961
rect 17681 18952 17693 18955
rect 17368 18924 17693 18952
rect 17368 18912 17374 18924
rect 17681 18921 17693 18924
rect 17727 18921 17739 18955
rect 17681 18915 17739 18921
rect 19245 18955 19303 18961
rect 19245 18921 19257 18955
rect 19291 18952 19303 18955
rect 19797 18955 19855 18961
rect 19797 18952 19809 18955
rect 19291 18924 19809 18952
rect 19291 18921 19303 18924
rect 19245 18915 19303 18921
rect 19797 18921 19809 18924
rect 19843 18921 19855 18955
rect 19797 18915 19855 18921
rect 10226 18884 10232 18896
rect 9640 18856 9720 18884
rect 9968 18856 10232 18884
rect 9640 18844 9646 18856
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18785 4123 18819
rect 4065 18779 4123 18785
rect 4332 18819 4390 18825
rect 4332 18785 4344 18819
rect 4378 18816 4390 18819
rect 4706 18816 4712 18828
rect 4378 18788 4712 18816
rect 4378 18785 4390 18788
rect 4332 18779 4390 18785
rect 4706 18776 4712 18788
rect 4764 18776 4770 18828
rect 6089 18819 6147 18825
rect 6089 18785 6101 18819
rect 6135 18816 6147 18819
rect 6362 18816 6368 18828
rect 6135 18788 6368 18816
rect 6135 18785 6147 18788
rect 6089 18779 6147 18785
rect 6362 18776 6368 18788
rect 6420 18776 6426 18828
rect 6730 18816 6736 18828
rect 6691 18788 6736 18816
rect 6730 18776 6736 18788
rect 6788 18776 6794 18828
rect 7098 18776 7104 18828
rect 7156 18816 7162 18828
rect 7377 18819 7435 18825
rect 7377 18816 7389 18819
rect 7156 18788 7389 18816
rect 7156 18776 7162 18788
rect 7377 18785 7389 18788
rect 7423 18785 7435 18819
rect 7377 18779 7435 18785
rect 7644 18819 7702 18825
rect 7644 18785 7656 18819
rect 7690 18816 7702 18819
rect 7690 18788 8616 18816
rect 7690 18785 7702 18788
rect 7644 18779 7702 18785
rect 2038 18708 2044 18760
rect 2096 18748 2102 18760
rect 2406 18748 2412 18760
rect 2096 18720 2412 18748
rect 2096 18708 2102 18720
rect 2406 18708 2412 18720
rect 2464 18708 2470 18760
rect 2593 18751 2651 18757
rect 2593 18717 2605 18751
rect 2639 18748 2651 18751
rect 2682 18748 2688 18760
rect 2639 18720 2688 18748
rect 2639 18717 2651 18720
rect 2593 18711 2651 18717
rect 2682 18708 2688 18720
rect 2740 18708 2746 18760
rect 3418 18748 3424 18760
rect 3379 18720 3424 18748
rect 3418 18708 3424 18720
rect 3476 18708 3482 18760
rect 3605 18751 3663 18757
rect 3605 18717 3617 18751
rect 3651 18717 3663 18751
rect 3605 18711 3663 18717
rect 1578 18612 1584 18624
rect 1539 18584 1584 18612
rect 1578 18572 1584 18584
rect 1636 18572 1642 18624
rect 1949 18615 2007 18621
rect 1949 18581 1961 18615
rect 1995 18612 2007 18615
rect 2866 18612 2872 18624
rect 1995 18584 2872 18612
rect 1995 18581 2007 18584
rect 1949 18575 2007 18581
rect 2866 18572 2872 18584
rect 2924 18572 2930 18624
rect 3620 18612 3648 18711
rect 5810 18708 5816 18760
rect 5868 18748 5874 18760
rect 6273 18751 6331 18757
rect 6273 18748 6285 18751
rect 5868 18720 6285 18748
rect 5868 18708 5874 18720
rect 6273 18717 6285 18720
rect 6319 18717 6331 18751
rect 8588 18748 8616 18788
rect 8662 18776 8668 18828
rect 8720 18816 8726 18828
rect 9033 18819 9091 18825
rect 9033 18816 9045 18819
rect 8720 18788 9045 18816
rect 8720 18776 8726 18788
rect 9033 18785 9045 18788
rect 9079 18785 9091 18819
rect 9692 18816 9720 18856
rect 10226 18844 10232 18856
rect 10284 18844 10290 18896
rect 12710 18884 12716 18896
rect 10704 18856 12716 18884
rect 9692 18788 9812 18816
rect 9033 18779 9091 18785
rect 9122 18748 9128 18760
rect 8588 18720 9128 18748
rect 6273 18711 6331 18717
rect 9122 18708 9128 18720
rect 9180 18708 9186 18760
rect 9784 18748 9812 18788
rect 9858 18776 9864 18828
rect 9916 18816 9922 18828
rect 9950 18816 9956 18828
rect 9916 18788 9956 18816
rect 9916 18776 9922 18788
rect 9950 18776 9956 18788
rect 10008 18776 10014 18828
rect 10704 18825 10732 18856
rect 12710 18844 12716 18856
rect 12768 18844 12774 18896
rect 12897 18887 12955 18893
rect 12897 18853 12909 18887
rect 12943 18884 12955 18887
rect 13078 18884 13084 18896
rect 12943 18856 13084 18884
rect 12943 18853 12955 18856
rect 12897 18847 12955 18853
rect 13078 18844 13084 18856
rect 13136 18884 13142 18896
rect 13326 18887 13384 18893
rect 13326 18884 13338 18887
rect 13136 18856 13338 18884
rect 13136 18844 13142 18856
rect 13326 18853 13338 18856
rect 13372 18853 13384 18887
rect 13326 18847 13384 18853
rect 13538 18844 13544 18896
rect 13596 18884 13602 18896
rect 15470 18884 15476 18896
rect 13596 18856 15476 18884
rect 13596 18844 13602 18856
rect 15470 18844 15476 18856
rect 15528 18844 15534 18896
rect 15749 18887 15807 18893
rect 15749 18853 15761 18887
rect 15795 18884 15807 18887
rect 17586 18884 17592 18896
rect 15795 18856 17592 18884
rect 15795 18853 15807 18856
rect 15749 18847 15807 18853
rect 17586 18844 17592 18856
rect 17644 18844 17650 18896
rect 18325 18887 18383 18893
rect 18325 18853 18337 18887
rect 18371 18884 18383 18887
rect 18782 18884 18788 18896
rect 18371 18856 18788 18884
rect 18371 18853 18383 18856
rect 18325 18847 18383 18853
rect 18782 18844 18788 18856
rect 18840 18844 18846 18896
rect 19334 18844 19340 18896
rect 19392 18884 19398 18896
rect 20165 18887 20223 18893
rect 20165 18884 20177 18887
rect 19392 18856 20177 18884
rect 19392 18844 19398 18856
rect 20165 18853 20177 18856
rect 20211 18853 20223 18887
rect 20165 18847 20223 18853
rect 10137 18819 10195 18825
rect 10137 18785 10149 18819
rect 10183 18816 10195 18819
rect 10689 18819 10747 18825
rect 10183 18788 10364 18816
rect 10183 18785 10195 18788
rect 10137 18779 10195 18785
rect 10229 18751 10287 18757
rect 10229 18748 10241 18751
rect 9784 18720 10241 18748
rect 10229 18717 10241 18720
rect 10275 18717 10287 18751
rect 10336 18748 10364 18788
rect 10689 18785 10701 18819
rect 10735 18785 10747 18819
rect 10689 18779 10747 18785
rect 11692 18819 11750 18825
rect 11692 18785 11704 18819
rect 11738 18816 11750 18819
rect 12066 18816 12072 18828
rect 11738 18788 12072 18816
rect 11738 18785 11750 18788
rect 11692 18779 11750 18785
rect 12066 18776 12072 18788
rect 12124 18776 12130 18828
rect 13630 18816 13636 18828
rect 13096 18788 13636 18816
rect 10778 18748 10784 18760
rect 10336 18720 10784 18748
rect 10229 18711 10287 18717
rect 10778 18708 10784 18720
rect 10836 18708 10842 18760
rect 10965 18751 11023 18757
rect 10965 18717 10977 18751
rect 11011 18748 11023 18751
rect 11146 18748 11152 18760
rect 11011 18720 11152 18748
rect 11011 18717 11023 18720
rect 10965 18711 11023 18717
rect 11146 18708 11152 18720
rect 11204 18708 11210 18760
rect 13096 18757 13124 18788
rect 13630 18776 13636 18788
rect 13688 18776 13694 18828
rect 13814 18776 13820 18828
rect 13872 18816 13878 18828
rect 15286 18816 15292 18828
rect 13872 18788 15292 18816
rect 13872 18776 13878 18788
rect 15286 18776 15292 18788
rect 15344 18776 15350 18828
rect 16114 18825 16120 18828
rect 16108 18816 16120 18825
rect 16027 18788 16120 18816
rect 16108 18779 16120 18788
rect 16172 18816 16178 18828
rect 16942 18816 16948 18828
rect 16172 18788 16948 18816
rect 16114 18776 16120 18779
rect 16172 18776 16178 18788
rect 16942 18776 16948 18788
rect 17000 18776 17006 18828
rect 17494 18816 17500 18828
rect 17455 18788 17500 18816
rect 17494 18776 17500 18788
rect 17552 18776 17558 18828
rect 18049 18819 18107 18825
rect 18049 18785 18061 18819
rect 18095 18816 18107 18819
rect 18966 18816 18972 18828
rect 18095 18788 18972 18816
rect 18095 18785 18107 18788
rect 18049 18779 18107 18785
rect 11425 18751 11483 18757
rect 11425 18717 11437 18751
rect 11471 18717 11483 18751
rect 11425 18711 11483 18717
rect 13081 18751 13139 18757
rect 13081 18717 13093 18751
rect 13127 18717 13139 18751
rect 13081 18711 13139 18717
rect 10502 18640 10508 18692
rect 10560 18680 10566 18692
rect 11440 18680 11468 18711
rect 15470 18708 15476 18760
rect 15528 18748 15534 18760
rect 15841 18751 15899 18757
rect 15841 18748 15853 18751
rect 15528 18720 15853 18748
rect 15528 18708 15534 18720
rect 15841 18717 15853 18720
rect 15887 18717 15899 18751
rect 15841 18711 15899 18717
rect 17034 18708 17040 18760
rect 17092 18748 17098 18760
rect 18064 18748 18092 18779
rect 18966 18776 18972 18788
rect 19024 18776 19030 18828
rect 19150 18816 19156 18828
rect 19111 18788 19156 18816
rect 19150 18776 19156 18788
rect 19208 18776 19214 18828
rect 17092 18720 18092 18748
rect 17092 18708 17098 18720
rect 18782 18708 18788 18760
rect 18840 18748 18846 18760
rect 19337 18751 19395 18757
rect 19337 18748 19349 18751
rect 18840 18720 19349 18748
rect 18840 18708 18846 18720
rect 19337 18717 19349 18720
rect 19383 18717 19395 18751
rect 19337 18711 19395 18717
rect 19794 18708 19800 18760
rect 19852 18748 19858 18760
rect 20257 18751 20315 18757
rect 20257 18748 20269 18751
rect 19852 18720 20269 18748
rect 19852 18708 19858 18720
rect 20257 18717 20269 18720
rect 20303 18717 20315 18751
rect 20438 18748 20444 18760
rect 20399 18720 20444 18748
rect 20257 18711 20315 18717
rect 20438 18708 20444 18720
rect 20496 18708 20502 18760
rect 10560 18652 11468 18680
rect 12805 18683 12863 18689
rect 10560 18640 10566 18652
rect 12805 18649 12817 18683
rect 12851 18680 12863 18683
rect 12897 18683 12955 18689
rect 12897 18680 12909 18683
rect 12851 18652 12909 18680
rect 12851 18649 12863 18652
rect 12805 18643 12863 18649
rect 12897 18649 12909 18652
rect 12943 18649 12955 18683
rect 12897 18643 12955 18649
rect 14274 18640 14280 18692
rect 14332 18680 14338 18692
rect 14332 18652 15884 18680
rect 14332 18640 14338 18652
rect 5350 18612 5356 18624
rect 3620 18584 5356 18612
rect 5350 18572 5356 18584
rect 5408 18612 5414 18624
rect 5445 18615 5503 18621
rect 5445 18612 5457 18615
rect 5408 18584 5457 18612
rect 5408 18572 5414 18584
rect 5445 18581 5457 18584
rect 5491 18581 5503 18615
rect 5718 18612 5724 18624
rect 5679 18584 5724 18612
rect 5445 18575 5503 18581
rect 5718 18572 5724 18584
rect 5776 18572 5782 18624
rect 5902 18572 5908 18624
rect 5960 18612 5966 18624
rect 7374 18612 7380 18624
rect 5960 18584 7380 18612
rect 5960 18572 5966 18584
rect 7374 18572 7380 18584
rect 7432 18572 7438 18624
rect 8018 18572 8024 18624
rect 8076 18612 8082 18624
rect 8757 18615 8815 18621
rect 8757 18612 8769 18615
rect 8076 18584 8769 18612
rect 8076 18572 8082 18584
rect 8757 18581 8769 18584
rect 8803 18581 8815 18615
rect 8757 18575 8815 18581
rect 9217 18615 9275 18621
rect 9217 18581 9229 18615
rect 9263 18612 9275 18615
rect 11606 18612 11612 18624
rect 9263 18584 11612 18612
rect 9263 18581 9275 18584
rect 9217 18575 9275 18581
rect 11606 18572 11612 18584
rect 11664 18572 11670 18624
rect 11698 18572 11704 18624
rect 11756 18612 11762 18624
rect 14090 18612 14096 18624
rect 11756 18584 14096 18612
rect 11756 18572 11762 18584
rect 14090 18572 14096 18584
rect 14148 18572 14154 18624
rect 14182 18572 14188 18624
rect 14240 18612 14246 18624
rect 14461 18615 14519 18621
rect 14461 18612 14473 18615
rect 14240 18584 14473 18612
rect 14240 18572 14246 18584
rect 14461 18581 14473 18584
rect 14507 18581 14519 18615
rect 14461 18575 14519 18581
rect 15473 18615 15531 18621
rect 15473 18581 15485 18615
rect 15519 18612 15531 18615
rect 15749 18615 15807 18621
rect 15749 18612 15761 18615
rect 15519 18584 15761 18612
rect 15519 18581 15531 18584
rect 15473 18575 15531 18581
rect 15749 18581 15761 18584
rect 15795 18581 15807 18615
rect 15856 18612 15884 18652
rect 16850 18640 16856 18692
rect 16908 18680 16914 18692
rect 20530 18680 20536 18692
rect 16908 18652 20536 18680
rect 16908 18640 16914 18652
rect 20530 18640 20536 18652
rect 20588 18640 20594 18692
rect 16758 18612 16764 18624
rect 15856 18584 16764 18612
rect 15749 18575 15807 18581
rect 16758 18572 16764 18584
rect 16816 18572 16822 18624
rect 17218 18612 17224 18624
rect 17179 18584 17224 18612
rect 17218 18572 17224 18584
rect 17276 18572 17282 18624
rect 18785 18615 18843 18621
rect 18785 18581 18797 18615
rect 18831 18612 18843 18615
rect 18966 18612 18972 18624
rect 18831 18584 18972 18612
rect 18831 18581 18843 18584
rect 18785 18575 18843 18581
rect 18966 18572 18972 18584
rect 19024 18572 19030 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 2406 18368 2412 18420
rect 2464 18408 2470 18420
rect 4798 18408 4804 18420
rect 2464 18380 4804 18408
rect 2464 18368 2470 18380
rect 4798 18368 4804 18380
rect 4856 18368 4862 18420
rect 4893 18411 4951 18417
rect 4893 18377 4905 18411
rect 4939 18408 4951 18411
rect 5718 18408 5724 18420
rect 4939 18380 5724 18408
rect 4939 18377 4951 18380
rect 4893 18371 4951 18377
rect 5718 18368 5724 18380
rect 5776 18368 5782 18420
rect 7466 18408 7472 18420
rect 7427 18380 7472 18408
rect 7466 18368 7472 18380
rect 7524 18368 7530 18420
rect 8481 18411 8539 18417
rect 8481 18377 8493 18411
rect 8527 18408 8539 18411
rect 9030 18408 9036 18420
rect 8527 18380 9036 18408
rect 8527 18377 8539 18380
rect 8481 18371 8539 18377
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 9493 18411 9551 18417
rect 9493 18377 9505 18411
rect 9539 18408 9551 18411
rect 10134 18408 10140 18420
rect 9539 18380 10140 18408
rect 9539 18377 9551 18380
rect 9493 18371 9551 18377
rect 10134 18368 10140 18380
rect 10192 18368 10198 18420
rect 12066 18408 12072 18420
rect 12027 18380 12072 18408
rect 12066 18368 12072 18380
rect 12124 18368 12130 18420
rect 12437 18411 12495 18417
rect 12437 18377 12449 18411
rect 12483 18408 12495 18411
rect 12618 18408 12624 18420
rect 12483 18380 12624 18408
rect 12483 18377 12495 18380
rect 12437 18371 12495 18377
rect 12618 18368 12624 18380
rect 12676 18368 12682 18420
rect 12710 18368 12716 18420
rect 12768 18408 12774 18420
rect 13262 18408 13268 18420
rect 12768 18380 13268 18408
rect 12768 18368 12774 18380
rect 13262 18368 13268 18380
rect 13320 18368 13326 18420
rect 14090 18368 14096 18420
rect 14148 18408 14154 18420
rect 15749 18411 15807 18417
rect 15749 18408 15761 18411
rect 14148 18380 15761 18408
rect 14148 18368 14154 18380
rect 15749 18377 15761 18380
rect 15795 18377 15807 18411
rect 17218 18408 17224 18420
rect 15749 18371 15807 18377
rect 16960 18380 17224 18408
rect 7101 18343 7159 18349
rect 3436 18312 4936 18340
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18204 1823 18207
rect 1946 18204 1952 18216
rect 1811 18176 1952 18204
rect 1811 18173 1823 18176
rect 1765 18167 1823 18173
rect 1946 18164 1952 18176
rect 2004 18164 2010 18216
rect 2038 18164 2044 18216
rect 2096 18204 2102 18216
rect 2409 18207 2467 18213
rect 2409 18204 2421 18207
rect 2096 18176 2421 18204
rect 2096 18164 2102 18176
rect 2409 18173 2421 18176
rect 2455 18173 2467 18207
rect 2409 18167 2467 18173
rect 3050 18164 3056 18216
rect 3108 18204 3114 18216
rect 3436 18204 3464 18312
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18272 4767 18275
rect 4798 18272 4804 18284
rect 4755 18244 4804 18272
rect 4755 18241 4767 18244
rect 4709 18235 4767 18241
rect 4798 18232 4804 18244
rect 4856 18232 4862 18284
rect 4908 18272 4936 18312
rect 7101 18309 7113 18343
rect 7147 18340 7159 18343
rect 7282 18340 7288 18352
rect 7147 18312 7288 18340
rect 7147 18309 7159 18312
rect 7101 18303 7159 18309
rect 7282 18300 7288 18312
rect 7340 18300 7346 18352
rect 7742 18300 7748 18352
rect 7800 18340 7806 18352
rect 7800 18312 10180 18340
rect 7800 18300 7806 18312
rect 4908 18244 5212 18272
rect 3108 18176 3464 18204
rect 3108 18164 3114 18176
rect 3786 18164 3792 18216
rect 3844 18204 3850 18216
rect 4433 18207 4491 18213
rect 4433 18204 4445 18207
rect 3844 18176 4445 18204
rect 3844 18164 3850 18176
rect 4433 18173 4445 18176
rect 4479 18173 4491 18207
rect 4433 18167 4491 18173
rect 4525 18207 4583 18213
rect 4525 18173 4537 18207
rect 4571 18204 4583 18207
rect 4893 18207 4951 18213
rect 4893 18204 4905 18207
rect 4571 18176 4905 18204
rect 4571 18173 4583 18176
rect 4525 18167 4583 18173
rect 4893 18173 4905 18176
rect 4939 18173 4951 18207
rect 4893 18167 4951 18173
rect 5077 18207 5135 18213
rect 5077 18173 5089 18207
rect 5123 18173 5135 18207
rect 5184 18204 5212 18244
rect 6270 18232 6276 18284
rect 6328 18272 6334 18284
rect 7558 18272 7564 18284
rect 6328 18244 7564 18272
rect 6328 18232 6334 18244
rect 7558 18232 7564 18244
rect 7616 18232 7622 18284
rect 7929 18275 7987 18281
rect 7929 18241 7941 18275
rect 7975 18272 7987 18275
rect 7975 18244 8064 18272
rect 7975 18241 7987 18244
rect 7929 18235 7987 18241
rect 6914 18204 6920 18216
rect 5184 18176 5488 18204
rect 6875 18176 6920 18204
rect 5077 18167 5135 18173
rect 2676 18139 2734 18145
rect 2676 18105 2688 18139
rect 2722 18136 2734 18139
rect 2958 18136 2964 18148
rect 2722 18108 2964 18136
rect 2722 18105 2734 18108
rect 2676 18099 2734 18105
rect 2958 18096 2964 18108
rect 3016 18096 3022 18148
rect 2774 18028 2780 18080
rect 2832 18068 2838 18080
rect 3068 18068 3096 18164
rect 4706 18136 4712 18148
rect 3804 18108 4712 18136
rect 3804 18077 3832 18108
rect 4706 18096 4712 18108
rect 4764 18096 4770 18148
rect 5092 18136 5120 18167
rect 5341 18136 5347 18148
rect 4908 18108 5120 18136
rect 5302 18108 5347 18136
rect 4908 18080 4936 18108
rect 5341 18096 5347 18108
rect 5399 18096 5405 18148
rect 5460 18136 5488 18176
rect 6914 18164 6920 18176
rect 6972 18164 6978 18216
rect 7837 18207 7895 18213
rect 7837 18173 7849 18207
rect 7883 18204 7895 18207
rect 8036 18204 8064 18244
rect 8110 18232 8116 18284
rect 8168 18272 8174 18284
rect 9033 18275 9091 18281
rect 9033 18272 9045 18275
rect 8168 18244 9045 18272
rect 8168 18232 8174 18244
rect 9033 18241 9045 18244
rect 9079 18241 9091 18275
rect 9033 18235 9091 18241
rect 9582 18232 9588 18284
rect 9640 18272 9646 18284
rect 10045 18275 10103 18281
rect 10045 18272 10057 18275
rect 9640 18244 10057 18272
rect 9640 18232 9646 18244
rect 10045 18241 10057 18244
rect 10091 18241 10103 18275
rect 10045 18235 10103 18241
rect 8941 18207 8999 18213
rect 7883 18176 7972 18204
rect 8036 18176 8800 18204
rect 7883 18173 7895 18176
rect 7837 18167 7895 18173
rect 5460 18108 6960 18136
rect 2832 18040 3096 18068
rect 3789 18071 3847 18077
rect 2832 18028 2838 18040
rect 3789 18037 3801 18071
rect 3835 18037 3847 18071
rect 3789 18031 3847 18037
rect 4065 18071 4123 18077
rect 4065 18037 4077 18071
rect 4111 18068 4123 18071
rect 4338 18068 4344 18080
rect 4111 18040 4344 18068
rect 4111 18037 4123 18040
rect 4065 18031 4123 18037
rect 4338 18028 4344 18040
rect 4396 18028 4402 18080
rect 4890 18028 4896 18080
rect 4948 18028 4954 18080
rect 5442 18028 5448 18080
rect 5500 18068 5506 18080
rect 5810 18068 5816 18080
rect 5500 18040 5816 18068
rect 5500 18028 5506 18040
rect 5810 18028 5816 18040
rect 5868 18028 5874 18080
rect 6270 18028 6276 18080
rect 6328 18068 6334 18080
rect 6457 18071 6515 18077
rect 6457 18068 6469 18071
rect 6328 18040 6469 18068
rect 6328 18028 6334 18040
rect 6457 18037 6469 18040
rect 6503 18068 6515 18071
rect 6822 18068 6828 18080
rect 6503 18040 6828 18068
rect 6503 18037 6515 18040
rect 6457 18031 6515 18037
rect 6822 18028 6828 18040
rect 6880 18028 6886 18080
rect 6932 18068 6960 18108
rect 7098 18096 7104 18148
rect 7156 18136 7162 18148
rect 7742 18136 7748 18148
rect 7156 18108 7748 18136
rect 7156 18096 7162 18108
rect 7742 18096 7748 18108
rect 7800 18096 7806 18148
rect 7944 18136 7972 18176
rect 8570 18136 8576 18148
rect 7944 18108 8576 18136
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 8772 18136 8800 18176
rect 8941 18173 8953 18207
rect 8987 18204 8999 18207
rect 9398 18204 9404 18216
rect 8987 18176 9404 18204
rect 8987 18173 8999 18176
rect 8941 18167 8999 18173
rect 9398 18164 9404 18176
rect 9456 18164 9462 18216
rect 9953 18207 10011 18213
rect 9953 18173 9965 18207
rect 9999 18204 10011 18207
rect 10152 18204 10180 18312
rect 11882 18300 11888 18352
rect 11940 18340 11946 18352
rect 13449 18343 13507 18349
rect 11940 18312 12940 18340
rect 11940 18300 11946 18312
rect 10410 18232 10416 18284
rect 10468 18272 10474 18284
rect 10468 18244 10815 18272
rect 10468 18232 10474 18244
rect 10318 18204 10324 18216
rect 9999 18176 10324 18204
rect 9999 18173 10011 18176
rect 9953 18167 10011 18173
rect 10318 18164 10324 18176
rect 10376 18164 10382 18216
rect 10502 18164 10508 18216
rect 10560 18204 10566 18216
rect 10689 18207 10747 18213
rect 10689 18204 10701 18207
rect 10560 18176 10701 18204
rect 10560 18164 10566 18176
rect 10689 18173 10701 18176
rect 10735 18173 10747 18207
rect 10787 18204 10815 18244
rect 12250 18232 12256 18284
rect 12308 18272 12314 18284
rect 12912 18281 12940 18312
rect 13449 18309 13461 18343
rect 13495 18340 13507 18343
rect 14550 18340 14556 18352
rect 13495 18312 14556 18340
rect 13495 18309 13507 18312
rect 13449 18303 13507 18309
rect 14550 18300 14556 18312
rect 14608 18300 14614 18352
rect 16960 18340 16988 18380
rect 17218 18368 17224 18380
rect 17276 18368 17282 18420
rect 19150 18368 19156 18420
rect 19208 18408 19214 18420
rect 20257 18411 20315 18417
rect 20257 18408 20269 18411
rect 19208 18380 20269 18408
rect 19208 18368 19214 18380
rect 20257 18377 20269 18380
rect 20303 18377 20315 18411
rect 20257 18371 20315 18377
rect 15028 18312 16988 18340
rect 17037 18343 17095 18349
rect 12897 18275 12955 18281
rect 12308 18244 12848 18272
rect 12308 18232 12314 18244
rect 12710 18204 12716 18216
rect 10787 18176 12716 18204
rect 10689 18167 10747 18173
rect 12710 18164 12716 18176
rect 12768 18164 12774 18216
rect 12820 18204 12848 18244
rect 12897 18241 12909 18275
rect 12943 18241 12955 18275
rect 13078 18272 13084 18284
rect 13039 18244 13084 18272
rect 12897 18235 12955 18241
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 14093 18275 14151 18281
rect 14093 18241 14105 18275
rect 14139 18272 14151 18275
rect 14182 18272 14188 18284
rect 14139 18244 14188 18272
rect 14139 18241 14151 18244
rect 14093 18235 14151 18241
rect 14182 18232 14188 18244
rect 14240 18232 14246 18284
rect 14274 18232 14280 18284
rect 14332 18272 14338 18284
rect 15028 18272 15056 18312
rect 15194 18272 15200 18284
rect 14332 18244 15056 18272
rect 15155 18244 15200 18272
rect 14332 18232 14338 18244
rect 15194 18232 15200 18244
rect 15252 18232 15258 18284
rect 15304 18281 15332 18312
rect 17037 18309 17049 18343
rect 17083 18340 17095 18343
rect 17954 18340 17960 18352
rect 17083 18312 17960 18340
rect 17083 18309 17095 18312
rect 17037 18303 17095 18309
rect 17954 18300 17960 18312
rect 18012 18300 18018 18352
rect 18598 18300 18604 18352
rect 18656 18340 18662 18352
rect 21818 18340 21824 18352
rect 18656 18312 21824 18340
rect 18656 18300 18662 18312
rect 21818 18300 21824 18312
rect 21876 18300 21882 18352
rect 15289 18275 15347 18281
rect 15289 18241 15301 18275
rect 15335 18241 15347 18275
rect 15289 18235 15347 18241
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18272 15623 18275
rect 16301 18275 16359 18281
rect 16301 18272 16313 18275
rect 15611 18244 16313 18272
rect 15611 18241 15623 18244
rect 15565 18235 15623 18241
rect 16301 18241 16313 18244
rect 16347 18241 16359 18275
rect 17310 18272 17316 18284
rect 16301 18235 16359 18241
rect 16868 18244 17316 18272
rect 13909 18207 13967 18213
rect 13909 18204 13921 18207
rect 12820 18176 13921 18204
rect 13909 18173 13921 18176
rect 13955 18173 13967 18207
rect 13909 18167 13967 18173
rect 15105 18207 15163 18213
rect 15105 18173 15117 18207
rect 15151 18204 15163 18207
rect 16114 18204 16120 18216
rect 15151 18176 15976 18204
rect 16075 18176 16120 18204
rect 15151 18173 15163 18176
rect 15105 18167 15163 18173
rect 10410 18136 10416 18148
rect 8772 18108 10416 18136
rect 10410 18096 10416 18108
rect 10468 18096 10474 18148
rect 10956 18139 11014 18145
rect 10956 18105 10968 18139
rect 11002 18136 11014 18139
rect 11882 18136 11888 18148
rect 11002 18108 11888 18136
rect 11002 18105 11014 18108
rect 10956 18099 11014 18105
rect 11882 18096 11888 18108
rect 11940 18096 11946 18148
rect 11974 18096 11980 18148
rect 12032 18136 12038 18148
rect 13817 18139 13875 18145
rect 13817 18136 13829 18139
rect 12032 18108 13829 18136
rect 12032 18096 12038 18108
rect 13817 18105 13829 18108
rect 13863 18105 13875 18139
rect 13817 18099 13875 18105
rect 13924 18108 14872 18136
rect 8294 18068 8300 18080
rect 6932 18040 8300 18068
rect 8294 18028 8300 18040
rect 8352 18028 8358 18080
rect 8846 18068 8852 18080
rect 8807 18040 8852 18068
rect 8846 18028 8852 18040
rect 8904 18028 8910 18080
rect 9030 18028 9036 18080
rect 9088 18068 9094 18080
rect 9858 18068 9864 18080
rect 9088 18040 9864 18068
rect 9088 18028 9094 18040
rect 9858 18028 9864 18040
rect 9916 18028 9922 18080
rect 12802 18068 12808 18080
rect 12763 18040 12808 18068
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 13078 18028 13084 18080
rect 13136 18068 13142 18080
rect 13924 18068 13952 18108
rect 13136 18040 13952 18068
rect 13136 18028 13142 18040
rect 14458 18028 14464 18080
rect 14516 18068 14522 18080
rect 14737 18071 14795 18077
rect 14737 18068 14749 18071
rect 14516 18040 14749 18068
rect 14516 18028 14522 18040
rect 14737 18037 14749 18040
rect 14783 18037 14795 18071
rect 14844 18068 14872 18108
rect 15378 18096 15384 18148
rect 15436 18136 15442 18148
rect 15948 18136 15976 18176
rect 16114 18164 16120 18176
rect 16172 18164 16178 18216
rect 16758 18204 16764 18216
rect 16224 18176 16764 18204
rect 16224 18136 16252 18176
rect 16758 18164 16764 18176
rect 16816 18164 16822 18216
rect 16868 18213 16896 18244
rect 17310 18232 17316 18244
rect 17368 18232 17374 18284
rect 17497 18275 17555 18281
rect 17497 18241 17509 18275
rect 17543 18272 17555 18275
rect 18506 18272 18512 18284
rect 17543 18244 18512 18272
rect 17543 18241 17555 18244
rect 17497 18235 17555 18241
rect 18506 18232 18512 18244
rect 18564 18232 18570 18284
rect 19061 18275 19119 18281
rect 19061 18241 19073 18275
rect 19107 18241 19119 18275
rect 19061 18235 19119 18241
rect 16853 18207 16911 18213
rect 16853 18173 16865 18207
rect 16899 18173 16911 18207
rect 17218 18204 17224 18216
rect 17179 18176 17224 18204
rect 16853 18167 16911 18173
rect 17218 18164 17224 18176
rect 17276 18164 17282 18216
rect 18049 18207 18107 18213
rect 18049 18204 18061 18207
rect 17788 18176 18061 18204
rect 15436 18108 15680 18136
rect 15948 18108 16252 18136
rect 15436 18096 15442 18108
rect 15565 18071 15623 18077
rect 15565 18068 15577 18071
rect 14844 18040 15577 18068
rect 14737 18031 14795 18037
rect 15565 18037 15577 18040
rect 15611 18037 15623 18071
rect 15652 18068 15680 18108
rect 16298 18096 16304 18148
rect 16356 18136 16362 18148
rect 17788 18136 17816 18176
rect 18049 18173 18061 18176
rect 18095 18173 18107 18207
rect 18049 18167 18107 18173
rect 16356 18108 17816 18136
rect 16356 18096 16362 18108
rect 17954 18096 17960 18148
rect 18012 18136 18018 18148
rect 18877 18139 18935 18145
rect 18877 18136 18889 18139
rect 18012 18108 18889 18136
rect 18012 18096 18018 18108
rect 18877 18105 18889 18108
rect 18923 18105 18935 18139
rect 19076 18136 19104 18235
rect 19242 18232 19248 18284
rect 19300 18272 19306 18284
rect 19705 18275 19763 18281
rect 19705 18272 19717 18275
rect 19300 18244 19717 18272
rect 19300 18232 19306 18244
rect 19705 18241 19717 18244
rect 19751 18241 19763 18275
rect 19705 18235 19763 18241
rect 20530 18232 20536 18284
rect 20588 18272 20594 18284
rect 20809 18275 20867 18281
rect 20809 18272 20821 18275
rect 20588 18244 20821 18272
rect 20588 18232 20594 18244
rect 20809 18241 20821 18244
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 19150 18164 19156 18216
rect 19208 18204 19214 18216
rect 19521 18207 19579 18213
rect 19521 18204 19533 18207
rect 19208 18176 19533 18204
rect 19208 18164 19214 18176
rect 19521 18173 19533 18176
rect 19567 18173 19579 18207
rect 20548 18204 20576 18232
rect 19521 18167 19579 18173
rect 19812 18176 20576 18204
rect 19812 18136 19840 18176
rect 19076 18108 19840 18136
rect 18877 18099 18935 18105
rect 19886 18096 19892 18148
rect 19944 18136 19950 18148
rect 20717 18139 20775 18145
rect 20717 18136 20729 18139
rect 19944 18108 20729 18136
rect 19944 18096 19950 18108
rect 20717 18105 20729 18108
rect 20763 18105 20775 18139
rect 20717 18099 20775 18105
rect 16209 18071 16267 18077
rect 16209 18068 16221 18071
rect 15652 18040 16221 18068
rect 15565 18031 15623 18037
rect 16209 18037 16221 18040
rect 16255 18037 16267 18071
rect 16209 18031 16267 18037
rect 16390 18028 16396 18080
rect 16448 18068 16454 18080
rect 17678 18068 17684 18080
rect 16448 18040 17684 18068
rect 16448 18028 16454 18040
rect 17678 18028 17684 18040
rect 17736 18028 17742 18080
rect 18230 18068 18236 18080
rect 18191 18040 18236 18068
rect 18230 18028 18236 18040
rect 18288 18028 18294 18080
rect 18414 18068 18420 18080
rect 18375 18040 18420 18068
rect 18414 18028 18420 18040
rect 18472 18028 18478 18080
rect 18785 18071 18843 18077
rect 18785 18037 18797 18071
rect 18831 18068 18843 18071
rect 19150 18068 19156 18080
rect 18831 18040 19156 18068
rect 18831 18037 18843 18040
rect 18785 18031 18843 18037
rect 19150 18028 19156 18040
rect 19208 18028 19214 18080
rect 20622 18068 20628 18080
rect 20583 18040 20628 18068
rect 20622 18028 20628 18040
rect 20680 18028 20686 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 1765 17867 1823 17873
rect 1765 17864 1777 17867
rect 1728 17836 1777 17864
rect 1728 17824 1734 17836
rect 1765 17833 1777 17836
rect 1811 17833 1823 17867
rect 1765 17827 1823 17833
rect 2409 17867 2467 17873
rect 2409 17833 2421 17867
rect 2455 17864 2467 17867
rect 2866 17864 2872 17876
rect 2455 17836 2636 17864
rect 2827 17836 2872 17864
rect 2455 17833 2467 17836
rect 2409 17827 2467 17833
rect 198 17756 204 17808
rect 256 17796 262 17808
rect 1854 17796 1860 17808
rect 256 17768 1860 17796
rect 256 17756 262 17768
rect 1854 17756 1860 17768
rect 1912 17756 1918 17808
rect 2608 17796 2636 17836
rect 2866 17824 2872 17836
rect 2924 17824 2930 17876
rect 3418 17824 3424 17876
rect 3476 17864 3482 17876
rect 4065 17867 4123 17873
rect 4065 17864 4077 17867
rect 3476 17836 4077 17864
rect 3476 17824 3482 17836
rect 4065 17833 4077 17836
rect 4111 17833 4123 17867
rect 4065 17827 4123 17833
rect 4338 17824 4344 17876
rect 4396 17864 4402 17876
rect 4525 17867 4583 17873
rect 4525 17864 4537 17867
rect 4396 17836 4537 17864
rect 4396 17824 4402 17836
rect 4525 17833 4537 17836
rect 4571 17833 4583 17867
rect 5074 17864 5080 17876
rect 5035 17836 5080 17864
rect 4525 17827 4583 17833
rect 5074 17824 5080 17836
rect 5132 17824 5138 17876
rect 5994 17864 6000 17876
rect 5184 17836 6000 17864
rect 4433 17799 4491 17805
rect 4433 17796 4445 17799
rect 2608 17768 4445 17796
rect 4433 17765 4445 17768
rect 4479 17765 4491 17799
rect 5184 17796 5212 17836
rect 5994 17824 6000 17836
rect 6052 17824 6058 17876
rect 6086 17824 6092 17876
rect 6144 17864 6150 17876
rect 7285 17867 7343 17873
rect 7285 17864 7297 17867
rect 6144 17836 7297 17864
rect 6144 17824 6150 17836
rect 7285 17833 7297 17836
rect 7331 17833 7343 17867
rect 8570 17864 8576 17876
rect 8531 17836 8576 17864
rect 7285 17827 7343 17833
rect 8570 17824 8576 17836
rect 8628 17824 8634 17876
rect 9214 17824 9220 17876
rect 9272 17864 9278 17876
rect 11333 17867 11391 17873
rect 9272 17836 11284 17864
rect 9272 17824 9278 17836
rect 4433 17759 4491 17765
rect 4540 17768 5212 17796
rect 2590 17688 2596 17740
rect 2648 17728 2654 17740
rect 2777 17731 2835 17737
rect 2777 17728 2789 17731
rect 2648 17700 2789 17728
rect 2648 17688 2654 17700
rect 2777 17697 2789 17700
rect 2823 17697 2835 17731
rect 2777 17691 2835 17697
rect 3050 17688 3056 17740
rect 3108 17728 3114 17740
rect 3326 17728 3332 17740
rect 3108 17700 3332 17728
rect 3108 17688 3114 17700
rect 3326 17688 3332 17700
rect 3384 17688 3390 17740
rect 3421 17731 3479 17737
rect 3421 17697 3433 17731
rect 3467 17728 3479 17731
rect 4540 17728 4568 17768
rect 5258 17756 5264 17808
rect 5316 17796 5322 17808
rect 7653 17799 7711 17805
rect 7653 17796 7665 17799
rect 5316 17768 7665 17796
rect 5316 17756 5322 17768
rect 7653 17765 7665 17768
rect 7699 17765 7711 17799
rect 7653 17759 7711 17765
rect 7926 17756 7932 17808
rect 7984 17796 7990 17808
rect 7984 17768 9628 17796
rect 7984 17756 7990 17768
rect 5442 17728 5448 17740
rect 3467 17700 4568 17728
rect 5403 17700 5448 17728
rect 3467 17697 3479 17700
rect 3421 17691 3479 17697
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 5810 17688 5816 17740
rect 5868 17728 5874 17740
rect 6641 17731 6699 17737
rect 6641 17728 6653 17731
rect 5868 17700 6653 17728
rect 5868 17688 5874 17700
rect 6641 17697 6653 17700
rect 6687 17697 6699 17731
rect 6641 17691 6699 17697
rect 6730 17688 6736 17740
rect 6788 17728 6794 17740
rect 6788 17700 6833 17728
rect 6788 17688 6794 17700
rect 7834 17688 7840 17740
rect 7892 17728 7898 17740
rect 8941 17731 8999 17737
rect 8941 17728 8953 17731
rect 7892 17700 8953 17728
rect 7892 17688 7898 17700
rect 8941 17697 8953 17700
rect 8987 17697 8999 17731
rect 8941 17691 8999 17697
rect 9033 17731 9091 17737
rect 9033 17697 9045 17731
rect 9079 17728 9091 17731
rect 9214 17728 9220 17740
rect 9079 17700 9220 17728
rect 9079 17697 9091 17700
rect 9033 17691 9091 17697
rect 9214 17688 9220 17700
rect 9272 17688 9278 17740
rect 9600 17728 9628 17768
rect 9766 17756 9772 17808
rect 9824 17796 9830 17808
rect 10413 17799 10471 17805
rect 10413 17796 10425 17799
rect 9824 17768 10425 17796
rect 9824 17756 9830 17768
rect 10413 17765 10425 17768
rect 10459 17765 10471 17799
rect 11256 17796 11284 17836
rect 11333 17833 11345 17867
rect 11379 17864 11391 17867
rect 12342 17864 12348 17876
rect 11379 17836 12348 17864
rect 11379 17833 11391 17836
rect 11333 17827 11391 17833
rect 12342 17824 12348 17836
rect 12400 17824 12406 17876
rect 12989 17867 13047 17873
rect 12989 17833 13001 17867
rect 13035 17864 13047 17867
rect 13354 17864 13360 17876
rect 13035 17836 13360 17864
rect 13035 17833 13047 17836
rect 12989 17827 13047 17833
rect 13354 17824 13360 17836
rect 13412 17824 13418 17876
rect 14550 17824 14556 17876
rect 14608 17864 14614 17876
rect 14645 17867 14703 17873
rect 14645 17864 14657 17867
rect 14608 17836 14657 17864
rect 14608 17824 14614 17836
rect 14645 17833 14657 17836
rect 14691 17833 14703 17867
rect 14645 17827 14703 17833
rect 15289 17867 15347 17873
rect 15289 17833 15301 17867
rect 15335 17833 15347 17867
rect 15289 17827 15347 17833
rect 11974 17796 11980 17808
rect 11256 17768 11980 17796
rect 10413 17759 10471 17765
rect 11974 17756 11980 17768
rect 12032 17756 12038 17808
rect 12069 17799 12127 17805
rect 12069 17765 12081 17799
rect 12115 17796 12127 17799
rect 12250 17796 12256 17808
rect 12115 17768 12256 17796
rect 12115 17765 12127 17768
rect 12069 17759 12127 17765
rect 12250 17756 12256 17768
rect 12308 17756 12314 17808
rect 13170 17756 13176 17808
rect 13228 17796 13234 17808
rect 13725 17799 13783 17805
rect 13725 17796 13737 17799
rect 13228 17768 13737 17796
rect 13228 17756 13234 17768
rect 13725 17765 13737 17768
rect 13771 17765 13783 17799
rect 15194 17796 15200 17808
rect 13725 17759 13783 17765
rect 14476 17768 15200 17796
rect 10042 17728 10048 17740
rect 9600 17700 10048 17728
rect 10042 17688 10048 17700
rect 10100 17688 10106 17740
rect 10318 17728 10324 17740
rect 10279 17700 10324 17728
rect 10318 17688 10324 17700
rect 10376 17688 10382 17740
rect 11146 17728 11152 17740
rect 10428 17700 10723 17728
rect 11107 17700 11152 17728
rect 2041 17663 2099 17669
rect 2041 17629 2053 17663
rect 2087 17660 2099 17663
rect 2222 17660 2228 17672
rect 2087 17632 2228 17660
rect 2087 17629 2099 17632
rect 2041 17623 2099 17629
rect 2222 17620 2228 17632
rect 2280 17620 2286 17672
rect 2958 17660 2964 17672
rect 2871 17632 2964 17660
rect 2958 17620 2964 17632
rect 3016 17660 3022 17672
rect 3234 17660 3240 17672
rect 3016 17632 3240 17660
rect 3016 17620 3022 17632
rect 3234 17620 3240 17632
rect 3292 17620 3298 17672
rect 4706 17660 4712 17672
rect 4619 17632 4712 17660
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 5534 17660 5540 17672
rect 5495 17632 5540 17660
rect 5534 17620 5540 17632
rect 5592 17620 5598 17672
rect 5629 17663 5687 17669
rect 5629 17629 5641 17663
rect 5675 17629 5687 17663
rect 5629 17623 5687 17629
rect 1397 17595 1455 17601
rect 1397 17561 1409 17595
rect 1443 17592 1455 17595
rect 3602 17592 3608 17604
rect 1443 17564 2544 17592
rect 3563 17564 3608 17592
rect 1443 17561 1455 17564
rect 1397 17555 1455 17561
rect 2516 17524 2544 17564
rect 3602 17552 3608 17564
rect 3660 17552 3666 17604
rect 4724 17592 4752 17620
rect 5644 17592 5672 17623
rect 6270 17620 6276 17672
rect 6328 17660 6334 17672
rect 6917 17663 6975 17669
rect 6917 17660 6929 17663
rect 6328 17632 6929 17660
rect 6328 17620 6334 17632
rect 6917 17629 6929 17632
rect 6963 17629 6975 17663
rect 6917 17623 6975 17629
rect 7466 17620 7472 17672
rect 7524 17660 7530 17672
rect 7745 17663 7803 17669
rect 7745 17660 7757 17663
rect 7524 17632 7757 17660
rect 7524 17620 7530 17632
rect 7745 17629 7757 17632
rect 7791 17629 7803 17663
rect 7745 17623 7803 17629
rect 7929 17663 7987 17669
rect 7929 17629 7941 17663
rect 7975 17660 7987 17663
rect 8294 17660 8300 17672
rect 7975 17632 8300 17660
rect 7975 17629 7987 17632
rect 7929 17623 7987 17629
rect 8294 17620 8300 17632
rect 8352 17620 8358 17672
rect 9122 17660 9128 17672
rect 9083 17632 9128 17660
rect 9122 17620 9128 17632
rect 9180 17620 9186 17672
rect 10428 17660 10456 17700
rect 9232 17632 10456 17660
rect 10597 17663 10655 17669
rect 4724 17564 5672 17592
rect 5994 17552 6000 17604
rect 6052 17592 6058 17604
rect 9232 17592 9260 17632
rect 10597 17629 10609 17663
rect 10643 17629 10655 17663
rect 10695 17660 10723 17700
rect 11146 17688 11152 17700
rect 11204 17688 11210 17740
rect 12805 17731 12863 17737
rect 12805 17697 12817 17731
rect 12851 17697 12863 17731
rect 13446 17728 13452 17740
rect 13407 17700 13452 17728
rect 12805 17691 12863 17697
rect 12158 17660 12164 17672
rect 10695 17632 12164 17660
rect 10597 17623 10655 17629
rect 6052 17564 9260 17592
rect 10612 17592 10640 17623
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 12253 17663 12311 17669
rect 12253 17629 12265 17663
rect 12299 17629 12311 17663
rect 12253 17623 12311 17629
rect 11790 17592 11796 17604
rect 10612 17564 11796 17592
rect 6052 17552 6058 17564
rect 11790 17552 11796 17564
rect 11848 17592 11854 17604
rect 12268 17592 12296 17623
rect 12342 17620 12348 17672
rect 12400 17660 12406 17672
rect 12820 17660 12848 17691
rect 13446 17688 13452 17700
rect 13504 17728 13510 17740
rect 14476 17728 14504 17768
rect 15194 17756 15200 17768
rect 15252 17756 15258 17808
rect 15304 17796 15332 17827
rect 15654 17824 15660 17876
rect 15712 17864 15718 17876
rect 15749 17867 15807 17873
rect 15749 17864 15761 17867
rect 15712 17836 15761 17864
rect 15712 17824 15718 17836
rect 15749 17833 15761 17836
rect 15795 17833 15807 17867
rect 15749 17827 15807 17833
rect 16301 17867 16359 17873
rect 16301 17833 16313 17867
rect 16347 17864 16359 17867
rect 17773 17867 17831 17873
rect 17773 17864 17785 17867
rect 16347 17836 17785 17864
rect 16347 17833 16359 17836
rect 16301 17827 16359 17833
rect 17773 17833 17785 17836
rect 17819 17833 17831 17867
rect 17773 17827 17831 17833
rect 17862 17824 17868 17876
rect 17920 17864 17926 17876
rect 18509 17867 18567 17873
rect 18509 17864 18521 17867
rect 17920 17836 18521 17864
rect 17920 17824 17926 17836
rect 18509 17833 18521 17836
rect 18555 17833 18567 17867
rect 18509 17827 18567 17833
rect 17681 17799 17739 17805
rect 17681 17796 17693 17799
rect 15304 17768 17693 17796
rect 17681 17765 17693 17768
rect 17727 17765 17739 17799
rect 17681 17759 17739 17765
rect 18046 17756 18052 17808
rect 18104 17796 18110 17808
rect 19702 17796 19708 17808
rect 18104 17768 19708 17796
rect 18104 17756 18110 17768
rect 19702 17756 19708 17768
rect 19760 17756 19766 17808
rect 19889 17799 19947 17805
rect 19889 17765 19901 17799
rect 19935 17796 19947 17799
rect 20346 17796 20352 17808
rect 19935 17768 20352 17796
rect 19935 17765 19947 17768
rect 19889 17759 19947 17765
rect 20346 17756 20352 17768
rect 20404 17756 20410 17808
rect 13504 17700 14504 17728
rect 14553 17731 14611 17737
rect 13504 17688 13510 17700
rect 14553 17697 14565 17731
rect 14599 17728 14611 17731
rect 15562 17728 15568 17740
rect 14599 17700 15568 17728
rect 14599 17697 14611 17700
rect 14553 17691 14611 17697
rect 15562 17688 15568 17700
rect 15620 17688 15626 17740
rect 15657 17731 15715 17737
rect 15657 17697 15669 17731
rect 15703 17697 15715 17731
rect 15657 17691 15715 17697
rect 12400 17632 12848 17660
rect 12400 17620 12406 17632
rect 14182 17620 14188 17672
rect 14240 17660 14246 17672
rect 14366 17660 14372 17672
rect 14240 17632 14372 17660
rect 14240 17620 14246 17632
rect 14366 17620 14372 17632
rect 14424 17620 14430 17672
rect 14826 17660 14832 17672
rect 14787 17632 14832 17660
rect 14826 17620 14832 17632
rect 14884 17620 14890 17672
rect 15286 17620 15292 17672
rect 15344 17660 15350 17672
rect 15672 17660 15700 17691
rect 16482 17688 16488 17740
rect 16540 17728 16546 17740
rect 16669 17731 16727 17737
rect 16669 17728 16681 17731
rect 16540 17700 16681 17728
rect 16540 17688 16546 17700
rect 16669 17697 16681 17700
rect 16715 17697 16727 17731
rect 16669 17691 16727 17697
rect 16761 17731 16819 17737
rect 16761 17697 16773 17731
rect 16807 17728 16819 17731
rect 16807 17700 16988 17728
rect 16807 17697 16819 17700
rect 16761 17691 16819 17697
rect 15838 17660 15844 17672
rect 15344 17632 15700 17660
rect 15799 17632 15844 17660
rect 15344 17620 15350 17632
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 16022 17620 16028 17672
rect 16080 17660 16086 17672
rect 16776 17660 16804 17691
rect 16080 17632 16804 17660
rect 16853 17663 16911 17669
rect 16080 17620 16086 17632
rect 16853 17629 16865 17663
rect 16899 17629 16911 17663
rect 16960 17660 16988 17700
rect 17034 17688 17040 17740
rect 17092 17728 17098 17740
rect 18877 17731 18935 17737
rect 18877 17728 18889 17731
rect 17092 17700 18889 17728
rect 17092 17688 17098 17700
rect 18877 17697 18889 17700
rect 18923 17697 18935 17731
rect 18877 17691 18935 17697
rect 19981 17731 20039 17737
rect 19981 17697 19993 17731
rect 20027 17728 20039 17731
rect 20254 17728 20260 17740
rect 20027 17700 20260 17728
rect 20027 17697 20039 17700
rect 19981 17691 20039 17697
rect 20254 17688 20260 17700
rect 20312 17688 20318 17740
rect 17494 17660 17500 17672
rect 16960 17632 17500 17660
rect 16853 17623 16911 17629
rect 15378 17592 15384 17604
rect 11848 17564 12296 17592
rect 14007 17564 15384 17592
rect 11848 17552 11854 17564
rect 4982 17524 4988 17536
rect 2516 17496 4988 17524
rect 4982 17484 4988 17496
rect 5040 17484 5046 17536
rect 6273 17527 6331 17533
rect 6273 17493 6285 17527
rect 6319 17524 6331 17527
rect 9858 17524 9864 17536
rect 6319 17496 9864 17524
rect 6319 17493 6331 17496
rect 6273 17487 6331 17493
rect 9858 17484 9864 17496
rect 9916 17484 9922 17536
rect 9953 17527 10011 17533
rect 9953 17493 9965 17527
rect 9999 17524 10011 17527
rect 11146 17524 11152 17536
rect 9999 17496 11152 17524
rect 9999 17493 10011 17496
rect 9953 17487 10011 17493
rect 11146 17484 11152 17496
rect 11204 17484 11210 17536
rect 11701 17527 11759 17533
rect 11701 17493 11713 17527
rect 11747 17524 11759 17527
rect 14007 17524 14035 17564
rect 15378 17552 15384 17564
rect 15436 17552 15442 17604
rect 15856 17592 15884 17620
rect 16868 17592 16896 17623
rect 17494 17620 17500 17632
rect 17552 17620 17558 17672
rect 17586 17620 17592 17672
rect 17644 17660 17650 17672
rect 17865 17663 17923 17669
rect 17865 17660 17877 17663
rect 17644 17632 17877 17660
rect 17644 17620 17650 17632
rect 17865 17629 17877 17632
rect 17911 17629 17923 17663
rect 17865 17623 17923 17629
rect 18969 17663 19027 17669
rect 18969 17629 18981 17663
rect 19015 17629 19027 17663
rect 18969 17623 19027 17629
rect 15856 17564 16896 17592
rect 11747 17496 14035 17524
rect 14185 17527 14243 17533
rect 11747 17493 11759 17496
rect 11701 17487 11759 17493
rect 14185 17493 14197 17527
rect 14231 17524 14243 17527
rect 15930 17524 15936 17536
rect 14231 17496 15936 17524
rect 14231 17493 14243 17496
rect 14185 17487 14243 17493
rect 15930 17484 15936 17496
rect 15988 17484 15994 17536
rect 17313 17527 17371 17533
rect 17313 17493 17325 17527
rect 17359 17524 17371 17527
rect 17586 17524 17592 17536
rect 17359 17496 17592 17524
rect 17359 17493 17371 17496
rect 17313 17487 17371 17493
rect 17586 17484 17592 17496
rect 17644 17484 17650 17536
rect 17862 17484 17868 17536
rect 17920 17524 17926 17536
rect 18325 17527 18383 17533
rect 18325 17524 18337 17527
rect 17920 17496 18337 17524
rect 17920 17484 17926 17496
rect 18325 17493 18337 17496
rect 18371 17524 18383 17527
rect 18984 17524 19012 17623
rect 19058 17620 19064 17672
rect 19116 17660 19122 17672
rect 20165 17663 20223 17669
rect 19116 17632 19161 17660
rect 19116 17620 19122 17632
rect 20165 17629 20177 17663
rect 20211 17660 20223 17663
rect 20530 17660 20536 17672
rect 20211 17632 20536 17660
rect 20211 17629 20223 17632
rect 20165 17623 20223 17629
rect 20530 17620 20536 17632
rect 20588 17620 20594 17672
rect 19518 17524 19524 17536
rect 18371 17496 19012 17524
rect 19479 17496 19524 17524
rect 18371 17493 18383 17496
rect 18325 17487 18383 17493
rect 19518 17484 19524 17496
rect 19576 17484 19582 17536
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 3418 17280 3424 17332
rect 3476 17320 3482 17332
rect 3513 17323 3571 17329
rect 3513 17320 3525 17323
rect 3476 17292 3525 17320
rect 3476 17280 3482 17292
rect 3513 17289 3525 17292
rect 3559 17320 3571 17323
rect 3602 17320 3608 17332
rect 3559 17292 3608 17320
rect 3559 17289 3571 17292
rect 3513 17283 3571 17289
rect 3602 17280 3608 17292
rect 3660 17280 3666 17332
rect 5169 17323 5227 17329
rect 5169 17289 5181 17323
rect 5215 17320 5227 17323
rect 5810 17320 5816 17332
rect 5215 17292 5816 17320
rect 5215 17289 5227 17292
rect 5169 17283 5227 17289
rect 5810 17280 5816 17292
rect 5868 17280 5874 17332
rect 6546 17280 6552 17332
rect 6604 17320 6610 17332
rect 7926 17320 7932 17332
rect 6604 17292 7932 17320
rect 6604 17280 6610 17292
rect 7926 17280 7932 17292
rect 7984 17280 7990 17332
rect 8389 17323 8447 17329
rect 8389 17289 8401 17323
rect 8435 17320 8447 17323
rect 8846 17320 8852 17332
rect 8435 17292 8852 17320
rect 8435 17289 8447 17292
rect 8389 17283 8447 17289
rect 8846 17280 8852 17292
rect 8904 17280 8910 17332
rect 9766 17280 9772 17332
rect 9824 17320 9830 17332
rect 10870 17320 10876 17332
rect 9824 17292 10876 17320
rect 9824 17280 9830 17292
rect 10870 17280 10876 17292
rect 10928 17280 10934 17332
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 12492 17292 12537 17320
rect 12492 17280 12498 17292
rect 14826 17280 14832 17332
rect 14884 17320 14890 17332
rect 15105 17323 15163 17329
rect 15105 17320 15117 17323
rect 14884 17292 15117 17320
rect 14884 17280 14890 17292
rect 15105 17289 15117 17292
rect 15151 17320 15163 17323
rect 15289 17323 15347 17329
rect 15289 17320 15301 17323
rect 15151 17292 15301 17320
rect 15151 17289 15163 17292
rect 15105 17283 15163 17289
rect 15289 17289 15301 17292
rect 15335 17289 15347 17323
rect 15289 17283 15347 17289
rect 15654 17280 15660 17332
rect 15712 17320 15718 17332
rect 16298 17320 16304 17332
rect 15712 17292 16304 17320
rect 15712 17280 15718 17292
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 16666 17280 16672 17332
rect 16724 17280 16730 17332
rect 17310 17280 17316 17332
rect 17368 17320 17374 17332
rect 17494 17320 17500 17332
rect 17368 17292 17500 17320
rect 17368 17280 17374 17292
rect 17494 17280 17500 17292
rect 17552 17280 17558 17332
rect 18049 17323 18107 17329
rect 18049 17289 18061 17323
rect 18095 17320 18107 17323
rect 19978 17320 19984 17332
rect 18095 17292 19984 17320
rect 18095 17289 18107 17292
rect 18049 17283 18107 17289
rect 19978 17280 19984 17292
rect 20036 17280 20042 17332
rect 20714 17280 20720 17332
rect 20772 17320 20778 17332
rect 21266 17320 21272 17332
rect 20772 17292 21272 17320
rect 20772 17280 20778 17292
rect 21266 17280 21272 17292
rect 21324 17280 21330 17332
rect 4065 17255 4123 17261
rect 4065 17221 4077 17255
rect 4111 17221 4123 17255
rect 4065 17215 4123 17221
rect 3786 17144 3792 17196
rect 3844 17184 3850 17196
rect 4080 17184 4108 17215
rect 4246 17212 4252 17264
rect 4304 17252 4310 17264
rect 5902 17252 5908 17264
rect 4304 17224 5908 17252
rect 4304 17212 4310 17224
rect 5902 17212 5908 17224
rect 5960 17212 5966 17264
rect 7834 17252 7840 17264
rect 6288 17224 7840 17252
rect 4706 17184 4712 17196
rect 3844 17156 4108 17184
rect 4667 17156 4712 17184
rect 3844 17144 3850 17156
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 5718 17144 5724 17196
rect 5776 17184 5782 17196
rect 6288 17193 6316 17224
rect 7834 17212 7840 17224
rect 7892 17212 7898 17264
rect 8018 17252 8024 17264
rect 7979 17224 8024 17252
rect 8018 17212 8024 17224
rect 8076 17212 8082 17264
rect 11977 17255 12035 17261
rect 9140 17224 11008 17252
rect 9140 17196 9168 17224
rect 5813 17187 5871 17193
rect 5813 17184 5825 17187
rect 5776 17156 5825 17184
rect 5776 17144 5782 17156
rect 5813 17153 5825 17156
rect 5859 17153 5871 17187
rect 5813 17147 5871 17153
rect 6273 17187 6331 17193
rect 6273 17153 6285 17187
rect 6319 17153 6331 17187
rect 6273 17147 6331 17153
rect 7190 17144 7196 17196
rect 7248 17184 7254 17196
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 7248 17156 7389 17184
rect 7248 17144 7254 17156
rect 7377 17153 7389 17156
rect 7423 17153 7435 17187
rect 7377 17147 7435 17153
rect 8386 17144 8392 17196
rect 8444 17184 8450 17196
rect 8846 17184 8852 17196
rect 8444 17156 8852 17184
rect 8444 17144 8450 17156
rect 8846 17144 8852 17156
rect 8904 17144 8910 17196
rect 9033 17187 9091 17193
rect 9033 17153 9045 17187
rect 9079 17184 9091 17187
rect 9122 17184 9128 17196
rect 9079 17156 9128 17184
rect 9079 17153 9091 17156
rect 9033 17147 9091 17153
rect 9122 17144 9128 17156
rect 9180 17144 9186 17196
rect 9582 17144 9588 17196
rect 9640 17184 9646 17196
rect 10980 17193 11008 17224
rect 11977 17221 11989 17255
rect 12023 17252 12035 17255
rect 12526 17252 12532 17264
rect 12023 17224 12532 17252
rect 12023 17221 12035 17224
rect 11977 17215 12035 17221
rect 12526 17212 12532 17224
rect 12584 17212 12590 17264
rect 12618 17212 12624 17264
rect 12676 17252 12682 17264
rect 16684 17252 16712 17280
rect 17129 17255 17187 17261
rect 17129 17252 17141 17255
rect 12676 17224 13768 17252
rect 16684 17224 17141 17252
rect 12676 17212 12682 17224
rect 9953 17187 10011 17193
rect 9953 17184 9965 17187
rect 9640 17156 9965 17184
rect 9640 17144 9646 17156
rect 9953 17153 9965 17156
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 10321 17187 10379 17193
rect 10321 17153 10333 17187
rect 10367 17184 10379 17187
rect 10965 17187 11023 17193
rect 10367 17156 10916 17184
rect 10367 17153 10379 17156
rect 10321 17147 10379 17153
rect 1210 17076 1216 17128
rect 1268 17116 1274 17128
rect 1397 17119 1455 17125
rect 1397 17116 1409 17119
rect 1268 17088 1409 17116
rect 1268 17076 1274 17088
rect 1397 17085 1409 17088
rect 1443 17085 1455 17119
rect 1397 17079 1455 17085
rect 1762 17076 1768 17128
rect 1820 17116 1826 17128
rect 2038 17116 2044 17128
rect 1820 17088 2044 17116
rect 1820 17076 1826 17088
rect 2038 17076 2044 17088
rect 2096 17116 2102 17128
rect 2133 17119 2191 17125
rect 2133 17116 2145 17119
rect 2096 17088 2145 17116
rect 2096 17076 2102 17088
rect 2133 17085 2145 17088
rect 2179 17085 2191 17119
rect 2133 17079 2191 17085
rect 2400 17119 2458 17125
rect 2400 17085 2412 17119
rect 2446 17116 2458 17119
rect 2682 17116 2688 17128
rect 2446 17088 2688 17116
rect 2446 17085 2458 17088
rect 2400 17079 2458 17085
rect 2682 17076 2688 17088
rect 2740 17076 2746 17128
rect 3142 17076 3148 17128
rect 3200 17116 3206 17128
rect 3970 17116 3976 17128
rect 3200 17088 3976 17116
rect 3200 17076 3206 17088
rect 3970 17076 3976 17088
rect 4028 17076 4034 17128
rect 4982 17076 4988 17128
rect 5040 17116 5046 17128
rect 7285 17119 7343 17125
rect 7285 17116 7297 17119
rect 5040 17088 7297 17116
rect 5040 17076 5046 17088
rect 7285 17085 7297 17088
rect 7331 17085 7343 17119
rect 7285 17079 7343 17085
rect 7837 17119 7895 17125
rect 7837 17085 7849 17119
rect 7883 17116 7895 17119
rect 10778 17116 10784 17128
rect 7883 17088 10784 17116
rect 7883 17085 7895 17088
rect 7837 17079 7895 17085
rect 10778 17076 10784 17088
rect 10836 17076 10842 17128
rect 10888 17116 10916 17156
rect 10965 17153 10977 17187
rect 11011 17153 11023 17187
rect 10965 17147 11023 17153
rect 11146 17144 11152 17196
rect 11204 17184 11210 17196
rect 12897 17187 12955 17193
rect 12897 17184 12909 17187
rect 11204 17156 12909 17184
rect 11204 17144 11210 17156
rect 12897 17153 12909 17156
rect 12943 17153 12955 17187
rect 13078 17184 13084 17196
rect 13039 17156 13084 17184
rect 12897 17147 12955 17153
rect 13078 17144 13084 17156
rect 13136 17144 13142 17196
rect 13740 17184 13768 17224
rect 17129 17221 17141 17224
rect 17175 17221 17187 17255
rect 17129 17215 17187 17221
rect 15378 17184 15384 17196
rect 13740 17156 13860 17184
rect 15339 17156 15384 17184
rect 11793 17119 11851 17125
rect 11793 17116 11805 17119
rect 10888 17088 11805 17116
rect 11793 17085 11805 17088
rect 11839 17085 11851 17119
rect 11793 17079 11851 17085
rect 11882 17076 11888 17128
rect 11940 17116 11946 17128
rect 13096 17116 13124 17144
rect 11940 17088 13124 17116
rect 11940 17076 11946 17088
rect 13630 17076 13636 17128
rect 13688 17116 13694 17128
rect 13725 17119 13783 17125
rect 13725 17116 13737 17119
rect 13688 17088 13737 17116
rect 13688 17076 13694 17088
rect 13725 17085 13737 17088
rect 13771 17085 13783 17119
rect 13832 17116 13860 17156
rect 15378 17144 15384 17156
rect 15436 17144 15442 17196
rect 16666 17144 16672 17196
rect 16724 17184 16730 17196
rect 17681 17187 17739 17193
rect 17681 17184 17693 17187
rect 16724 17156 17693 17184
rect 16724 17144 16730 17156
rect 17681 17153 17693 17156
rect 17727 17153 17739 17187
rect 17681 17147 17739 17153
rect 18693 17187 18751 17193
rect 18693 17153 18705 17187
rect 18739 17184 18751 17187
rect 18874 17184 18880 17196
rect 18739 17156 18880 17184
rect 18739 17153 18751 17156
rect 18693 17147 18751 17153
rect 18874 17144 18880 17156
rect 18932 17144 18938 17196
rect 19702 17184 19708 17196
rect 19663 17156 19708 17184
rect 19702 17144 19708 17156
rect 19760 17144 19766 17196
rect 20530 17144 20536 17196
rect 20588 17184 20594 17196
rect 20717 17187 20775 17193
rect 20717 17184 20729 17187
rect 20588 17156 20729 17184
rect 20588 17144 20594 17156
rect 20717 17153 20729 17156
rect 20763 17184 20775 17187
rect 21542 17184 21548 17196
rect 20763 17156 21548 17184
rect 20763 17153 20775 17156
rect 20717 17147 20775 17153
rect 21542 17144 21548 17156
rect 21600 17144 21606 17196
rect 17034 17116 17040 17128
rect 13832 17088 17040 17116
rect 13725 17079 13783 17085
rect 17034 17076 17040 17088
rect 17092 17076 17098 17128
rect 17586 17076 17592 17128
rect 17644 17116 17650 17128
rect 19429 17119 19487 17125
rect 19429 17116 19441 17119
rect 17644 17088 19441 17116
rect 17644 17076 17650 17088
rect 19429 17085 19441 17088
rect 19475 17085 19487 17119
rect 19429 17079 19487 17085
rect 1673 17051 1731 17057
rect 1673 17017 1685 17051
rect 1719 17017 1731 17051
rect 1673 17011 1731 17017
rect 1688 16980 1716 17011
rect 2498 17008 2504 17060
rect 2556 17048 2562 17060
rect 4433 17051 4491 17057
rect 4433 17048 4445 17051
rect 2556 17020 4445 17048
rect 2556 17008 2562 17020
rect 4433 17017 4445 17020
rect 4479 17017 4491 17051
rect 4433 17011 4491 17017
rect 4525 17051 4583 17057
rect 4525 17017 4537 17051
rect 4571 17048 4583 17051
rect 4571 17020 5304 17048
rect 4571 17017 4583 17020
rect 4525 17011 4583 17017
rect 5074 16980 5080 16992
rect 1688 16952 5080 16980
rect 5074 16940 5080 16952
rect 5132 16940 5138 16992
rect 5276 16989 5304 17020
rect 6638 17008 6644 17060
rect 6696 17048 6702 17060
rect 7193 17051 7251 17057
rect 7193 17048 7205 17051
rect 6696 17020 7205 17048
rect 6696 17008 6702 17020
rect 7193 17017 7205 17020
rect 7239 17017 7251 17051
rect 7193 17011 7251 17017
rect 8757 17051 8815 17057
rect 8757 17017 8769 17051
rect 8803 17048 8815 17051
rect 8803 17020 9444 17048
rect 8803 17017 8815 17020
rect 8757 17011 8815 17017
rect 5261 16983 5319 16989
rect 5261 16949 5273 16983
rect 5307 16949 5319 16983
rect 5626 16980 5632 16992
rect 5587 16952 5632 16980
rect 5261 16943 5319 16949
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 5721 16983 5779 16989
rect 5721 16949 5733 16983
rect 5767 16980 5779 16983
rect 5810 16980 5816 16992
rect 5767 16952 5816 16980
rect 5767 16949 5779 16952
rect 5721 16943 5779 16949
rect 5810 16940 5816 16952
rect 5868 16940 5874 16992
rect 6822 16980 6828 16992
rect 6783 16952 6828 16980
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 8846 16980 8852 16992
rect 8807 16952 8852 16980
rect 8846 16940 8852 16952
rect 8904 16940 8910 16992
rect 9416 16989 9444 17020
rect 9674 17008 9680 17060
rect 9732 17048 9738 17060
rect 9861 17051 9919 17057
rect 9861 17048 9873 17051
rect 9732 17020 9873 17048
rect 9732 17008 9738 17020
rect 9861 17017 9873 17020
rect 9907 17017 9919 17051
rect 9861 17011 9919 17017
rect 10873 17051 10931 17057
rect 10873 17017 10885 17051
rect 10919 17048 10931 17051
rect 11146 17048 11152 17060
rect 10919 17020 11152 17048
rect 10919 17017 10931 17020
rect 10873 17011 10931 17017
rect 11146 17008 11152 17020
rect 11204 17008 11210 17060
rect 12526 17008 12532 17060
rect 12584 17048 12590 17060
rect 13814 17048 13820 17060
rect 12584 17020 13820 17048
rect 12584 17008 12590 17020
rect 13814 17008 13820 17020
rect 13872 17008 13878 17060
rect 13998 17057 14004 17060
rect 13992 17048 14004 17057
rect 13959 17020 14004 17048
rect 13992 17011 14004 17020
rect 13998 17008 14004 17011
rect 14056 17008 14062 17060
rect 15194 17008 15200 17060
rect 15252 17048 15258 17060
rect 15289 17051 15347 17057
rect 15289 17048 15301 17051
rect 15252 17020 15301 17048
rect 15252 17008 15258 17020
rect 15289 17017 15301 17020
rect 15335 17048 15347 17051
rect 15626 17051 15684 17057
rect 15626 17048 15638 17051
rect 15335 17020 15638 17048
rect 15335 17017 15347 17020
rect 15289 17011 15347 17017
rect 15626 17017 15638 17020
rect 15672 17017 15684 17051
rect 18322 17048 18328 17060
rect 15626 17011 15684 17017
rect 15764 17020 18328 17048
rect 9401 16983 9459 16989
rect 9401 16949 9413 16983
rect 9447 16949 9459 16983
rect 9401 16943 9459 16949
rect 9490 16940 9496 16992
rect 9548 16980 9554 16992
rect 9769 16983 9827 16989
rect 9769 16980 9781 16983
rect 9548 16952 9781 16980
rect 9548 16940 9554 16952
rect 9769 16949 9781 16952
rect 9815 16980 9827 16983
rect 10321 16983 10379 16989
rect 10321 16980 10333 16983
rect 9815 16952 10333 16980
rect 9815 16949 9827 16952
rect 9769 16943 9827 16949
rect 10321 16949 10333 16952
rect 10367 16949 10379 16983
rect 10321 16943 10379 16949
rect 10410 16940 10416 16992
rect 10468 16980 10474 16992
rect 10781 16983 10839 16989
rect 10468 16952 10513 16980
rect 10468 16940 10474 16952
rect 10781 16949 10793 16983
rect 10827 16980 10839 16983
rect 11974 16980 11980 16992
rect 10827 16952 11980 16980
rect 10827 16949 10839 16952
rect 10781 16943 10839 16949
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 12802 16980 12808 16992
rect 12763 16952 12808 16980
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 13078 16940 13084 16992
rect 13136 16980 13142 16992
rect 15764 16980 15792 17020
rect 18322 17008 18328 17020
rect 18380 17008 18386 17060
rect 18509 17051 18567 17057
rect 18509 17017 18521 17051
rect 18555 17048 18567 17051
rect 19150 17048 19156 17060
rect 18555 17020 19156 17048
rect 18555 17017 18567 17020
rect 18509 17011 18567 17017
rect 19150 17008 19156 17020
rect 19208 17008 19214 17060
rect 19242 17008 19248 17060
rect 19300 17048 19306 17060
rect 19521 17051 19579 17057
rect 19521 17048 19533 17051
rect 19300 17020 19533 17048
rect 19300 17008 19306 17020
rect 19521 17017 19533 17020
rect 19567 17017 19579 17051
rect 19521 17011 19579 17017
rect 20441 17051 20499 17057
rect 20441 17017 20453 17051
rect 20487 17048 20499 17051
rect 21082 17048 21088 17060
rect 20487 17020 21088 17048
rect 20487 17017 20499 17020
rect 20441 17011 20499 17017
rect 21082 17008 21088 17020
rect 21140 17008 21146 17060
rect 13136 16952 15792 16980
rect 16761 16983 16819 16989
rect 13136 16940 13142 16952
rect 16761 16949 16773 16983
rect 16807 16980 16819 16983
rect 16942 16980 16948 16992
rect 16807 16952 16948 16980
rect 16807 16949 16819 16952
rect 16761 16943 16819 16949
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17034 16940 17040 16992
rect 17092 16980 17098 16992
rect 17497 16983 17555 16989
rect 17497 16980 17509 16983
rect 17092 16952 17509 16980
rect 17092 16940 17098 16952
rect 17497 16949 17509 16952
rect 17543 16949 17555 16983
rect 17497 16943 17555 16949
rect 17589 16983 17647 16989
rect 17589 16949 17601 16983
rect 17635 16980 17647 16983
rect 17954 16980 17960 16992
rect 17635 16952 17960 16980
rect 17635 16949 17647 16952
rect 17589 16943 17647 16949
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 18414 16980 18420 16992
rect 18375 16952 18420 16980
rect 18414 16940 18420 16952
rect 18472 16940 18478 16992
rect 18874 16940 18880 16992
rect 18932 16980 18938 16992
rect 19061 16983 19119 16989
rect 19061 16980 19073 16983
rect 18932 16952 19073 16980
rect 18932 16940 18938 16952
rect 19061 16949 19073 16952
rect 19107 16949 19119 16983
rect 20070 16980 20076 16992
rect 20031 16952 20076 16980
rect 19061 16943 19119 16949
rect 20070 16940 20076 16952
rect 20128 16940 20134 16992
rect 20530 16980 20536 16992
rect 20491 16952 20536 16980
rect 20530 16940 20536 16952
rect 20588 16940 20594 16992
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1949 16779 2007 16785
rect 1949 16745 1961 16779
rect 1995 16776 2007 16779
rect 2498 16776 2504 16788
rect 1995 16748 2504 16776
rect 1995 16745 2007 16748
rect 1949 16739 2007 16745
rect 2498 16736 2504 16748
rect 2556 16736 2562 16788
rect 2961 16779 3019 16785
rect 2961 16745 2973 16779
rect 3007 16776 3019 16779
rect 4246 16776 4252 16788
rect 3007 16748 4252 16776
rect 3007 16745 3019 16748
rect 2961 16739 3019 16745
rect 4246 16736 4252 16748
rect 4304 16736 4310 16788
rect 4522 16776 4528 16788
rect 4483 16748 4528 16776
rect 4522 16736 4528 16748
rect 4580 16736 4586 16788
rect 5074 16736 5080 16788
rect 5132 16776 5138 16788
rect 5350 16776 5356 16788
rect 5132 16748 5356 16776
rect 5132 16736 5138 16748
rect 5350 16736 5356 16748
rect 5408 16736 5414 16788
rect 6362 16736 6368 16788
rect 6420 16776 6426 16788
rect 6638 16776 6644 16788
rect 6420 16748 6644 16776
rect 6420 16736 6426 16748
rect 6638 16736 6644 16748
rect 6696 16736 6702 16788
rect 6822 16736 6828 16788
rect 6880 16776 6886 16788
rect 7377 16779 7435 16785
rect 7377 16776 7389 16779
rect 6880 16748 7389 16776
rect 6880 16736 6886 16748
rect 7377 16745 7389 16748
rect 7423 16745 7435 16779
rect 7377 16739 7435 16745
rect 9309 16779 9367 16785
rect 9309 16745 9321 16779
rect 9355 16776 9367 16779
rect 9582 16776 9588 16788
rect 9355 16748 9588 16776
rect 9355 16745 9367 16748
rect 9309 16739 9367 16745
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 10137 16779 10195 16785
rect 10137 16745 10149 16779
rect 10183 16776 10195 16779
rect 11054 16776 11060 16788
rect 10183 16748 11060 16776
rect 10183 16745 10195 16748
rect 10137 16739 10195 16745
rect 11054 16736 11060 16748
rect 11112 16736 11118 16788
rect 11882 16776 11888 16788
rect 11843 16748 11888 16776
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 13078 16776 13084 16788
rect 11992 16748 13084 16776
rect 1857 16711 1915 16717
rect 1857 16677 1869 16711
rect 1903 16708 1915 16711
rect 2314 16708 2320 16720
rect 1903 16680 2320 16708
rect 1903 16677 1915 16680
rect 1857 16671 1915 16677
rect 2314 16668 2320 16680
rect 2372 16668 2378 16720
rect 2406 16668 2412 16720
rect 2464 16708 2470 16720
rect 2464 16680 2509 16708
rect 2464 16668 2470 16680
rect 3694 16668 3700 16720
rect 3752 16708 3758 16720
rect 4982 16708 4988 16720
rect 3752 16680 4988 16708
rect 3752 16668 3758 16680
rect 4982 16668 4988 16680
rect 5040 16668 5046 16720
rect 5718 16708 5724 16720
rect 5184 16680 5724 16708
rect 3326 16640 3332 16652
rect 3287 16612 3332 16640
rect 3326 16600 3332 16612
rect 3384 16600 3390 16652
rect 3418 16600 3424 16652
rect 3476 16640 3482 16652
rect 4433 16643 4491 16649
rect 3476 16612 3521 16640
rect 3476 16600 3482 16612
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 4798 16640 4804 16652
rect 4479 16612 4804 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 4798 16600 4804 16612
rect 4856 16600 4862 16652
rect 4890 16600 4896 16652
rect 4948 16640 4954 16652
rect 5074 16640 5080 16652
rect 4948 16612 5080 16640
rect 4948 16600 4954 16612
rect 5074 16600 5080 16612
rect 5132 16600 5138 16652
rect 2593 16575 2651 16581
rect 2593 16541 2605 16575
rect 2639 16572 2651 16575
rect 2682 16572 2688 16584
rect 2639 16544 2688 16572
rect 2639 16541 2651 16544
rect 2593 16535 2651 16541
rect 2682 16532 2688 16544
rect 2740 16572 2746 16584
rect 3513 16575 3571 16581
rect 3513 16572 3525 16575
rect 2740 16544 3525 16572
rect 2740 16532 2746 16544
rect 3513 16541 3525 16544
rect 3559 16572 3571 16575
rect 4617 16575 4675 16581
rect 4617 16572 4629 16575
rect 3559 16544 4629 16572
rect 3559 16541 3571 16544
rect 3513 16535 3571 16541
rect 4617 16541 4629 16544
rect 4663 16572 4675 16575
rect 5184 16572 5212 16680
rect 5718 16668 5724 16680
rect 5776 16668 5782 16720
rect 6914 16668 6920 16720
rect 6972 16708 6978 16720
rect 7466 16708 7472 16720
rect 6972 16680 7472 16708
rect 6972 16668 6978 16680
rect 7466 16668 7472 16680
rect 7524 16668 7530 16720
rect 8196 16711 8254 16717
rect 8196 16677 8208 16711
rect 8242 16708 8254 16711
rect 8294 16708 8300 16720
rect 8242 16680 8300 16708
rect 8242 16677 8254 16680
rect 8196 16671 8254 16677
rect 8294 16668 8300 16680
rect 8352 16668 8358 16720
rect 8662 16668 8668 16720
rect 8720 16708 8726 16720
rect 9490 16708 9496 16720
rect 8720 16680 9496 16708
rect 8720 16668 8726 16680
rect 9490 16668 9496 16680
rect 9548 16668 9554 16720
rect 11992 16708 12020 16748
rect 13078 16736 13084 16748
rect 13136 16736 13142 16788
rect 13722 16736 13728 16788
rect 13780 16776 13786 16788
rect 14369 16779 14427 16785
rect 14369 16776 14381 16779
rect 13780 16748 14381 16776
rect 13780 16736 13786 16748
rect 14369 16745 14381 16748
rect 14415 16745 14427 16779
rect 14369 16739 14427 16745
rect 14829 16779 14887 16785
rect 14829 16745 14841 16779
rect 14875 16776 14887 16779
rect 15013 16779 15071 16785
rect 15013 16776 15025 16779
rect 14875 16748 15025 16776
rect 14875 16745 14887 16748
rect 14829 16739 14887 16745
rect 15013 16745 15025 16748
rect 15059 16745 15071 16779
rect 15562 16776 15568 16788
rect 15523 16748 15568 16776
rect 15013 16739 15071 16745
rect 15562 16736 15568 16748
rect 15620 16736 15626 16788
rect 15930 16776 15936 16788
rect 15891 16748 15936 16776
rect 15930 16736 15936 16748
rect 15988 16736 15994 16788
rect 16025 16779 16083 16785
rect 16025 16745 16037 16779
rect 16071 16776 16083 16779
rect 16298 16776 16304 16788
rect 16071 16748 16304 16776
rect 16071 16745 16083 16748
rect 16025 16739 16083 16745
rect 16298 16736 16304 16748
rect 16356 16736 16362 16788
rect 16574 16776 16580 16788
rect 16535 16748 16580 16776
rect 16574 16736 16580 16748
rect 16632 16736 16638 16788
rect 16945 16779 17003 16785
rect 16945 16745 16957 16779
rect 16991 16776 17003 16779
rect 17126 16776 17132 16788
rect 16991 16748 17132 16776
rect 16991 16745 17003 16748
rect 16945 16739 17003 16745
rect 17126 16736 17132 16748
rect 17184 16736 17190 16788
rect 17586 16776 17592 16788
rect 17236 16748 17448 16776
rect 17547 16748 17592 16776
rect 12710 16708 12716 16720
rect 9600 16680 12020 16708
rect 12084 16680 12716 16708
rect 5528 16643 5586 16649
rect 5528 16609 5540 16643
rect 5574 16640 5586 16643
rect 5902 16640 5908 16652
rect 5574 16612 5908 16640
rect 5574 16609 5586 16612
rect 5528 16603 5586 16609
rect 5902 16600 5908 16612
rect 5960 16600 5966 16652
rect 5994 16600 6000 16652
rect 6052 16640 6058 16652
rect 6822 16640 6828 16652
rect 6052 16612 6828 16640
rect 6052 16600 6058 16612
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 7285 16643 7343 16649
rect 7285 16609 7297 16643
rect 7331 16640 7343 16643
rect 8570 16640 8576 16652
rect 7331 16612 8576 16640
rect 7331 16609 7343 16612
rect 7285 16603 7343 16609
rect 8570 16600 8576 16612
rect 8628 16600 8634 16652
rect 9030 16600 9036 16652
rect 9088 16640 9094 16652
rect 9306 16640 9312 16652
rect 9088 16612 9312 16640
rect 9088 16600 9094 16612
rect 9306 16600 9312 16612
rect 9364 16640 9370 16652
rect 9600 16640 9628 16680
rect 9950 16640 9956 16652
rect 9364 16612 9628 16640
rect 9911 16612 9956 16640
rect 9364 16600 9370 16612
rect 9950 16600 9956 16612
rect 10008 16600 10014 16652
rect 10772 16643 10830 16649
rect 10772 16609 10784 16643
rect 10818 16640 10830 16643
rect 11790 16640 11796 16652
rect 10818 16612 11796 16640
rect 10818 16609 10830 16612
rect 10772 16603 10830 16609
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 11974 16600 11980 16652
rect 12032 16640 12038 16652
rect 12084 16640 12112 16680
rect 12710 16668 12716 16680
rect 12768 16708 12774 16720
rect 13256 16711 13314 16717
rect 12768 16680 13216 16708
rect 12768 16668 12774 16680
rect 12032 16612 12112 16640
rect 12253 16643 12311 16649
rect 12032 16600 12038 16612
rect 12253 16609 12265 16643
rect 12299 16640 12311 16643
rect 12434 16640 12440 16652
rect 12299 16612 12440 16640
rect 12299 16609 12311 16612
rect 12253 16603 12311 16609
rect 12434 16600 12440 16612
rect 12492 16600 12498 16652
rect 12529 16643 12587 16649
rect 12529 16609 12541 16643
rect 12575 16640 12587 16643
rect 13078 16640 13084 16652
rect 12575 16612 13084 16640
rect 12575 16609 12587 16612
rect 12529 16603 12587 16609
rect 13078 16600 13084 16612
rect 13136 16600 13142 16652
rect 13188 16640 13216 16680
rect 13256 16677 13268 16711
rect 13302 16708 13314 16711
rect 14274 16708 14280 16720
rect 13302 16680 14280 16708
rect 13302 16677 13314 16680
rect 13256 16671 13314 16677
rect 14274 16668 14280 16680
rect 14332 16668 14338 16720
rect 17236 16708 17264 16748
rect 14752 16680 17264 16708
rect 14645 16643 14703 16649
rect 14645 16640 14657 16643
rect 13188 16612 14657 16640
rect 14645 16609 14657 16612
rect 14691 16609 14703 16643
rect 14645 16603 14703 16609
rect 4663 16544 5212 16572
rect 5261 16575 5319 16581
rect 4663 16541 4675 16544
rect 4617 16535 4675 16541
rect 5261 16541 5273 16575
rect 5307 16541 5319 16575
rect 7466 16572 7472 16584
rect 5261 16535 5319 16541
rect 6564 16544 7328 16572
rect 7427 16544 7472 16572
rect 4522 16464 4528 16516
rect 4580 16464 4586 16516
rect 5074 16464 5080 16516
rect 5132 16504 5138 16516
rect 5276 16504 5304 16535
rect 5132 16476 5304 16504
rect 5132 16464 5138 16476
rect 3970 16396 3976 16448
rect 4028 16436 4034 16448
rect 4065 16439 4123 16445
rect 4065 16436 4077 16439
rect 4028 16408 4077 16436
rect 4028 16396 4034 16408
rect 4065 16405 4077 16408
rect 4111 16405 4123 16439
rect 4540 16436 4568 16464
rect 4890 16436 4896 16448
rect 4540 16408 4896 16436
rect 4065 16399 4123 16405
rect 4890 16396 4896 16408
rect 4948 16396 4954 16448
rect 5534 16396 5540 16448
rect 5592 16436 5598 16448
rect 6564 16436 6592 16544
rect 6914 16504 6920 16516
rect 6875 16476 6920 16504
rect 6914 16464 6920 16476
rect 6972 16464 6978 16516
rect 5592 16408 6592 16436
rect 6641 16439 6699 16445
rect 5592 16396 5598 16408
rect 6641 16405 6653 16439
rect 6687 16436 6699 16439
rect 7190 16436 7196 16448
rect 6687 16408 7196 16436
rect 6687 16405 6699 16408
rect 6641 16399 6699 16405
rect 7190 16396 7196 16408
rect 7248 16396 7254 16448
rect 7300 16436 7328 16544
rect 7466 16532 7472 16544
rect 7524 16532 7530 16584
rect 7742 16532 7748 16584
rect 7800 16572 7806 16584
rect 7929 16575 7987 16581
rect 7929 16572 7941 16575
rect 7800 16544 7941 16572
rect 7800 16532 7806 16544
rect 7929 16541 7941 16544
rect 7975 16541 7987 16575
rect 10502 16572 10508 16584
rect 10463 16544 10508 16572
rect 7929 16535 7987 16541
rect 10502 16532 10508 16544
rect 10560 16532 10566 16584
rect 12066 16532 12072 16584
rect 12124 16572 12130 16584
rect 12989 16575 13047 16581
rect 12989 16572 13001 16575
rect 12124 16544 13001 16572
rect 12124 16532 12130 16544
rect 12989 16541 13001 16544
rect 13035 16541 13047 16575
rect 12989 16535 13047 16541
rect 10686 16436 10692 16448
rect 7300 16408 10692 16436
rect 10686 16396 10692 16408
rect 10744 16436 10750 16448
rect 12526 16436 12532 16448
rect 10744 16408 12532 16436
rect 10744 16396 10750 16408
rect 12526 16396 12532 16408
rect 12584 16396 12590 16448
rect 13004 16436 13032 16535
rect 14090 16532 14096 16584
rect 14148 16572 14154 16584
rect 14752 16572 14780 16680
rect 17310 16668 17316 16720
rect 17368 16668 17374 16720
rect 17420 16708 17448 16748
rect 17586 16736 17592 16748
rect 17644 16736 17650 16788
rect 18969 16779 19027 16785
rect 18969 16745 18981 16779
rect 19015 16776 19027 16779
rect 19242 16776 19248 16788
rect 19015 16748 19248 16776
rect 19015 16745 19027 16748
rect 18969 16739 19027 16745
rect 19242 16736 19248 16748
rect 19300 16776 19306 16788
rect 19610 16776 19616 16788
rect 19300 16748 19616 16776
rect 19300 16736 19306 16748
rect 19610 16736 19616 16748
rect 19668 16736 19674 16788
rect 19981 16779 20039 16785
rect 19981 16745 19993 16779
rect 20027 16776 20039 16779
rect 20162 16776 20168 16788
rect 20027 16748 20168 16776
rect 20027 16745 20039 16748
rect 19981 16739 20039 16745
rect 20162 16736 20168 16748
rect 20220 16736 20226 16788
rect 18049 16711 18107 16717
rect 18049 16708 18061 16711
rect 17420 16680 18061 16708
rect 18049 16677 18061 16680
rect 18095 16677 18107 16711
rect 20073 16711 20131 16717
rect 20073 16708 20085 16711
rect 18049 16671 18107 16677
rect 18156 16680 20085 16708
rect 15013 16643 15071 16649
rect 15013 16609 15025 16643
rect 15059 16609 15071 16643
rect 15013 16603 15071 16609
rect 14148 16544 14780 16572
rect 15028 16572 15056 16603
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 15470 16640 15476 16652
rect 15252 16612 15476 16640
rect 15252 16600 15258 16612
rect 15470 16600 15476 16612
rect 15528 16640 15534 16652
rect 17328 16640 17356 16668
rect 17957 16643 18015 16649
rect 17957 16640 17969 16643
rect 15528 16612 17264 16640
rect 17328 16612 17969 16640
rect 15528 16600 15534 16612
rect 16022 16572 16028 16584
rect 15028 16544 16028 16572
rect 14148 16532 14154 16544
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 16209 16575 16267 16581
rect 16209 16541 16221 16575
rect 16255 16572 16267 16575
rect 16390 16572 16396 16584
rect 16255 16544 16396 16572
rect 16255 16541 16267 16544
rect 16209 16535 16267 16541
rect 13998 16464 14004 16516
rect 14056 16504 14062 16516
rect 16224 16504 16252 16535
rect 16390 16532 16396 16544
rect 16448 16532 16454 16584
rect 17236 16581 17264 16612
rect 17957 16609 17969 16612
rect 18003 16609 18015 16643
rect 17957 16603 18015 16609
rect 17037 16575 17095 16581
rect 17037 16541 17049 16575
rect 17083 16541 17095 16575
rect 17037 16535 17095 16541
rect 17221 16575 17279 16581
rect 17221 16541 17233 16575
rect 17267 16541 17279 16575
rect 17221 16535 17279 16541
rect 14056 16476 16252 16504
rect 14056 16464 14062 16476
rect 16574 16464 16580 16516
rect 16632 16504 16638 16516
rect 16850 16504 16856 16516
rect 16632 16476 16856 16504
rect 16632 16464 16638 16476
rect 16850 16464 16856 16476
rect 16908 16464 16914 16516
rect 13630 16436 13636 16448
rect 13004 16408 13636 16436
rect 13630 16396 13636 16408
rect 13688 16396 13694 16448
rect 15838 16396 15844 16448
rect 15896 16436 15902 16448
rect 17052 16436 17080 16535
rect 17770 16532 17776 16584
rect 17828 16572 17834 16584
rect 18156 16572 18184 16680
rect 20073 16677 20085 16680
rect 20119 16677 20131 16711
rect 20073 16671 20131 16677
rect 18322 16600 18328 16652
rect 18380 16640 18386 16652
rect 19061 16643 19119 16649
rect 19061 16640 19073 16643
rect 18380 16612 19073 16640
rect 18380 16600 18386 16612
rect 19061 16609 19073 16612
rect 19107 16609 19119 16643
rect 20901 16643 20959 16649
rect 20901 16640 20913 16643
rect 19061 16603 19119 16609
rect 19352 16612 20913 16640
rect 17828 16544 18184 16572
rect 18233 16575 18291 16581
rect 17828 16532 17834 16544
rect 18233 16541 18245 16575
rect 18279 16572 18291 16575
rect 19153 16575 19211 16581
rect 19153 16572 19165 16575
rect 18279 16544 19165 16572
rect 18279 16541 18291 16544
rect 18233 16535 18291 16541
rect 19153 16541 19165 16544
rect 19199 16541 19211 16575
rect 19153 16535 19211 16541
rect 17862 16464 17868 16516
rect 17920 16504 17926 16516
rect 18248 16504 18276 16535
rect 19242 16532 19248 16584
rect 19300 16572 19306 16584
rect 19352 16572 19380 16612
rect 20901 16609 20913 16612
rect 20947 16609 20959 16643
rect 20901 16603 20959 16609
rect 19300 16544 19380 16572
rect 20165 16575 20223 16581
rect 19300 16532 19306 16544
rect 20165 16541 20177 16575
rect 20211 16541 20223 16575
rect 20165 16535 20223 16541
rect 17920 16476 18276 16504
rect 17920 16464 17926 16476
rect 18414 16464 18420 16516
rect 18472 16464 18478 16516
rect 18598 16504 18604 16516
rect 18559 16476 18604 16504
rect 18598 16464 18604 16476
rect 18656 16464 18662 16516
rect 18782 16464 18788 16516
rect 18840 16504 18846 16516
rect 20180 16504 20208 16535
rect 18840 16476 20208 16504
rect 18840 16464 18846 16476
rect 15896 16408 17080 16436
rect 15896 16396 15902 16408
rect 17586 16396 17592 16448
rect 17644 16436 17650 16448
rect 18432 16436 18460 16464
rect 19610 16436 19616 16448
rect 17644 16408 18460 16436
rect 19571 16408 19616 16436
rect 17644 16396 17650 16408
rect 19610 16396 19616 16408
rect 19668 16396 19674 16448
rect 20162 16396 20168 16448
rect 20220 16436 20226 16448
rect 20622 16436 20628 16448
rect 20220 16408 20628 16436
rect 20220 16396 20226 16408
rect 20622 16396 20628 16408
rect 20680 16396 20686 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 1486 16192 1492 16244
rect 1544 16232 1550 16244
rect 1581 16235 1639 16241
rect 1581 16232 1593 16235
rect 1544 16204 1593 16232
rect 1544 16192 1550 16204
rect 1581 16201 1593 16204
rect 1627 16201 1639 16235
rect 2590 16232 2596 16244
rect 2551 16204 2596 16232
rect 1581 16195 1639 16201
rect 2590 16192 2596 16204
rect 2648 16192 2654 16244
rect 3789 16235 3847 16241
rect 3789 16201 3801 16235
rect 3835 16232 3847 16235
rect 5442 16232 5448 16244
rect 3835 16204 5448 16232
rect 3835 16201 3847 16204
rect 3789 16195 3847 16201
rect 5442 16192 5448 16204
rect 5500 16192 5506 16244
rect 6641 16235 6699 16241
rect 6641 16201 6653 16235
rect 6687 16232 6699 16235
rect 7742 16232 7748 16244
rect 6687 16204 7748 16232
rect 6687 16201 6699 16204
rect 6641 16195 6699 16201
rect 7742 16192 7748 16204
rect 7800 16192 7806 16244
rect 8846 16192 8852 16244
rect 8904 16232 8910 16244
rect 12437 16235 12495 16241
rect 8904 16204 9352 16232
rect 8904 16192 8910 16204
rect 4614 16164 4620 16176
rect 4448 16136 4620 16164
rect 2682 16056 2688 16108
rect 2740 16096 2746 16108
rect 3145 16099 3203 16105
rect 3145 16096 3157 16099
rect 2740 16068 3157 16096
rect 2740 16056 2746 16068
rect 3145 16065 3157 16068
rect 3191 16065 3203 16099
rect 3145 16059 3203 16065
rect 3970 16056 3976 16108
rect 4028 16056 4034 16108
rect 4246 16096 4252 16108
rect 4207 16068 4252 16096
rect 4246 16056 4252 16068
rect 4304 16056 4310 16108
rect 4448 16105 4476 16136
rect 4614 16124 4620 16136
rect 4672 16124 4678 16176
rect 6178 16164 6184 16176
rect 5828 16136 6184 16164
rect 4433 16099 4491 16105
rect 4433 16065 4445 16099
rect 4479 16065 4491 16099
rect 4433 16059 4491 16065
rect 4798 16056 4804 16108
rect 4856 16096 4862 16108
rect 5828 16105 5856 16136
rect 6178 16124 6184 16136
rect 6236 16124 6242 16176
rect 9033 16167 9091 16173
rect 9033 16164 9045 16167
rect 8680 16136 9045 16164
rect 5813 16099 5871 16105
rect 4856 16068 4901 16096
rect 4856 16056 4862 16068
rect 5813 16065 5825 16099
rect 5859 16065 5871 16099
rect 5813 16059 5871 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1670 16028 1676 16040
rect 1443 16000 1676 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1670 15988 1676 16000
rect 1728 15988 1734 16040
rect 1857 16031 1915 16037
rect 1857 15997 1869 16031
rect 1903 16028 1915 16031
rect 2038 16028 2044 16040
rect 1903 16000 2044 16028
rect 1903 15997 1915 16000
rect 1857 15991 1915 15997
rect 2038 15988 2044 16000
rect 2096 15988 2102 16040
rect 2130 15988 2136 16040
rect 2188 16028 2194 16040
rect 2188 16000 2233 16028
rect 2188 15988 2194 16000
rect 2774 15988 2780 16040
rect 2832 16028 2838 16040
rect 3053 16031 3111 16037
rect 3053 16028 3065 16031
rect 2832 16000 3065 16028
rect 2832 15988 2838 16000
rect 3053 15997 3065 16000
rect 3099 15997 3111 16031
rect 3988 16028 4016 16056
rect 8680 16037 8708 16136
rect 9033 16133 9045 16136
rect 9079 16133 9091 16167
rect 9324 16164 9352 16204
rect 10435 16204 12388 16232
rect 9401 16167 9459 16173
rect 9401 16164 9413 16167
rect 9324 16136 9413 16164
rect 9033 16127 9091 16133
rect 9401 16133 9413 16136
rect 9447 16133 9459 16167
rect 10435 16164 10463 16204
rect 9401 16127 9459 16133
rect 9508 16136 10463 16164
rect 8754 16056 8760 16108
rect 8812 16096 8818 16108
rect 9306 16096 9312 16108
rect 8812 16068 9312 16096
rect 8812 16056 8818 16068
rect 9306 16056 9312 16068
rect 9364 16056 9370 16108
rect 4157 16031 4215 16037
rect 4157 16028 4169 16031
rect 3988 16000 4169 16028
rect 3053 15991 3111 15997
rect 4157 15997 4169 16000
rect 4203 15997 4215 16031
rect 4157 15991 4215 15997
rect 6641 16031 6699 16037
rect 6641 15997 6653 16031
rect 6687 16028 6699 16031
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 6687 16000 6837 16028
rect 6687 15997 6699 16000
rect 6641 15991 6699 15997
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 6825 15991 6883 15997
rect 8665 16031 8723 16037
rect 8665 15997 8677 16031
rect 8711 15997 8723 16031
rect 8665 15991 8723 15997
rect 8938 15988 8944 16040
rect 8996 16028 9002 16040
rect 9508 16028 9536 16136
rect 9582 16056 9588 16108
rect 9640 16096 9646 16108
rect 9953 16099 10011 16105
rect 9953 16096 9965 16099
rect 9640 16068 9965 16096
rect 9640 16056 9646 16068
rect 9953 16065 9965 16068
rect 9999 16065 10011 16099
rect 9953 16059 10011 16065
rect 8996 16000 9536 16028
rect 10413 16031 10471 16037
rect 8996 15988 9002 16000
rect 10413 15997 10425 16031
rect 10459 16028 10471 16031
rect 10502 16028 10508 16040
rect 10459 16000 10508 16028
rect 10459 15997 10471 16000
rect 10413 15991 10471 15997
rect 10502 15988 10508 16000
rect 10560 15988 10566 16040
rect 12360 16028 12388 16204
rect 12437 16201 12449 16235
rect 12483 16232 12495 16235
rect 12894 16232 12900 16244
rect 12483 16204 12900 16232
rect 12483 16201 12495 16204
rect 12437 16195 12495 16201
rect 12894 16192 12900 16204
rect 12952 16192 12958 16244
rect 12986 16192 12992 16244
rect 13044 16232 13050 16244
rect 13449 16235 13507 16241
rect 13449 16232 13461 16235
rect 13044 16204 13461 16232
rect 13044 16192 13050 16204
rect 13449 16201 13461 16204
rect 13495 16201 13507 16235
rect 13449 16195 13507 16201
rect 14182 16192 14188 16244
rect 14240 16232 14246 16244
rect 15102 16232 15108 16244
rect 14240 16204 15108 16232
rect 14240 16192 14246 16204
rect 15102 16192 15108 16204
rect 15160 16192 15166 16244
rect 15838 16232 15844 16244
rect 15799 16204 15844 16232
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 17954 16192 17960 16244
rect 18012 16232 18018 16244
rect 18233 16235 18291 16241
rect 18233 16232 18245 16235
rect 18012 16204 18245 16232
rect 18012 16192 18018 16204
rect 18233 16201 18245 16204
rect 18279 16201 18291 16235
rect 18233 16195 18291 16201
rect 18506 16192 18512 16244
rect 18564 16232 18570 16244
rect 18782 16232 18788 16244
rect 18564 16204 18788 16232
rect 18564 16192 18570 16204
rect 18782 16192 18788 16204
rect 18840 16192 18846 16244
rect 14829 16167 14887 16173
rect 14829 16133 14841 16167
rect 14875 16133 14887 16167
rect 14829 16127 14887 16133
rect 16132 16136 16528 16164
rect 13081 16099 13139 16105
rect 13081 16065 13093 16099
rect 13127 16096 13139 16099
rect 13262 16096 13268 16108
rect 13127 16068 13268 16096
rect 13127 16065 13139 16068
rect 13081 16059 13139 16065
rect 13262 16056 13268 16068
rect 13320 16096 13326 16108
rect 14001 16099 14059 16105
rect 14001 16096 14013 16099
rect 13320 16068 14013 16096
rect 13320 16056 13326 16068
rect 14001 16065 14013 16068
rect 14047 16065 14059 16099
rect 14001 16059 14059 16065
rect 13909 16031 13967 16037
rect 13909 16028 13921 16031
rect 12360 16000 13921 16028
rect 13909 15997 13921 16000
rect 13955 15997 13967 16031
rect 14844 16028 14872 16127
rect 15102 16056 15108 16108
rect 15160 16096 15166 16108
rect 15289 16099 15347 16105
rect 15289 16096 15301 16099
rect 15160 16068 15301 16096
rect 15160 16056 15166 16068
rect 15289 16065 15301 16068
rect 15335 16065 15347 16099
rect 15470 16096 15476 16108
rect 15431 16068 15476 16096
rect 15289 16059 15347 16065
rect 15470 16056 15476 16068
rect 15528 16056 15534 16108
rect 15197 16031 15255 16037
rect 14844 16000 15148 16028
rect 13909 15991 13967 15997
rect 4614 15920 4620 15972
rect 4672 15960 4678 15972
rect 5534 15960 5540 15972
rect 4672 15932 5540 15960
rect 4672 15920 4678 15932
rect 5534 15920 5540 15932
rect 5592 15920 5598 15972
rect 5721 15963 5779 15969
rect 5721 15929 5733 15963
rect 5767 15960 5779 15963
rect 6914 15960 6920 15972
rect 5767 15932 6920 15960
rect 5767 15929 5779 15932
rect 5721 15923 5779 15929
rect 6914 15920 6920 15932
rect 6972 15920 6978 15972
rect 7092 15963 7150 15969
rect 7092 15929 7104 15963
rect 7138 15960 7150 15963
rect 7190 15960 7196 15972
rect 7138 15932 7196 15960
rect 7138 15929 7150 15932
rect 7092 15923 7150 15929
rect 7190 15920 7196 15932
rect 7248 15960 7254 15972
rect 9122 15960 9128 15972
rect 7248 15932 9128 15960
rect 7248 15920 7254 15932
rect 9122 15920 9128 15932
rect 9180 15920 9186 15972
rect 9309 15963 9367 15969
rect 9309 15929 9321 15963
rect 9355 15960 9367 15963
rect 9861 15963 9919 15969
rect 9861 15960 9873 15963
rect 9355 15932 9873 15960
rect 9355 15929 9367 15932
rect 9309 15923 9367 15929
rect 9861 15929 9873 15932
rect 9907 15960 9919 15963
rect 10042 15960 10048 15972
rect 9907 15932 10048 15960
rect 9907 15929 9919 15932
rect 9861 15923 9919 15929
rect 10042 15920 10048 15932
rect 10100 15920 10106 15972
rect 10680 15963 10738 15969
rect 10680 15929 10692 15963
rect 10726 15960 10738 15963
rect 11606 15960 11612 15972
rect 10726 15932 11612 15960
rect 10726 15929 10738 15932
rect 10680 15923 10738 15929
rect 11606 15920 11612 15932
rect 11664 15920 11670 15972
rect 12805 15963 12863 15969
rect 12805 15929 12817 15963
rect 12851 15960 12863 15963
rect 13262 15960 13268 15972
rect 12851 15932 13268 15960
rect 12851 15929 12863 15932
rect 12805 15923 12863 15929
rect 13262 15920 13268 15932
rect 13320 15920 13326 15972
rect 2406 15852 2412 15904
rect 2464 15892 2470 15904
rect 2961 15895 3019 15901
rect 2961 15892 2973 15895
rect 2464 15864 2973 15892
rect 2464 15852 2470 15864
rect 2961 15861 2973 15864
rect 3007 15861 3019 15895
rect 2961 15855 3019 15861
rect 4706 15852 4712 15904
rect 4764 15892 4770 15904
rect 5261 15895 5319 15901
rect 5261 15892 5273 15895
rect 4764 15864 5273 15892
rect 4764 15852 4770 15864
rect 5261 15861 5273 15864
rect 5307 15861 5319 15895
rect 5626 15892 5632 15904
rect 5587 15864 5632 15892
rect 5261 15855 5319 15861
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 6270 15892 6276 15904
rect 6231 15864 6276 15892
rect 6270 15852 6276 15864
rect 6328 15852 6334 15904
rect 6362 15852 6368 15904
rect 6420 15892 6426 15904
rect 7282 15892 7288 15904
rect 6420 15864 7288 15892
rect 6420 15852 6426 15864
rect 7282 15852 7288 15864
rect 7340 15892 7346 15904
rect 7466 15892 7472 15904
rect 7340 15864 7472 15892
rect 7340 15852 7346 15864
rect 7466 15852 7472 15864
rect 7524 15892 7530 15904
rect 8205 15895 8263 15901
rect 8205 15892 8217 15895
rect 7524 15864 8217 15892
rect 7524 15852 7530 15864
rect 8205 15861 8217 15864
rect 8251 15861 8263 15895
rect 8846 15892 8852 15904
rect 8807 15864 8852 15892
rect 8205 15855 8263 15861
rect 8846 15852 8852 15864
rect 8904 15852 8910 15904
rect 9033 15895 9091 15901
rect 9033 15861 9045 15895
rect 9079 15892 9091 15895
rect 9674 15892 9680 15904
rect 9079 15864 9680 15892
rect 9079 15861 9091 15864
rect 9033 15855 9091 15861
rect 9674 15852 9680 15864
rect 9732 15852 9738 15904
rect 9769 15895 9827 15901
rect 9769 15861 9781 15895
rect 9815 15892 9827 15895
rect 10962 15892 10968 15904
rect 9815 15864 10968 15892
rect 9815 15861 9827 15864
rect 9769 15855 9827 15861
rect 10962 15852 10968 15864
rect 11020 15852 11026 15904
rect 11790 15892 11796 15904
rect 11703 15864 11796 15892
rect 11790 15852 11796 15864
rect 11848 15892 11854 15904
rect 12710 15892 12716 15904
rect 11848 15864 12716 15892
rect 11848 15852 11854 15864
rect 12710 15852 12716 15864
rect 12768 15852 12774 15904
rect 12894 15892 12900 15904
rect 12855 15864 12900 15892
rect 12894 15852 12900 15864
rect 12952 15852 12958 15904
rect 13814 15892 13820 15904
rect 13775 15864 13820 15892
rect 13814 15852 13820 15864
rect 13872 15852 13878 15904
rect 13924 15892 13952 15991
rect 15120 15960 15148 16000
rect 15197 15997 15209 16031
rect 15243 16028 15255 16031
rect 16132 16028 16160 16136
rect 16390 16096 16396 16108
rect 16351 16068 16396 16096
rect 16390 16056 16396 16068
rect 16448 16056 16454 16108
rect 15243 16000 16160 16028
rect 15243 15997 15255 16000
rect 15197 15991 15255 15997
rect 16206 15988 16212 16040
rect 16264 16028 16270 16040
rect 16301 16031 16359 16037
rect 16301 16028 16313 16031
rect 16264 16000 16313 16028
rect 16264 15988 16270 16000
rect 16301 15997 16313 16000
rect 16347 15997 16359 16031
rect 16500 16028 16528 16136
rect 16758 16124 16764 16176
rect 16816 16164 16822 16176
rect 16853 16167 16911 16173
rect 16853 16164 16865 16167
rect 16816 16136 16865 16164
rect 16816 16124 16822 16136
rect 16853 16133 16865 16136
rect 16899 16133 16911 16167
rect 16853 16127 16911 16133
rect 17126 16124 17132 16176
rect 17184 16164 17190 16176
rect 17184 16136 18828 16164
rect 17184 16124 17190 16136
rect 16942 16056 16948 16108
rect 17000 16096 17006 16108
rect 17405 16099 17463 16105
rect 17405 16096 17417 16099
rect 17000 16068 17417 16096
rect 17000 16056 17006 16068
rect 17405 16065 17417 16068
rect 17451 16065 17463 16099
rect 17405 16059 17463 16065
rect 17678 16056 17684 16108
rect 17736 16096 17742 16108
rect 18800 16105 18828 16136
rect 18966 16124 18972 16176
rect 19024 16164 19030 16176
rect 20438 16164 20444 16176
rect 19024 16136 20444 16164
rect 19024 16124 19030 16136
rect 20438 16124 20444 16136
rect 20496 16124 20502 16176
rect 18693 16099 18751 16105
rect 18693 16096 18705 16099
rect 17736 16068 18705 16096
rect 17736 16056 17742 16068
rect 18693 16065 18705 16068
rect 18739 16065 18751 16099
rect 18693 16059 18751 16065
rect 18785 16099 18843 16105
rect 18785 16065 18797 16099
rect 18831 16065 18843 16099
rect 19702 16096 19708 16108
rect 19663 16068 19708 16096
rect 18785 16059 18843 16065
rect 19702 16056 19708 16068
rect 19760 16056 19766 16108
rect 20622 16096 20628 16108
rect 20583 16068 20628 16096
rect 20622 16056 20628 16068
rect 20680 16056 20686 16108
rect 19242 16028 19248 16040
rect 16500 16000 19248 16028
rect 16301 15991 16359 15997
rect 19242 15988 19248 16000
rect 19300 15988 19306 16040
rect 17221 15963 17279 15969
rect 17221 15960 17233 15963
rect 15120 15932 17233 15960
rect 17221 15929 17233 15932
rect 17267 15929 17279 15963
rect 20441 15963 20499 15969
rect 20441 15960 20453 15963
rect 17221 15923 17279 15929
rect 19076 15932 20453 15960
rect 16022 15892 16028 15904
rect 13924 15864 16028 15892
rect 16022 15852 16028 15864
rect 16080 15852 16086 15904
rect 16114 15852 16120 15904
rect 16172 15892 16178 15904
rect 16209 15895 16267 15901
rect 16209 15892 16221 15895
rect 16172 15864 16221 15892
rect 16172 15852 16178 15864
rect 16209 15861 16221 15864
rect 16255 15861 16267 15895
rect 16209 15855 16267 15861
rect 16298 15852 16304 15904
rect 16356 15892 16362 15904
rect 17126 15892 17132 15904
rect 16356 15864 17132 15892
rect 16356 15852 16362 15864
rect 17126 15852 17132 15864
rect 17184 15852 17190 15904
rect 17310 15892 17316 15904
rect 17271 15864 17316 15892
rect 17310 15852 17316 15864
rect 17368 15852 17374 15904
rect 18598 15892 18604 15904
rect 18559 15864 18604 15892
rect 18598 15852 18604 15864
rect 18656 15852 18662 15904
rect 19076 15901 19104 15932
rect 20441 15929 20453 15932
rect 20487 15929 20499 15963
rect 20441 15923 20499 15929
rect 19061 15895 19119 15901
rect 19061 15861 19073 15895
rect 19107 15861 19119 15895
rect 19426 15892 19432 15904
rect 19387 15864 19432 15892
rect 19061 15855 19119 15861
rect 19426 15852 19432 15864
rect 19484 15852 19490 15904
rect 19518 15852 19524 15904
rect 19576 15892 19582 15904
rect 19576 15864 19621 15892
rect 19576 15852 19582 15864
rect 19978 15852 19984 15904
rect 20036 15892 20042 15904
rect 20073 15895 20131 15901
rect 20073 15892 20085 15895
rect 20036 15864 20085 15892
rect 20036 15852 20042 15864
rect 20073 15861 20085 15864
rect 20119 15861 20131 15895
rect 20530 15892 20536 15904
rect 20491 15864 20536 15892
rect 20073 15855 20131 15861
rect 20530 15852 20536 15864
rect 20588 15852 20594 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 2314 15688 2320 15700
rect 2275 15660 2320 15688
rect 2314 15648 2320 15660
rect 2372 15648 2378 15700
rect 4062 15648 4068 15700
rect 4120 15688 4126 15700
rect 6086 15688 6092 15700
rect 4120 15660 6092 15688
rect 4120 15648 4126 15660
rect 6086 15648 6092 15660
rect 6144 15648 6150 15700
rect 6270 15648 6276 15700
rect 6328 15688 6334 15700
rect 8941 15691 8999 15697
rect 8941 15688 8953 15691
rect 6328 15660 8953 15688
rect 6328 15648 6334 15660
rect 8941 15657 8953 15660
rect 8987 15657 8999 15691
rect 8941 15651 8999 15657
rect 9674 15648 9680 15700
rect 9732 15688 9738 15700
rect 10689 15691 10747 15697
rect 9732 15660 9777 15688
rect 9732 15648 9738 15660
rect 10689 15657 10701 15691
rect 10735 15688 10747 15691
rect 13814 15688 13820 15700
rect 10735 15660 13820 15688
rect 10735 15657 10747 15660
rect 10689 15651 10747 15657
rect 13814 15648 13820 15660
rect 13872 15648 13878 15700
rect 16298 15688 16304 15700
rect 14384 15660 16304 15688
rect 3421 15623 3479 15629
rect 3421 15589 3433 15623
rect 3467 15620 3479 15623
rect 4614 15620 4620 15632
rect 3467 15592 4620 15620
rect 3467 15589 3479 15592
rect 3421 15583 3479 15589
rect 4614 15580 4620 15592
rect 4672 15580 4678 15632
rect 4893 15623 4951 15629
rect 4893 15589 4905 15623
rect 4939 15620 4951 15623
rect 4939 15592 8524 15620
rect 4939 15589 4951 15592
rect 4893 15583 4951 15589
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15521 1455 15555
rect 1397 15515 1455 15521
rect 1412 15416 1440 15515
rect 2222 15512 2228 15564
rect 2280 15552 2286 15564
rect 2590 15552 2596 15564
rect 2280 15524 2596 15552
rect 2280 15512 2286 15524
rect 1486 15444 1492 15496
rect 1544 15484 1550 15496
rect 2516 15493 2544 15524
rect 2590 15512 2596 15524
rect 2648 15512 2654 15564
rect 3329 15555 3387 15561
rect 3329 15521 3341 15555
rect 3375 15552 3387 15555
rect 4798 15552 4804 15564
rect 3375 15524 4804 15552
rect 3375 15521 3387 15524
rect 3329 15515 3387 15521
rect 4798 15512 4804 15524
rect 4856 15512 4862 15564
rect 4985 15555 5043 15561
rect 4985 15521 4997 15555
rect 5031 15552 5043 15555
rect 5442 15552 5448 15564
rect 5031 15524 5448 15552
rect 5031 15521 5043 15524
rect 4985 15515 5043 15521
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 5905 15555 5963 15561
rect 5905 15521 5917 15555
rect 5951 15552 5963 15555
rect 6454 15552 6460 15564
rect 5951 15524 6460 15552
rect 5951 15521 5963 15524
rect 5905 15515 5963 15521
rect 6454 15512 6460 15524
rect 6512 15512 6518 15564
rect 7190 15561 7196 15564
rect 6733 15555 6791 15561
rect 6733 15552 6745 15555
rect 6656 15524 6745 15552
rect 2409 15487 2467 15493
rect 2409 15484 2421 15487
rect 1544 15456 2421 15484
rect 1544 15444 1550 15456
rect 2409 15453 2421 15456
rect 2455 15453 2467 15487
rect 2409 15447 2467 15453
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15453 2559 15487
rect 2501 15447 2559 15453
rect 2774 15444 2780 15496
rect 2832 15484 2838 15496
rect 3513 15487 3571 15493
rect 3513 15484 3525 15487
rect 2832 15456 3525 15484
rect 2832 15444 2838 15456
rect 3513 15453 3525 15456
rect 3559 15453 3571 15487
rect 3513 15447 3571 15453
rect 3786 15444 3792 15496
rect 3844 15484 3850 15496
rect 4065 15487 4123 15493
rect 4065 15484 4077 15487
rect 3844 15456 4077 15484
rect 3844 15444 3850 15456
rect 4065 15453 4077 15456
rect 4111 15453 4123 15487
rect 4065 15447 4123 15453
rect 5169 15487 5227 15493
rect 5169 15453 5181 15487
rect 5215 15453 5227 15487
rect 5994 15484 6000 15496
rect 5955 15456 6000 15484
rect 5169 15447 5227 15453
rect 4890 15416 4896 15428
rect 1412 15388 4896 15416
rect 4890 15376 4896 15388
rect 4948 15376 4954 15428
rect 5184 15416 5212 15447
rect 5994 15444 6000 15456
rect 6052 15444 6058 15496
rect 6178 15484 6184 15496
rect 6139 15456 6184 15484
rect 6178 15444 6184 15456
rect 6236 15444 6242 15496
rect 6270 15416 6276 15428
rect 5184 15388 6276 15416
rect 6270 15376 6276 15388
rect 6328 15376 6334 15428
rect 6656 15360 6684 15524
rect 6733 15521 6745 15524
rect 6779 15521 6791 15555
rect 6733 15515 6791 15521
rect 7184 15515 7196 15561
rect 7248 15552 7254 15564
rect 7248 15524 7284 15552
rect 7190 15512 7196 15515
rect 7248 15512 7254 15524
rect 7466 15512 7472 15564
rect 7524 15552 7530 15564
rect 7524 15524 8432 15552
rect 7524 15512 7530 15524
rect 6917 15487 6975 15493
rect 6917 15453 6929 15487
rect 6963 15453 6975 15487
rect 6917 15447 6975 15453
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 1949 15351 2007 15357
rect 1949 15317 1961 15351
rect 1995 15348 2007 15351
rect 2406 15348 2412 15360
rect 1995 15320 2412 15348
rect 1995 15317 2007 15320
rect 1949 15311 2007 15317
rect 2406 15308 2412 15320
rect 2464 15308 2470 15360
rect 2958 15348 2964 15360
rect 2919 15320 2964 15348
rect 2958 15308 2964 15320
rect 3016 15308 3022 15360
rect 4525 15351 4583 15357
rect 4525 15317 4537 15351
rect 4571 15348 4583 15351
rect 5258 15348 5264 15360
rect 4571 15320 5264 15348
rect 4571 15317 4583 15320
rect 4525 15311 4583 15317
rect 5258 15308 5264 15320
rect 5316 15308 5322 15360
rect 5534 15348 5540 15360
rect 5495 15320 5540 15348
rect 5534 15308 5540 15320
rect 5592 15308 5598 15360
rect 6362 15308 6368 15360
rect 6420 15348 6426 15360
rect 6549 15351 6607 15357
rect 6549 15348 6561 15351
rect 6420 15320 6561 15348
rect 6420 15308 6426 15320
rect 6549 15317 6561 15320
rect 6595 15317 6607 15351
rect 6549 15311 6607 15317
rect 6638 15308 6644 15360
rect 6696 15308 6702 15360
rect 6932 15348 6960 15447
rect 8294 15416 8300 15428
rect 8255 15388 8300 15416
rect 8294 15376 8300 15388
rect 8352 15376 8358 15428
rect 7834 15348 7840 15360
rect 6932 15320 7840 15348
rect 7834 15308 7840 15320
rect 7892 15348 7898 15360
rect 8110 15348 8116 15360
rect 7892 15320 8116 15348
rect 7892 15308 7898 15320
rect 8110 15308 8116 15320
rect 8168 15308 8174 15360
rect 8404 15348 8432 15524
rect 8496 15416 8524 15592
rect 10502 15580 10508 15632
rect 10560 15620 10566 15632
rect 12066 15620 12072 15632
rect 10560 15592 12072 15620
rect 10560 15580 10566 15592
rect 9033 15555 9091 15561
rect 9033 15521 9045 15555
rect 9079 15552 9091 15555
rect 9582 15552 9588 15564
rect 9079 15524 9588 15552
rect 9079 15521 9091 15524
rect 9033 15515 9091 15521
rect 9582 15512 9588 15524
rect 9640 15512 9646 15564
rect 10045 15555 10103 15561
rect 10045 15521 10057 15555
rect 10091 15552 10103 15555
rect 10686 15552 10692 15564
rect 10091 15524 10692 15552
rect 10091 15521 10103 15524
rect 10045 15515 10103 15521
rect 10686 15512 10692 15524
rect 10744 15512 10750 15564
rect 11164 15561 11192 15592
rect 12066 15580 12072 15592
rect 12124 15620 12130 15632
rect 12621 15623 12679 15629
rect 12124 15592 12572 15620
rect 12124 15580 12130 15592
rect 11149 15555 11207 15561
rect 11149 15521 11161 15555
rect 11195 15521 11207 15555
rect 11149 15515 11207 15521
rect 11416 15555 11474 15561
rect 11416 15521 11428 15555
rect 11462 15552 11474 15555
rect 12544 15552 12572 15592
rect 12621 15589 12633 15623
rect 12667 15620 12679 15623
rect 13072 15623 13130 15629
rect 13072 15620 13084 15623
rect 12667 15592 13084 15620
rect 12667 15589 12679 15592
rect 12621 15583 12679 15589
rect 13072 15589 13084 15592
rect 13118 15620 13130 15623
rect 13538 15620 13544 15632
rect 13118 15592 13544 15620
rect 13118 15589 13130 15592
rect 13072 15583 13130 15589
rect 13538 15580 13544 15592
rect 13596 15620 13602 15632
rect 14384 15620 14412 15660
rect 16298 15648 16304 15660
rect 16356 15648 16362 15700
rect 16393 15691 16451 15697
rect 16393 15657 16405 15691
rect 16439 15688 16451 15691
rect 18693 15691 18751 15697
rect 18693 15688 18705 15691
rect 16439 15660 18705 15688
rect 16439 15657 16451 15660
rect 16393 15651 16451 15657
rect 18693 15657 18705 15660
rect 18739 15657 18751 15691
rect 18693 15651 18751 15657
rect 19429 15691 19487 15697
rect 19429 15657 19441 15691
rect 19475 15657 19487 15691
rect 19429 15651 19487 15657
rect 17310 15620 17316 15632
rect 13596 15592 14412 15620
rect 15120 15592 17316 15620
rect 13596 15580 13602 15592
rect 12805 15555 12863 15561
rect 12805 15552 12817 15555
rect 11462 15524 12487 15552
rect 12544 15524 12817 15552
rect 11462 15521 11474 15524
rect 11416 15515 11474 15521
rect 9122 15484 9128 15496
rect 9083 15456 9128 15484
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 9950 15444 9956 15496
rect 10008 15484 10014 15496
rect 10137 15487 10195 15493
rect 10137 15484 10149 15487
rect 10008 15456 10149 15484
rect 10008 15444 10014 15456
rect 10137 15453 10149 15456
rect 10183 15453 10195 15487
rect 10137 15447 10195 15453
rect 10229 15487 10287 15493
rect 10229 15453 10241 15487
rect 10275 15453 10287 15487
rect 12459 15484 12487 15524
rect 12805 15521 12817 15524
rect 12851 15521 12863 15555
rect 13630 15552 13636 15564
rect 12805 15515 12863 15521
rect 12912 15524 13636 15552
rect 12912 15484 12940 15524
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 14090 15512 14096 15564
rect 14148 15552 14154 15564
rect 14461 15555 14519 15561
rect 14461 15552 14473 15555
rect 14148 15524 14473 15552
rect 14148 15512 14154 15524
rect 14461 15521 14473 15524
rect 14507 15521 14519 15555
rect 14461 15515 14519 15521
rect 12459 15456 12940 15484
rect 10229 15447 10287 15453
rect 8573 15419 8631 15425
rect 8573 15416 8585 15419
rect 8496 15388 8585 15416
rect 8573 15385 8585 15388
rect 8619 15385 8631 15419
rect 8573 15379 8631 15385
rect 9490 15376 9496 15428
rect 9548 15416 9554 15428
rect 10244 15416 10272 15447
rect 14274 15444 14280 15496
rect 14332 15484 14338 15496
rect 14645 15487 14703 15493
rect 14645 15484 14657 15487
rect 14332 15456 14657 15484
rect 14332 15444 14338 15456
rect 14645 15453 14657 15456
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 9548 15388 10272 15416
rect 12529 15419 12587 15425
rect 9548 15376 9554 15388
rect 12529 15385 12541 15419
rect 12575 15416 12587 15419
rect 12621 15419 12679 15425
rect 12621 15416 12633 15419
rect 12575 15388 12633 15416
rect 12575 15385 12587 15388
rect 12529 15379 12587 15385
rect 12621 15385 12633 15388
rect 12667 15385 12679 15419
rect 15120 15416 15148 15592
rect 17310 15580 17316 15592
rect 17368 15580 17374 15632
rect 17773 15623 17831 15629
rect 17773 15589 17785 15623
rect 17819 15620 17831 15623
rect 18966 15620 18972 15632
rect 17819 15592 18972 15620
rect 17819 15589 17831 15592
rect 17773 15583 17831 15589
rect 18966 15580 18972 15592
rect 19024 15580 19030 15632
rect 19444 15620 19472 15651
rect 19610 15648 19616 15700
rect 19668 15688 19674 15700
rect 19889 15691 19947 15697
rect 19889 15688 19901 15691
rect 19668 15660 19901 15688
rect 19668 15648 19674 15660
rect 19889 15657 19901 15660
rect 19935 15657 19947 15691
rect 19889 15651 19947 15657
rect 20530 15620 20536 15632
rect 19444 15592 20536 15620
rect 20530 15580 20536 15592
rect 20588 15580 20594 15632
rect 15194 15512 15200 15564
rect 15252 15552 15258 15564
rect 15657 15555 15715 15561
rect 15657 15552 15669 15555
rect 15252 15524 15669 15552
rect 15252 15512 15258 15524
rect 15657 15521 15669 15524
rect 15703 15521 15715 15555
rect 16117 15555 16175 15561
rect 16117 15552 16129 15555
rect 15657 15515 15715 15521
rect 15764 15524 16129 15552
rect 15562 15444 15568 15496
rect 15620 15484 15626 15496
rect 15764 15493 15792 15524
rect 16117 15521 16129 15524
rect 16163 15521 16175 15555
rect 16758 15552 16764 15564
rect 16719 15524 16764 15552
rect 16117 15515 16175 15521
rect 16758 15512 16764 15524
rect 16816 15512 16822 15564
rect 17494 15552 17500 15564
rect 16960 15524 17500 15552
rect 15749 15487 15807 15493
rect 15749 15484 15761 15487
rect 15620 15456 15761 15484
rect 15620 15444 15626 15456
rect 15749 15453 15761 15456
rect 15795 15453 15807 15487
rect 15749 15447 15807 15453
rect 15841 15487 15899 15493
rect 15841 15453 15853 15487
rect 15887 15453 15899 15487
rect 16850 15484 16856 15496
rect 16811 15456 16856 15484
rect 15841 15447 15899 15453
rect 15289 15419 15347 15425
rect 15289 15416 15301 15419
rect 15120 15388 15301 15416
rect 12621 15379 12679 15385
rect 15289 15385 15301 15388
rect 15335 15385 15347 15419
rect 15289 15379 15347 15385
rect 15470 15376 15476 15428
rect 15528 15416 15534 15428
rect 15856 15416 15884 15447
rect 16850 15444 16856 15456
rect 16908 15444 16914 15496
rect 16666 15416 16672 15428
rect 15528 15388 15884 15416
rect 15948 15388 16672 15416
rect 15528 15376 15534 15388
rect 8754 15348 8760 15360
rect 8404 15320 8760 15348
rect 8754 15308 8760 15320
rect 8812 15348 8818 15360
rect 12250 15348 12256 15360
rect 8812 15320 12256 15348
rect 8812 15308 8818 15320
rect 12250 15308 12256 15320
rect 12308 15308 12314 15360
rect 14185 15351 14243 15357
rect 14185 15317 14197 15351
rect 14231 15348 14243 15351
rect 14642 15348 14648 15360
rect 14231 15320 14648 15348
rect 14231 15317 14243 15320
rect 14185 15311 14243 15317
rect 14642 15308 14648 15320
rect 14700 15348 14706 15360
rect 15948 15348 15976 15388
rect 16666 15376 16672 15388
rect 16724 15376 16730 15428
rect 14700 15320 15976 15348
rect 14700 15308 14706 15320
rect 16022 15308 16028 15360
rect 16080 15348 16086 15360
rect 16960 15348 16988 15524
rect 17494 15512 17500 15524
rect 17552 15552 17558 15564
rect 17865 15555 17923 15561
rect 17865 15552 17877 15555
rect 17552 15524 17877 15552
rect 17552 15512 17558 15524
rect 17865 15521 17877 15524
rect 17911 15552 17923 15555
rect 18598 15552 18604 15564
rect 17911 15524 18359 15552
rect 18559 15524 18604 15552
rect 17911 15521 17923 15524
rect 17865 15515 17923 15521
rect 17037 15487 17095 15493
rect 17037 15453 17049 15487
rect 17083 15484 17095 15487
rect 17310 15484 17316 15496
rect 17083 15456 17316 15484
rect 17083 15453 17095 15456
rect 17037 15447 17095 15453
rect 17310 15444 17316 15456
rect 17368 15444 17374 15496
rect 17954 15444 17960 15496
rect 18012 15484 18018 15496
rect 18331 15484 18359 15524
rect 18598 15512 18604 15524
rect 18656 15512 18662 15564
rect 19797 15555 19855 15561
rect 18708 15524 19104 15552
rect 18708 15484 18736 15524
rect 18874 15484 18880 15496
rect 18012 15456 18057 15484
rect 18331 15456 18736 15484
rect 18835 15456 18880 15484
rect 18012 15444 18018 15456
rect 18874 15444 18880 15456
rect 18932 15444 18938 15496
rect 19076 15484 19104 15524
rect 19797 15521 19809 15555
rect 19843 15552 19855 15555
rect 20438 15552 20444 15564
rect 19843 15524 20444 15552
rect 19843 15521 19855 15524
rect 19797 15515 19855 15521
rect 20438 15512 20444 15524
rect 20496 15512 20502 15564
rect 19076 15456 19196 15484
rect 17402 15348 17408 15360
rect 16080 15320 16988 15348
rect 17363 15320 17408 15348
rect 16080 15308 16086 15320
rect 17402 15308 17408 15320
rect 17460 15308 17466 15360
rect 17954 15308 17960 15360
rect 18012 15348 18018 15360
rect 18233 15351 18291 15357
rect 18233 15348 18245 15351
rect 18012 15320 18245 15348
rect 18012 15308 18018 15320
rect 18233 15317 18245 15320
rect 18279 15317 18291 15351
rect 19168 15348 19196 15456
rect 19610 15444 19616 15496
rect 19668 15484 19674 15496
rect 19981 15487 20039 15493
rect 19981 15484 19993 15487
rect 19668 15456 19993 15484
rect 19668 15444 19674 15456
rect 19981 15453 19993 15456
rect 20027 15453 20039 15487
rect 19981 15447 20039 15453
rect 21358 15348 21364 15360
rect 19168 15320 21364 15348
rect 18233 15311 18291 15317
rect 21358 15308 21364 15320
rect 21416 15308 21422 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 2406 15104 2412 15156
rect 2464 15144 2470 15156
rect 5258 15144 5264 15156
rect 2464 15116 5264 15144
rect 2464 15104 2470 15116
rect 5258 15104 5264 15116
rect 5316 15104 5322 15156
rect 5626 15104 5632 15156
rect 5684 15144 5690 15156
rect 6825 15147 6883 15153
rect 6825 15144 6837 15147
rect 5684 15116 6837 15144
rect 5684 15104 5690 15116
rect 6825 15113 6837 15116
rect 6871 15113 6883 15147
rect 6825 15107 6883 15113
rect 7190 15104 7196 15156
rect 7248 15144 7254 15156
rect 7248 15116 11560 15144
rect 7248 15104 7254 15116
rect 3053 15079 3111 15085
rect 3053 15045 3065 15079
rect 3099 15076 3111 15079
rect 3237 15079 3295 15085
rect 3237 15076 3249 15079
rect 3099 15048 3249 15076
rect 3099 15045 3111 15048
rect 3053 15039 3111 15045
rect 3237 15045 3249 15048
rect 3283 15045 3295 15079
rect 3237 15039 3295 15045
rect 6086 15036 6092 15088
rect 6144 15076 6150 15088
rect 8021 15079 8079 15085
rect 8021 15076 8033 15079
rect 6144 15048 8033 15076
rect 6144 15036 6150 15048
rect 8021 15045 8033 15048
rect 8067 15045 8079 15079
rect 8021 15039 8079 15045
rect 8110 15036 8116 15088
rect 8168 15076 8174 15088
rect 8389 15079 8447 15085
rect 8389 15076 8401 15079
rect 8168 15048 8401 15076
rect 8168 15036 8174 15048
rect 8389 15045 8401 15048
rect 8435 15076 8447 15079
rect 10045 15079 10103 15085
rect 8435 15048 8708 15076
rect 8435 15045 8447 15048
rect 8389 15039 8447 15045
rect 6454 14968 6460 15020
rect 6512 15008 6518 15020
rect 6638 15008 6644 15020
rect 6512 14980 6644 15008
rect 6512 14968 6518 14980
rect 6638 14968 6644 14980
rect 6696 14968 6702 15020
rect 8680 15017 8708 15048
rect 10045 15045 10057 15079
rect 10091 15076 10103 15079
rect 10229 15079 10287 15085
rect 10229 15076 10241 15079
rect 10091 15048 10241 15076
rect 10091 15045 10103 15048
rect 10045 15039 10103 15045
rect 10229 15045 10241 15048
rect 10275 15045 10287 15079
rect 11532 15076 11560 15116
rect 11606 15104 11612 15156
rect 11664 15144 11670 15156
rect 11701 15147 11759 15153
rect 11701 15144 11713 15147
rect 11664 15116 11713 15144
rect 11664 15104 11670 15116
rect 11701 15113 11713 15116
rect 11747 15113 11759 15147
rect 11701 15107 11759 15113
rect 12437 15147 12495 15153
rect 12437 15113 12449 15147
rect 12483 15144 12495 15147
rect 12802 15144 12808 15156
rect 12483 15116 12808 15144
rect 12483 15113 12495 15116
rect 12437 15107 12495 15113
rect 12802 15104 12808 15116
rect 12860 15104 12866 15156
rect 15010 15104 15016 15156
rect 15068 15144 15074 15156
rect 18785 15147 18843 15153
rect 18785 15144 18797 15147
rect 15068 15116 18797 15144
rect 15068 15104 15074 15116
rect 18785 15113 18797 15116
rect 18831 15113 18843 15147
rect 18785 15107 18843 15113
rect 18892 15116 19196 15144
rect 11532 15048 13115 15076
rect 10229 15039 10287 15045
rect 7469 15011 7527 15017
rect 7469 14977 7481 15011
rect 7515 14977 7527 15011
rect 7469 14971 7527 14977
rect 8665 15011 8723 15017
rect 8665 14977 8677 15011
rect 8711 14977 8723 15011
rect 8665 14971 8723 14977
rect 1673 14943 1731 14949
rect 1673 14909 1685 14943
rect 1719 14940 1731 14943
rect 1762 14940 1768 14952
rect 1719 14912 1768 14940
rect 1719 14909 1731 14912
rect 1673 14903 1731 14909
rect 1762 14900 1768 14912
rect 1820 14940 1826 14952
rect 2406 14940 2412 14952
rect 1820 14912 2412 14940
rect 1820 14900 1826 14912
rect 2406 14900 2412 14912
rect 2464 14940 2470 14952
rect 3329 14943 3387 14949
rect 3329 14940 3341 14943
rect 2464 14912 3341 14940
rect 2464 14900 2470 14912
rect 3329 14909 3341 14912
rect 3375 14940 3387 14943
rect 4985 14943 5043 14949
rect 4985 14940 4997 14943
rect 3375 14912 4997 14940
rect 3375 14909 3387 14912
rect 3329 14903 3387 14909
rect 4985 14909 4997 14912
rect 5031 14940 5043 14943
rect 5074 14940 5080 14952
rect 5031 14912 5080 14940
rect 5031 14909 5043 14912
rect 4985 14903 5043 14909
rect 5074 14900 5080 14912
rect 5132 14940 5138 14952
rect 6362 14940 6368 14952
rect 5132 14912 6368 14940
rect 5132 14900 5138 14912
rect 6362 14900 6368 14912
rect 6420 14900 6426 14952
rect 1940 14875 1998 14881
rect 1940 14841 1952 14875
rect 1986 14872 1998 14875
rect 2774 14872 2780 14884
rect 1986 14844 2780 14872
rect 1986 14841 1998 14844
rect 1940 14835 1998 14841
rect 2774 14832 2780 14844
rect 2832 14832 2838 14884
rect 3237 14875 3295 14881
rect 3237 14841 3249 14875
rect 3283 14872 3295 14875
rect 3510 14872 3516 14884
rect 3283 14844 3516 14872
rect 3283 14841 3295 14844
rect 3237 14835 3295 14841
rect 3510 14832 3516 14844
rect 3568 14881 3574 14884
rect 5258 14881 5264 14884
rect 3568 14875 3632 14881
rect 3568 14841 3586 14875
rect 3620 14841 3632 14875
rect 5252 14872 5264 14881
rect 3568 14835 3632 14841
rect 4540 14844 5120 14872
rect 5219 14844 5264 14872
rect 3568 14832 3574 14835
rect 2792 14804 2820 14832
rect 4540 14804 4568 14844
rect 2792 14776 4568 14804
rect 4614 14764 4620 14816
rect 4672 14804 4678 14816
rect 4709 14807 4767 14813
rect 4709 14804 4721 14807
rect 4672 14776 4721 14804
rect 4672 14764 4678 14776
rect 4709 14773 4721 14776
rect 4755 14773 4767 14807
rect 5092 14804 5120 14844
rect 5252 14835 5264 14844
rect 5258 14832 5264 14835
rect 5316 14832 5322 14884
rect 6270 14832 6276 14884
rect 6328 14872 6334 14884
rect 6656 14872 6684 14968
rect 7484 14940 7512 14971
rect 7742 14940 7748 14952
rect 7484 14912 7748 14940
rect 7742 14900 7748 14912
rect 7800 14900 7806 14952
rect 7837 14943 7895 14949
rect 7837 14909 7849 14943
rect 7883 14940 7895 14943
rect 7926 14940 7932 14952
rect 7883 14912 7932 14940
rect 7883 14909 7895 14912
rect 7837 14903 7895 14909
rect 7926 14900 7932 14912
rect 7984 14900 7990 14952
rect 8573 14943 8631 14949
rect 8573 14909 8585 14943
rect 8619 14909 8631 14943
rect 8680 14940 8708 14971
rect 12158 14968 12164 15020
rect 12216 15008 12222 15020
rect 12342 15008 12348 15020
rect 12216 14980 12348 15008
rect 12216 14968 12222 14980
rect 12342 14968 12348 14980
rect 12400 14968 12406 15020
rect 12710 14968 12716 15020
rect 12768 15008 12774 15020
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12768 14980 13001 15008
rect 12768 14968 12774 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 13087 15008 13115 15048
rect 17494 15036 17500 15088
rect 17552 15076 17558 15088
rect 18892 15076 18920 15116
rect 17552 15048 18920 15076
rect 19168 15076 19196 15116
rect 19426 15104 19432 15156
rect 19484 15144 19490 15156
rect 19484 15116 20760 15144
rect 19484 15104 19490 15116
rect 20073 15079 20131 15085
rect 20073 15076 20085 15079
rect 19168 15048 20085 15076
rect 17552 15036 17558 15048
rect 20073 15045 20085 15048
rect 20119 15045 20131 15079
rect 20073 15039 20131 15045
rect 14090 15008 14096 15020
rect 13087 14980 13952 15008
rect 14051 14980 14096 15008
rect 12989 14971 13047 14977
rect 10321 14943 10379 14949
rect 10321 14940 10333 14943
rect 8680 14912 10333 14940
rect 8573 14903 8631 14909
rect 10321 14909 10333 14912
rect 10367 14909 10379 14943
rect 10321 14903 10379 14909
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 12434 14940 12440 14952
rect 12299 14912 12440 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 8588 14872 8616 14903
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 12805 14943 12863 14949
rect 12805 14909 12817 14943
rect 12851 14940 12863 14943
rect 13078 14940 13084 14952
rect 12851 14912 13084 14940
rect 12851 14909 12863 14912
rect 12805 14903 12863 14909
rect 13078 14900 13084 14912
rect 13136 14900 13142 14952
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14940 13599 14943
rect 13722 14940 13728 14952
rect 13587 14912 13728 14940
rect 13587 14909 13599 14912
rect 13541 14903 13599 14909
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 13924 14940 13952 14980
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 15378 14968 15384 15020
rect 15436 15008 15442 15020
rect 16209 15011 16267 15017
rect 16209 15008 16221 15011
rect 15436 14980 16221 15008
rect 15436 14968 15442 14980
rect 16209 14977 16221 14980
rect 16255 14977 16267 15011
rect 16209 14971 16267 14977
rect 15470 14940 15476 14952
rect 13924 14912 15476 14940
rect 15470 14900 15476 14912
rect 15528 14900 15534 14952
rect 16224 14940 16252 14971
rect 18230 14968 18236 15020
rect 18288 15008 18294 15020
rect 19521 15011 19579 15017
rect 19521 15008 19533 15011
rect 18288 14980 19533 15008
rect 18288 14968 18294 14980
rect 19521 14977 19533 14980
rect 19567 14977 19579 15011
rect 19702 15008 19708 15020
rect 19663 14980 19708 15008
rect 19521 14971 19579 14977
rect 19702 14968 19708 14980
rect 19760 14968 19766 15020
rect 20530 14968 20536 15020
rect 20588 15008 20594 15020
rect 20732 15017 20760 15116
rect 20717 15011 20775 15017
rect 20588 14980 20633 15008
rect 20588 14968 20594 14980
rect 20717 14977 20729 15011
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 17034 14940 17040 14952
rect 16224 14912 17040 14940
rect 17034 14900 17040 14912
rect 17092 14900 17098 14952
rect 18785 14943 18843 14949
rect 18785 14909 18797 14943
rect 18831 14940 18843 14943
rect 18877 14943 18935 14949
rect 18877 14940 18889 14943
rect 18831 14912 18889 14940
rect 18831 14909 18843 14912
rect 18785 14903 18843 14909
rect 18877 14909 18889 14912
rect 18923 14940 18935 14943
rect 19429 14943 19487 14949
rect 19429 14940 19441 14943
rect 18923 14912 19441 14940
rect 18923 14909 18935 14912
rect 18877 14903 18935 14909
rect 19429 14909 19441 14912
rect 19475 14909 19487 14943
rect 19429 14903 19487 14909
rect 6328 14844 6592 14872
rect 6656 14844 8616 14872
rect 8932 14875 8990 14881
rect 6328 14832 6334 14844
rect 6178 14804 6184 14816
rect 5092 14776 6184 14804
rect 4709 14767 4767 14773
rect 6178 14764 6184 14776
rect 6236 14804 6242 14816
rect 6365 14807 6423 14813
rect 6365 14804 6377 14807
rect 6236 14776 6377 14804
rect 6236 14764 6242 14776
rect 6365 14773 6377 14776
rect 6411 14773 6423 14807
rect 6564 14804 6592 14844
rect 8932 14841 8944 14875
rect 8978 14872 8990 14875
rect 9674 14872 9680 14884
rect 8978 14844 9680 14872
rect 8978 14841 8990 14844
rect 8932 14835 8990 14841
rect 9674 14832 9680 14844
rect 9732 14832 9738 14884
rect 10229 14875 10287 14881
rect 10229 14841 10241 14875
rect 10275 14872 10287 14875
rect 10566 14875 10624 14881
rect 10566 14872 10578 14875
rect 10275 14844 10578 14872
rect 10275 14841 10287 14844
rect 10229 14835 10287 14841
rect 10566 14841 10578 14844
rect 10612 14872 10624 14875
rect 11422 14872 11428 14884
rect 10612 14844 11428 14872
rect 10612 14841 10624 14844
rect 10566 14835 10624 14841
rect 11422 14832 11428 14844
rect 11480 14832 11486 14884
rect 14360 14875 14418 14881
rect 14360 14841 14372 14875
rect 14406 14872 14418 14875
rect 14642 14872 14648 14884
rect 14406 14844 14648 14872
rect 14406 14841 14418 14844
rect 14360 14835 14418 14841
rect 14642 14832 14648 14844
rect 14700 14832 14706 14884
rect 15838 14872 15844 14884
rect 15396 14844 15844 14872
rect 7193 14807 7251 14813
rect 7193 14804 7205 14807
rect 6564 14776 7205 14804
rect 6365 14767 6423 14773
rect 7193 14773 7205 14776
rect 7239 14773 7251 14807
rect 7193 14767 7251 14773
rect 7285 14807 7343 14813
rect 7285 14773 7297 14807
rect 7331 14804 7343 14807
rect 9398 14804 9404 14816
rect 7331 14776 9404 14804
rect 7331 14773 7343 14776
rect 7285 14767 7343 14773
rect 9398 14764 9404 14776
rect 9456 14804 9462 14816
rect 10870 14804 10876 14816
rect 9456 14776 10876 14804
rect 9456 14764 9462 14776
rect 10870 14764 10876 14776
rect 10928 14764 10934 14816
rect 12069 14807 12127 14813
rect 12069 14773 12081 14807
rect 12115 14804 12127 14807
rect 12158 14804 12164 14816
rect 12115 14776 12164 14804
rect 12115 14773 12127 14776
rect 12069 14767 12127 14773
rect 12158 14764 12164 14776
rect 12216 14764 12222 14816
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 12897 14807 12955 14813
rect 12897 14804 12909 14807
rect 12860 14776 12909 14804
rect 12860 14764 12866 14776
rect 12897 14773 12909 14776
rect 12943 14773 12955 14807
rect 12897 14767 12955 14773
rect 13725 14807 13783 14813
rect 13725 14773 13737 14807
rect 13771 14804 13783 14807
rect 15396 14804 15424 14844
rect 15838 14832 15844 14844
rect 15896 14832 15902 14884
rect 16476 14875 16534 14881
rect 16476 14841 16488 14875
rect 16522 14872 16534 14875
rect 16666 14872 16672 14884
rect 16522 14844 16672 14872
rect 16522 14841 16534 14844
rect 16476 14835 16534 14841
rect 16666 14832 16672 14844
rect 16724 14832 16730 14884
rect 16942 14832 16948 14884
rect 17000 14872 17006 14884
rect 17000 14844 17724 14872
rect 17000 14832 17006 14844
rect 13771 14776 15424 14804
rect 13771 14773 13783 14776
rect 13725 14767 13783 14773
rect 15470 14764 15476 14816
rect 15528 14804 15534 14816
rect 15746 14804 15752 14816
rect 15528 14776 15573 14804
rect 15707 14776 15752 14804
rect 15528 14764 15534 14776
rect 15746 14764 15752 14776
rect 15804 14764 15810 14816
rect 17310 14764 17316 14816
rect 17368 14804 17374 14816
rect 17589 14807 17647 14813
rect 17589 14804 17601 14807
rect 17368 14776 17601 14804
rect 17368 14764 17374 14776
rect 17589 14773 17601 14776
rect 17635 14773 17647 14807
rect 17696 14804 17724 14844
rect 18414 14832 18420 14884
rect 18472 14872 18478 14884
rect 20070 14872 20076 14884
rect 18472 14844 20076 14872
rect 18472 14832 18478 14844
rect 20070 14832 20076 14844
rect 20128 14832 20134 14884
rect 18506 14804 18512 14816
rect 17696 14776 18512 14804
rect 17589 14767 17647 14773
rect 18506 14764 18512 14776
rect 18564 14764 18570 14816
rect 19058 14804 19064 14816
rect 19019 14776 19064 14804
rect 19058 14764 19064 14776
rect 19116 14764 19122 14816
rect 19334 14764 19340 14816
rect 19392 14804 19398 14816
rect 20441 14807 20499 14813
rect 20441 14804 20453 14807
rect 19392 14776 20453 14804
rect 19392 14764 19398 14776
rect 20441 14773 20453 14776
rect 20487 14773 20499 14807
rect 20441 14767 20499 14773
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 3329 14603 3387 14609
rect 3329 14569 3341 14603
rect 3375 14600 3387 14603
rect 4249 14603 4307 14609
rect 4249 14600 4261 14603
rect 3375 14572 4261 14600
rect 3375 14569 3387 14572
rect 3329 14563 3387 14569
rect 4249 14569 4261 14572
rect 4295 14569 4307 14603
rect 4249 14563 4307 14569
rect 4617 14603 4675 14609
rect 4617 14569 4629 14603
rect 4663 14600 4675 14603
rect 5534 14600 5540 14612
rect 4663 14572 5540 14600
rect 4663 14569 4675 14572
rect 4617 14563 4675 14569
rect 5534 14560 5540 14572
rect 5592 14560 5598 14612
rect 6914 14560 6920 14612
rect 6972 14600 6978 14612
rect 7561 14603 7619 14609
rect 7561 14600 7573 14603
rect 6972 14572 7573 14600
rect 6972 14560 6978 14572
rect 7561 14569 7573 14572
rect 7607 14569 7619 14603
rect 8570 14600 8576 14612
rect 8531 14572 8576 14600
rect 7561 14563 7619 14569
rect 8570 14560 8576 14572
rect 8628 14560 8634 14612
rect 8846 14560 8852 14612
rect 8904 14600 8910 14612
rect 9490 14600 9496 14612
rect 8904 14572 9496 14600
rect 8904 14560 8910 14572
rect 9490 14560 9496 14572
rect 9548 14560 9554 14612
rect 9861 14603 9919 14609
rect 9861 14569 9873 14603
rect 9907 14600 9919 14603
rect 10226 14600 10232 14612
rect 9907 14572 10232 14600
rect 9907 14569 9919 14572
rect 9861 14563 9919 14569
rect 10226 14560 10232 14572
rect 10284 14560 10290 14612
rect 10321 14603 10379 14609
rect 10321 14569 10333 14603
rect 10367 14600 10379 14603
rect 12805 14603 12863 14609
rect 12805 14600 12817 14603
rect 10367 14572 12020 14600
rect 10367 14569 10379 14572
rect 10321 14563 10379 14569
rect 3602 14492 3608 14544
rect 3660 14532 3666 14544
rect 4522 14532 4528 14544
rect 3660 14504 4528 14532
rect 3660 14492 3666 14504
rect 4522 14492 4528 14504
rect 4580 14492 4586 14544
rect 6150 14535 6208 14541
rect 6150 14532 6162 14535
rect 4632 14504 6162 14532
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 2225 14467 2283 14473
rect 2225 14464 2237 14467
rect 1443 14436 2237 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 2225 14433 2237 14436
rect 2271 14433 2283 14467
rect 2225 14427 2283 14433
rect 2866 14424 2872 14476
rect 2924 14464 2930 14476
rect 3237 14467 3295 14473
rect 3237 14464 3249 14467
rect 2924 14436 3249 14464
rect 2924 14424 2930 14436
rect 3237 14433 3249 14436
rect 3283 14433 3295 14467
rect 3237 14427 3295 14433
rect 4632 14408 4660 14504
rect 6150 14501 6162 14504
rect 6196 14501 6208 14535
rect 7282 14532 7288 14544
rect 6150 14495 6208 14501
rect 6840 14504 7288 14532
rect 4706 14424 4712 14476
rect 4764 14464 4770 14476
rect 5261 14467 5319 14473
rect 4764 14436 4809 14464
rect 4764 14424 4770 14436
rect 5261 14433 5273 14467
rect 5307 14464 5319 14467
rect 5350 14464 5356 14476
rect 5307 14436 5356 14464
rect 5307 14433 5319 14436
rect 5261 14427 5319 14433
rect 5350 14424 5356 14436
rect 5408 14424 5414 14476
rect 5905 14467 5963 14473
rect 5905 14433 5917 14467
rect 5951 14464 5963 14467
rect 6840 14464 6868 14504
rect 7282 14492 7288 14504
rect 7340 14492 7346 14544
rect 7742 14492 7748 14544
rect 7800 14532 7806 14544
rect 7800 14504 8156 14532
rect 7800 14492 7806 14504
rect 5951 14436 6868 14464
rect 5951 14433 5963 14436
rect 5905 14427 5963 14433
rect 6914 14424 6920 14476
rect 6972 14464 6978 14476
rect 7650 14464 7656 14476
rect 6972 14436 7656 14464
rect 6972 14424 6978 14436
rect 7650 14424 7656 14436
rect 7708 14424 7714 14476
rect 7926 14464 7932 14476
rect 7887 14436 7932 14464
rect 7926 14424 7932 14436
rect 7984 14424 7990 14476
rect 8128 14408 8156 14504
rect 8478 14492 8484 14544
rect 8536 14532 8542 14544
rect 8941 14535 8999 14541
rect 8941 14532 8953 14535
rect 8536 14504 8953 14532
rect 8536 14492 8542 14504
rect 8941 14501 8953 14504
rect 8987 14501 8999 14535
rect 8941 14495 8999 14501
rect 11701 14535 11759 14541
rect 11701 14501 11713 14535
rect 11747 14532 11759 14535
rect 11882 14532 11888 14544
rect 11747 14504 11888 14532
rect 11747 14501 11759 14504
rect 11701 14495 11759 14501
rect 11882 14492 11888 14504
rect 11940 14492 11946 14544
rect 11992 14532 12020 14572
rect 12544 14572 12817 14600
rect 12544 14532 12572 14572
rect 12805 14569 12817 14572
rect 12851 14569 12863 14603
rect 12805 14563 12863 14569
rect 13173 14603 13231 14609
rect 13173 14569 13185 14603
rect 13219 14600 13231 14603
rect 13725 14603 13783 14609
rect 13725 14600 13737 14603
rect 13219 14572 13737 14600
rect 13219 14569 13231 14572
rect 13173 14563 13231 14569
rect 13725 14569 13737 14572
rect 13771 14569 13783 14603
rect 13725 14563 13783 14569
rect 16025 14603 16083 14609
rect 16025 14569 16037 14603
rect 16071 14600 16083 14603
rect 16758 14600 16764 14612
rect 16071 14572 16764 14600
rect 16071 14569 16083 14572
rect 16025 14563 16083 14569
rect 16758 14560 16764 14572
rect 16816 14560 16822 14612
rect 17770 14560 17776 14612
rect 17828 14600 17834 14612
rect 18969 14603 19027 14609
rect 18969 14600 18981 14603
rect 17828 14572 18981 14600
rect 17828 14560 17834 14572
rect 18969 14569 18981 14572
rect 19015 14569 19027 14603
rect 18969 14563 19027 14569
rect 19613 14603 19671 14609
rect 19613 14569 19625 14603
rect 19659 14600 19671 14603
rect 20070 14600 20076 14612
rect 19659 14572 20076 14600
rect 19659 14569 19671 14572
rect 19613 14563 19671 14569
rect 20070 14560 20076 14572
rect 20128 14560 20134 14612
rect 20806 14560 20812 14612
rect 20864 14600 20870 14612
rect 20901 14603 20959 14609
rect 20901 14600 20913 14603
rect 20864 14572 20913 14600
rect 20864 14560 20870 14572
rect 20901 14569 20913 14572
rect 20947 14569 20959 14603
rect 20901 14563 20959 14569
rect 12710 14532 12716 14544
rect 11992 14504 12572 14532
rect 12671 14504 12716 14532
rect 12710 14492 12716 14504
rect 12768 14492 12774 14544
rect 17954 14532 17960 14544
rect 12820 14504 13952 14532
rect 9677 14467 9735 14473
rect 9677 14433 9689 14467
rect 9723 14464 9735 14467
rect 9766 14464 9772 14476
rect 9723 14436 9772 14464
rect 9723 14433 9735 14436
rect 9677 14427 9735 14433
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 10689 14467 10747 14473
rect 10689 14433 10701 14467
rect 10735 14464 10747 14467
rect 11054 14464 11060 14476
rect 10735 14436 11060 14464
rect 10735 14433 10747 14436
rect 10689 14427 10747 14433
rect 11054 14424 11060 14436
rect 11112 14424 11118 14476
rect 11606 14424 11612 14476
rect 11664 14464 11670 14476
rect 12820 14464 12848 14504
rect 13817 14467 13875 14473
rect 13817 14464 13829 14467
rect 11664 14436 12848 14464
rect 12912 14436 13829 14464
rect 11664 14424 11670 14436
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14365 2375 14399
rect 2317 14359 2375 14365
rect 2501 14399 2559 14405
rect 2501 14365 2513 14399
rect 2547 14396 2559 14399
rect 2774 14396 2780 14408
rect 2547 14368 2780 14396
rect 2547 14365 2559 14368
rect 2501 14359 2559 14365
rect 2332 14328 2360 14359
rect 2774 14356 2780 14368
rect 2832 14356 2838 14408
rect 3513 14399 3571 14405
rect 3513 14365 3525 14399
rect 3559 14396 3571 14399
rect 4614 14396 4620 14408
rect 3559 14368 4620 14396
rect 3559 14365 3571 14368
rect 3513 14359 3571 14365
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 4801 14399 4859 14405
rect 4801 14365 4813 14399
rect 4847 14365 4859 14399
rect 4801 14359 4859 14365
rect 3326 14328 3332 14340
rect 2332 14300 3332 14328
rect 3326 14288 3332 14300
rect 3384 14288 3390 14340
rect 3602 14288 3608 14340
rect 3660 14328 3666 14340
rect 4816 14328 4844 14359
rect 4982 14356 4988 14408
rect 5040 14396 5046 14408
rect 5040 14368 5488 14396
rect 5040 14356 5046 14368
rect 3660 14300 4844 14328
rect 3660 14288 3666 14300
rect 1857 14263 1915 14269
rect 1857 14229 1869 14263
rect 1903 14260 1915 14263
rect 2774 14260 2780 14272
rect 1903 14232 2780 14260
rect 1903 14229 1915 14232
rect 1857 14223 1915 14229
rect 2774 14220 2780 14232
rect 2832 14220 2838 14272
rect 2869 14263 2927 14269
rect 2869 14229 2881 14263
rect 2915 14260 2927 14263
rect 5350 14260 5356 14272
rect 2915 14232 5356 14260
rect 2915 14229 2927 14232
rect 2869 14223 2927 14229
rect 5350 14220 5356 14232
rect 5408 14220 5414 14272
rect 5460 14269 5488 14368
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 8021 14399 8079 14405
rect 8021 14396 8033 14399
rect 7432 14368 8033 14396
rect 7432 14356 7438 14368
rect 8021 14365 8033 14368
rect 8067 14365 8079 14399
rect 8021 14359 8079 14365
rect 8110 14356 8116 14408
rect 8168 14396 8174 14408
rect 8168 14368 8213 14396
rect 8168 14356 8174 14368
rect 8570 14356 8576 14408
rect 8628 14396 8634 14408
rect 8754 14396 8760 14408
rect 8628 14368 8760 14396
rect 8628 14356 8634 14368
rect 8754 14356 8760 14368
rect 8812 14356 8818 14408
rect 9033 14399 9091 14405
rect 9033 14365 9045 14399
rect 9079 14365 9091 14399
rect 9033 14359 9091 14365
rect 9048 14328 9076 14359
rect 9122 14356 9128 14408
rect 9180 14396 9186 14408
rect 9180 14368 9273 14396
rect 9180 14356 9186 14368
rect 9858 14356 9864 14408
rect 9916 14396 9922 14408
rect 10781 14399 10839 14405
rect 10781 14396 10793 14399
rect 9916 14368 10793 14396
rect 9916 14356 9922 14368
rect 10781 14365 10793 14368
rect 10827 14365 10839 14399
rect 10781 14359 10839 14365
rect 10870 14356 10876 14408
rect 10928 14396 10934 14408
rect 10928 14368 10973 14396
rect 10928 14356 10934 14368
rect 11514 14356 11520 14408
rect 11572 14396 11578 14408
rect 11793 14399 11851 14405
rect 11793 14396 11805 14399
rect 11572 14368 11805 14396
rect 11572 14356 11578 14368
rect 11793 14365 11805 14368
rect 11839 14365 11851 14399
rect 11793 14359 11851 14365
rect 11885 14399 11943 14405
rect 11885 14365 11897 14399
rect 11931 14365 11943 14399
rect 11885 14359 11943 14365
rect 6840 14300 9076 14328
rect 5445 14263 5503 14269
rect 5445 14229 5457 14263
rect 5491 14229 5503 14263
rect 5445 14223 5503 14229
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 6840 14260 6868 14300
rect 5592 14232 6868 14260
rect 7285 14263 7343 14269
rect 5592 14220 5598 14232
rect 7285 14229 7297 14263
rect 7331 14260 7343 14263
rect 7466 14260 7472 14272
rect 7331 14232 7472 14260
rect 7331 14229 7343 14232
rect 7285 14223 7343 14229
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 8294 14220 8300 14272
rect 8352 14260 8358 14272
rect 9140 14260 9168 14356
rect 10888 14328 10916 14356
rect 11900 14328 11928 14359
rect 10888 14300 11928 14328
rect 12345 14331 12403 14337
rect 12345 14297 12357 14331
rect 12391 14328 12403 14331
rect 12912 14328 12940 14436
rect 13817 14433 13829 14436
rect 13863 14433 13875 14467
rect 13817 14427 13875 14433
rect 12989 14399 13047 14405
rect 12989 14365 13001 14399
rect 13035 14396 13047 14399
rect 13078 14396 13084 14408
rect 13035 14368 13084 14396
rect 13035 14365 13047 14368
rect 12989 14359 13047 14365
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 13924 14405 13952 14504
rect 14476 14504 17960 14532
rect 14476 14473 14504 14504
rect 17954 14492 17960 14504
rect 18012 14492 18018 14544
rect 18046 14492 18052 14544
rect 18104 14532 18110 14544
rect 20165 14535 20223 14541
rect 18104 14504 19104 14532
rect 18104 14492 18110 14504
rect 14461 14467 14519 14473
rect 14461 14433 14473 14467
rect 14507 14433 14519 14467
rect 14461 14427 14519 14433
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14464 15347 14467
rect 15838 14464 15844 14476
rect 15335 14436 15844 14464
rect 15335 14433 15347 14436
rect 15289 14427 15347 14433
rect 15838 14424 15844 14436
rect 15896 14424 15902 14476
rect 16022 14424 16028 14476
rect 16080 14464 16086 14476
rect 16393 14467 16451 14473
rect 16393 14464 16405 14467
rect 16080 14436 16405 14464
rect 16080 14424 16086 14436
rect 16393 14433 16405 14436
rect 16439 14433 16451 14467
rect 17034 14464 17040 14476
rect 16995 14436 17040 14464
rect 16393 14427 16451 14433
rect 17034 14424 17040 14436
rect 17092 14424 17098 14476
rect 17310 14473 17316 14476
rect 17304 14464 17316 14473
rect 17271 14436 17316 14464
rect 17304 14427 17316 14436
rect 17310 14424 17316 14427
rect 17368 14424 17374 14476
rect 17586 14424 17592 14476
rect 17644 14464 17650 14476
rect 17644 14436 18092 14464
rect 17644 14424 17650 14436
rect 13909 14399 13967 14405
rect 13909 14365 13921 14399
rect 13955 14365 13967 14399
rect 13909 14359 13967 14365
rect 14737 14399 14795 14405
rect 14737 14365 14749 14399
rect 14783 14396 14795 14399
rect 15194 14396 15200 14408
rect 14783 14368 15200 14396
rect 14783 14365 14795 14368
rect 14737 14359 14795 14365
rect 15194 14356 15200 14368
rect 15252 14356 15258 14408
rect 15565 14399 15623 14405
rect 15565 14365 15577 14399
rect 15611 14365 15623 14399
rect 15565 14359 15623 14365
rect 13354 14328 13360 14340
rect 12391 14300 12940 14328
rect 13315 14300 13360 14328
rect 12391 14297 12403 14300
rect 12345 14291 12403 14297
rect 13354 14288 13360 14300
rect 13412 14288 13418 14340
rect 13538 14288 13544 14340
rect 13596 14328 13602 14340
rect 14918 14328 14924 14340
rect 13596 14300 14924 14328
rect 13596 14288 13602 14300
rect 14918 14288 14924 14300
rect 14976 14288 14982 14340
rect 15580 14328 15608 14359
rect 16482 14356 16488 14408
rect 16540 14396 16546 14408
rect 16666 14396 16672 14408
rect 16540 14368 16585 14396
rect 16627 14368 16672 14396
rect 16540 14356 16546 14368
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 18064 14396 18092 14436
rect 18230 14424 18236 14476
rect 18288 14464 18294 14476
rect 18877 14467 18935 14473
rect 18877 14464 18889 14467
rect 18288 14436 18889 14464
rect 18288 14424 18294 14436
rect 18877 14433 18889 14436
rect 18923 14433 18935 14467
rect 18877 14427 18935 14433
rect 19076 14405 19104 14504
rect 20165 14501 20177 14535
rect 20211 14532 20223 14535
rect 21358 14532 21364 14544
rect 20211 14504 21364 14532
rect 20211 14501 20223 14504
rect 20165 14495 20223 14501
rect 21358 14492 21364 14504
rect 21416 14492 21422 14544
rect 19061 14399 19119 14405
rect 18064 14368 18543 14396
rect 16758 14328 16764 14340
rect 15580 14300 16764 14328
rect 16758 14288 16764 14300
rect 16816 14288 16822 14340
rect 18138 14288 18144 14340
rect 18196 14328 18202 14340
rect 18417 14331 18475 14337
rect 18417 14328 18429 14331
rect 18196 14300 18429 14328
rect 18196 14288 18202 14300
rect 18417 14297 18429 14300
rect 18463 14297 18475 14331
rect 18515 14328 18543 14368
rect 19061 14365 19073 14399
rect 19107 14365 19119 14399
rect 19061 14359 19119 14365
rect 19702 14356 19708 14408
rect 19760 14396 19766 14408
rect 20349 14399 20407 14405
rect 20349 14396 20361 14399
rect 19760 14368 20361 14396
rect 19760 14356 19766 14368
rect 20349 14365 20361 14368
rect 20395 14396 20407 14399
rect 20806 14396 20812 14408
rect 20395 14368 20812 14396
rect 20395 14365 20407 14368
rect 20349 14359 20407 14365
rect 20806 14356 20812 14368
rect 20864 14356 20870 14408
rect 19334 14328 19340 14340
rect 18515 14300 19340 14328
rect 18417 14291 18475 14297
rect 19334 14288 19340 14300
rect 19392 14288 19398 14340
rect 8352 14232 9168 14260
rect 8352 14220 8358 14232
rect 11146 14220 11152 14272
rect 11204 14260 11210 14272
rect 11333 14263 11391 14269
rect 11333 14260 11345 14263
rect 11204 14232 11345 14260
rect 11204 14220 11210 14232
rect 11333 14229 11345 14232
rect 11379 14229 11391 14263
rect 11333 14223 11391 14229
rect 11606 14220 11612 14272
rect 11664 14260 11670 14272
rect 13173 14263 13231 14269
rect 13173 14260 13185 14263
rect 11664 14232 13185 14260
rect 11664 14220 11670 14232
rect 13173 14229 13185 14232
rect 13219 14229 13231 14263
rect 13173 14223 13231 14229
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 15930 14260 15936 14272
rect 13504 14232 15936 14260
rect 13504 14220 13510 14232
rect 15930 14220 15936 14232
rect 15988 14220 15994 14272
rect 16022 14220 16028 14272
rect 16080 14260 16086 14272
rect 17678 14260 17684 14272
rect 16080 14232 17684 14260
rect 16080 14220 16086 14232
rect 17678 14220 17684 14232
rect 17736 14220 17742 14272
rect 17770 14220 17776 14272
rect 17828 14260 17834 14272
rect 18509 14263 18567 14269
rect 18509 14260 18521 14263
rect 17828 14232 18521 14260
rect 17828 14220 17834 14232
rect 18509 14229 18521 14232
rect 18555 14229 18567 14263
rect 19702 14260 19708 14272
rect 19663 14232 19708 14260
rect 18509 14223 18567 14229
rect 19702 14220 19708 14232
rect 19760 14220 19766 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 1857 14059 1915 14065
rect 1857 14025 1869 14059
rect 1903 14056 1915 14059
rect 5534 14056 5540 14068
rect 1903 14028 5540 14056
rect 1903 14025 1915 14028
rect 1857 14019 1915 14025
rect 5534 14016 5540 14028
rect 5592 14016 5598 14068
rect 5721 14059 5779 14065
rect 5721 14025 5733 14059
rect 5767 14056 5779 14059
rect 5994 14056 6000 14068
rect 5767 14028 6000 14056
rect 5767 14025 5779 14028
rect 5721 14019 5779 14025
rect 5994 14016 6000 14028
rect 6052 14016 6058 14068
rect 6730 14016 6736 14068
rect 6788 14056 6794 14068
rect 9125 14059 9183 14065
rect 6788 14028 7144 14056
rect 6788 14016 6794 14028
rect 2866 13948 2872 14000
rect 2924 13988 2930 14000
rect 2924 13960 2969 13988
rect 2924 13948 2930 13960
rect 4890 13948 4896 14000
rect 4948 13988 4954 14000
rect 4948 13960 7052 13988
rect 4948 13948 4954 13960
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13920 2559 13923
rect 2590 13920 2596 13932
rect 2547 13892 2596 13920
rect 2547 13889 2559 13892
rect 2501 13883 2559 13889
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 3510 13920 3516 13932
rect 3471 13892 3516 13920
rect 3510 13880 3516 13892
rect 3568 13880 3574 13932
rect 6086 13920 6092 13932
rect 5276 13892 6092 13920
rect 5276 13864 5304 13892
rect 6086 13880 6092 13892
rect 6144 13920 6150 13932
rect 6273 13923 6331 13929
rect 6273 13920 6285 13923
rect 6144 13892 6285 13920
rect 6144 13880 6150 13892
rect 6273 13889 6285 13892
rect 6319 13889 6331 13923
rect 6730 13920 6736 13932
rect 6273 13883 6331 13889
rect 6380 13892 6736 13920
rect 2958 13812 2964 13864
rect 3016 13852 3022 13864
rect 3881 13855 3939 13861
rect 3881 13852 3893 13855
rect 3016 13824 3280 13852
rect 3016 13812 3022 13824
rect 2774 13744 2780 13796
rect 2832 13744 2838 13796
rect 3252 13784 3280 13824
rect 3528 13824 3893 13852
rect 3528 13796 3556 13824
rect 3881 13821 3893 13824
rect 3927 13821 3939 13855
rect 4137 13855 4195 13861
rect 4137 13852 4149 13855
rect 3881 13815 3939 13821
rect 3988 13824 4149 13852
rect 3329 13787 3387 13793
rect 3329 13784 3341 13787
rect 3252 13756 3341 13784
rect 3329 13753 3341 13756
rect 3375 13753 3387 13787
rect 3329 13747 3387 13753
rect 3510 13744 3516 13796
rect 3568 13744 3574 13796
rect 3694 13744 3700 13796
rect 3752 13784 3758 13796
rect 3988 13784 4016 13824
rect 4137 13821 4149 13824
rect 4183 13821 4195 13855
rect 4982 13852 4988 13864
rect 4137 13815 4195 13821
rect 4264 13824 4988 13852
rect 3752 13756 4016 13784
rect 3752 13744 3758 13756
rect 1394 13716 1400 13728
rect 1355 13688 1400 13716
rect 1394 13676 1400 13688
rect 1452 13676 1458 13728
rect 1854 13676 1860 13728
rect 1912 13716 1918 13728
rect 2225 13719 2283 13725
rect 2225 13716 2237 13719
rect 1912 13688 2237 13716
rect 1912 13676 1918 13688
rect 2225 13685 2237 13688
rect 2271 13685 2283 13719
rect 2225 13679 2283 13685
rect 2317 13719 2375 13725
rect 2317 13685 2329 13719
rect 2363 13716 2375 13719
rect 2590 13716 2596 13728
rect 2363 13688 2596 13716
rect 2363 13685 2375 13688
rect 2317 13679 2375 13685
rect 2590 13676 2596 13688
rect 2648 13676 2654 13728
rect 2792 13716 2820 13744
rect 3237 13719 3295 13725
rect 3237 13716 3249 13719
rect 2792 13688 3249 13716
rect 3237 13685 3249 13688
rect 3283 13685 3295 13719
rect 3237 13679 3295 13685
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 4264 13716 4292 13824
rect 4982 13812 4988 13824
rect 5040 13812 5046 13864
rect 5258 13812 5264 13864
rect 5316 13812 5322 13864
rect 5350 13812 5356 13864
rect 5408 13852 5414 13864
rect 6181 13855 6239 13861
rect 5408 13824 6132 13852
rect 5408 13812 5414 13824
rect 5276 13725 5304 13812
rect 6104 13784 6132 13824
rect 6181 13821 6193 13855
rect 6227 13852 6239 13855
rect 6380 13852 6408 13892
rect 6730 13880 6736 13892
rect 6788 13880 6794 13932
rect 7024 13929 7052 13960
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13889 7067 13923
rect 7116 13920 7144 14028
rect 9125 14025 9137 14059
rect 9171 14056 9183 14059
rect 9674 14056 9680 14068
rect 9171 14028 9680 14056
rect 9171 14025 9183 14028
rect 9125 14019 9183 14025
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 9953 14059 10011 14065
rect 9953 14025 9965 14059
rect 9999 14056 10011 14059
rect 12710 14056 12716 14068
rect 9999 14028 12716 14056
rect 9999 14025 10011 14028
rect 9953 14019 10011 14025
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 12802 14016 12808 14068
rect 12860 14056 12866 14068
rect 13170 14056 13176 14068
rect 12860 14028 13176 14056
rect 12860 14016 12866 14028
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 14366 14056 14372 14068
rect 13780 14028 14372 14056
rect 13780 14016 13786 14028
rect 14366 14016 14372 14028
rect 14424 14016 14430 14068
rect 14737 14059 14795 14065
rect 14737 14025 14749 14059
rect 14783 14056 14795 14059
rect 16298 14056 16304 14068
rect 14783 14028 16304 14056
rect 14783 14025 14795 14028
rect 14737 14019 14795 14025
rect 16298 14016 16304 14028
rect 16356 14016 16362 14068
rect 16761 14059 16819 14065
rect 16761 14025 16773 14059
rect 16807 14056 16819 14059
rect 16850 14056 16856 14068
rect 16807 14028 16856 14056
rect 16807 14025 16819 14028
rect 16761 14019 16819 14025
rect 16850 14016 16856 14028
rect 16908 14016 16914 14068
rect 17034 14016 17040 14068
rect 17092 14016 17098 14068
rect 17494 14016 17500 14068
rect 17552 14056 17558 14068
rect 20898 14056 20904 14068
rect 17552 14028 19104 14056
rect 20859 14028 20904 14056
rect 17552 14016 17558 14028
rect 9585 13991 9643 13997
rect 9585 13957 9597 13991
rect 9631 13988 9643 13991
rect 12526 13988 12532 14000
rect 9631 13960 12532 13988
rect 9631 13957 9643 13960
rect 9585 13951 9643 13957
rect 12526 13948 12532 13960
rect 12584 13948 12590 14000
rect 14185 13991 14243 13997
rect 14185 13957 14197 13991
rect 14231 13957 14243 13991
rect 14185 13951 14243 13957
rect 16485 13991 16543 13997
rect 16485 13957 16497 13991
rect 16531 13957 16543 13991
rect 17052 13988 17080 14016
rect 17052 13960 17540 13988
rect 16485 13951 16543 13957
rect 7116 13892 7880 13920
rect 7009 13883 7067 13889
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6227 13824 6408 13852
rect 6472 13824 6837 13852
rect 6227 13821 6239 13824
rect 6181 13815 6239 13821
rect 6472 13784 6500 13824
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 7282 13812 7288 13864
rect 7340 13852 7346 13864
rect 7745 13855 7803 13861
rect 7745 13852 7757 13855
rect 7340 13824 7757 13852
rect 7340 13812 7346 13824
rect 7745 13821 7757 13824
rect 7791 13821 7803 13855
rect 7852 13852 7880 13892
rect 8772 13892 9628 13920
rect 8012 13855 8070 13861
rect 8012 13852 8024 13855
rect 7852 13824 8024 13852
rect 7745 13815 7803 13821
rect 8012 13821 8024 13824
rect 8058 13852 8070 13855
rect 8772 13852 8800 13892
rect 8058 13824 8800 13852
rect 8058 13821 8070 13824
rect 8012 13815 8070 13821
rect 8846 13812 8852 13864
rect 8904 13852 8910 13864
rect 9401 13855 9459 13861
rect 8904 13824 9260 13852
rect 8904 13812 8910 13824
rect 6104 13756 6500 13784
rect 6546 13744 6552 13796
rect 6604 13784 6610 13796
rect 9232 13784 9260 13824
rect 9401 13821 9413 13855
rect 9447 13852 9459 13855
rect 9490 13852 9496 13864
rect 9447 13824 9496 13852
rect 9447 13821 9459 13824
rect 9401 13815 9459 13821
rect 9490 13812 9496 13824
rect 9548 13812 9554 13864
rect 9600 13852 9628 13892
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 10226 13920 10232 13932
rect 9732 13892 10232 13920
rect 9732 13880 9738 13892
rect 10226 13880 10232 13892
rect 10284 13920 10290 13932
rect 10505 13923 10563 13929
rect 10505 13920 10517 13923
rect 10284 13892 10517 13920
rect 10284 13880 10290 13892
rect 10505 13889 10517 13892
rect 10551 13920 10563 13923
rect 10870 13920 10876 13932
rect 10551 13892 10876 13920
rect 10551 13889 10563 13892
rect 10505 13883 10563 13889
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 11517 13923 11575 13929
rect 11517 13889 11529 13923
rect 11563 13889 11575 13923
rect 14200 13920 14228 13951
rect 14274 13920 14280 13932
rect 14187 13892 14280 13920
rect 11517 13883 11575 13889
rect 11532 13852 11560 13883
rect 14274 13880 14280 13892
rect 14332 13920 14338 13932
rect 16500 13920 16528 13951
rect 16666 13920 16672 13932
rect 14332 13892 15240 13920
rect 16500 13892 16672 13920
rect 14332 13880 14338 13892
rect 12066 13852 12072 13864
rect 9600 13824 12072 13852
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 12805 13855 12863 13861
rect 12805 13821 12817 13855
rect 12851 13821 12863 13855
rect 12805 13815 12863 13821
rect 13072 13855 13130 13861
rect 13072 13821 13084 13855
rect 13118 13852 13130 13855
rect 14182 13852 14188 13864
rect 13118 13824 14188 13852
rect 13118 13821 13130 13824
rect 13072 13815 13130 13821
rect 11333 13787 11391 13793
rect 11333 13784 11345 13787
rect 6604 13756 8975 13784
rect 9232 13756 11345 13784
rect 6604 13744 6610 13756
rect 4028 13688 4292 13716
rect 5261 13719 5319 13725
rect 4028 13676 4034 13688
rect 5261 13685 5273 13719
rect 5307 13685 5319 13719
rect 5261 13679 5319 13685
rect 5994 13676 6000 13728
rect 6052 13716 6058 13728
rect 6089 13719 6147 13725
rect 6089 13716 6101 13719
rect 6052 13688 6101 13716
rect 6052 13676 6058 13688
rect 6089 13685 6101 13688
rect 6135 13685 6147 13719
rect 6089 13679 6147 13685
rect 6270 13676 6276 13728
rect 6328 13716 6334 13728
rect 8846 13716 8852 13728
rect 6328 13688 8852 13716
rect 6328 13676 6334 13688
rect 8846 13676 8852 13688
rect 8904 13676 8910 13728
rect 8947 13716 8975 13756
rect 11333 13753 11345 13756
rect 11379 13784 11391 13787
rect 12250 13784 12256 13796
rect 11379 13756 12256 13784
rect 11379 13753 11391 13756
rect 11333 13747 11391 13753
rect 12250 13744 12256 13756
rect 12308 13744 12314 13796
rect 12820 13784 12848 13815
rect 14182 13812 14188 13824
rect 14240 13812 14246 13864
rect 14553 13855 14611 13861
rect 14553 13821 14565 13855
rect 14599 13852 14611 13855
rect 14642 13852 14648 13864
rect 14599 13824 14648 13852
rect 14599 13821 14611 13824
rect 14553 13815 14611 13821
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 15010 13812 15016 13864
rect 15068 13852 15074 13864
rect 15105 13855 15163 13861
rect 15105 13852 15117 13855
rect 15068 13824 15117 13852
rect 15068 13812 15074 13824
rect 15105 13821 15117 13824
rect 15151 13821 15163 13855
rect 15212 13852 15240 13892
rect 16666 13880 16672 13892
rect 16724 13920 16730 13932
rect 17405 13923 17463 13929
rect 17405 13920 17417 13923
rect 16724 13892 17417 13920
rect 16724 13880 16730 13892
rect 17405 13889 17417 13892
rect 17451 13889 17463 13923
rect 17405 13883 17463 13889
rect 15212 13824 17347 13852
rect 15105 13815 15163 13821
rect 13538 13784 13544 13796
rect 12820 13756 13544 13784
rect 13538 13744 13544 13756
rect 13596 13784 13602 13796
rect 15028 13784 15056 13812
rect 13596 13756 15056 13784
rect 13596 13744 13602 13756
rect 15194 13744 15200 13796
rect 15252 13784 15258 13796
rect 15350 13787 15408 13793
rect 15350 13784 15362 13787
rect 15252 13756 15362 13784
rect 15252 13744 15258 13756
rect 15350 13753 15362 13756
rect 15396 13753 15408 13787
rect 15350 13747 15408 13753
rect 16850 13744 16856 13796
rect 16908 13784 16914 13796
rect 17221 13787 17279 13793
rect 17221 13784 17233 13787
rect 16908 13756 17233 13784
rect 16908 13744 16914 13756
rect 17221 13753 17233 13756
rect 17267 13753 17279 13787
rect 17221 13747 17279 13753
rect 10318 13716 10324 13728
rect 8947 13688 10324 13716
rect 10318 13676 10324 13688
rect 10376 13676 10382 13728
rect 10413 13719 10471 13725
rect 10413 13685 10425 13719
rect 10459 13716 10471 13719
rect 10965 13719 11023 13725
rect 10965 13716 10977 13719
rect 10459 13688 10977 13716
rect 10459 13685 10471 13688
rect 10413 13679 10471 13685
rect 10965 13685 10977 13688
rect 11011 13685 11023 13719
rect 11422 13716 11428 13728
rect 11383 13688 11428 13716
rect 10965 13679 11023 13685
rect 11422 13676 11428 13688
rect 11480 13676 11486 13728
rect 11698 13676 11704 13728
rect 11756 13716 11762 13728
rect 15470 13716 15476 13728
rect 11756 13688 15476 13716
rect 11756 13676 11762 13688
rect 15470 13676 15476 13688
rect 15528 13676 15534 13728
rect 17126 13716 17132 13728
rect 17087 13688 17132 13716
rect 17126 13676 17132 13688
rect 17184 13676 17190 13728
rect 17319 13716 17347 13824
rect 17420 13784 17448 13883
rect 17512 13852 17540 13960
rect 17954 13880 17960 13932
rect 18012 13920 18018 13932
rect 18012 13892 18184 13920
rect 18012 13880 18018 13892
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 17512 13824 18061 13852
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18156 13852 18184 13892
rect 18305 13855 18363 13861
rect 18305 13852 18317 13855
rect 18156 13824 18317 13852
rect 18049 13815 18107 13821
rect 18305 13821 18317 13824
rect 18351 13821 18363 13855
rect 19076 13852 19104 14028
rect 20898 14016 20904 14028
rect 20956 14016 20962 14068
rect 19426 13948 19432 14000
rect 19484 13988 19490 14000
rect 19705 13991 19763 13997
rect 19705 13988 19717 13991
rect 19484 13960 19717 13988
rect 19484 13948 19490 13960
rect 19705 13957 19717 13960
rect 19751 13957 19763 13991
rect 19705 13951 19763 13957
rect 19334 13880 19340 13932
rect 19392 13920 19398 13932
rect 20257 13923 20315 13929
rect 20257 13920 20269 13923
rect 19392 13892 20269 13920
rect 19392 13880 19398 13892
rect 20257 13889 20269 13892
rect 20303 13889 20315 13923
rect 20257 13883 20315 13889
rect 20162 13852 20168 13864
rect 19076 13824 19472 13852
rect 20123 13824 20168 13852
rect 18305 13815 18363 13821
rect 17862 13784 17868 13796
rect 17420 13756 17868 13784
rect 17862 13744 17868 13756
rect 17920 13744 17926 13796
rect 17586 13716 17592 13728
rect 17319 13688 17592 13716
rect 17586 13676 17592 13688
rect 17644 13676 17650 13728
rect 17954 13676 17960 13728
rect 18012 13716 18018 13728
rect 19242 13716 19248 13728
rect 18012 13688 19248 13716
rect 18012 13676 18018 13688
rect 19242 13676 19248 13688
rect 19300 13676 19306 13728
rect 19444 13725 19472 13824
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 20714 13852 20720 13864
rect 20675 13824 20720 13852
rect 20714 13812 20720 13824
rect 20772 13812 20778 13864
rect 19429 13719 19487 13725
rect 19429 13685 19441 13719
rect 19475 13685 19487 13719
rect 20070 13716 20076 13728
rect 20031 13688 20076 13716
rect 19429 13679 19487 13685
rect 20070 13676 20076 13688
rect 20128 13676 20134 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 2406 13472 2412 13524
rect 2464 13512 2470 13524
rect 3510 13512 3516 13524
rect 2464 13484 3516 13512
rect 2464 13472 2470 13484
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 4525 13515 4583 13521
rect 4525 13481 4537 13515
rect 4571 13512 4583 13515
rect 5169 13515 5227 13521
rect 5169 13512 5181 13515
rect 4571 13484 5181 13512
rect 4571 13481 4583 13484
rect 4525 13475 4583 13481
rect 5169 13481 5181 13484
rect 5215 13481 5227 13515
rect 5169 13475 5227 13481
rect 5442 13472 5448 13524
rect 5500 13512 5506 13524
rect 6825 13515 6883 13521
rect 6825 13512 6837 13515
rect 5500 13484 6837 13512
rect 5500 13472 5506 13484
rect 6825 13481 6837 13484
rect 6871 13481 6883 13515
rect 6825 13475 6883 13481
rect 7374 13472 7380 13524
rect 7432 13512 7438 13524
rect 7432 13484 11008 13512
rect 7432 13472 7438 13484
rect 1857 13447 1915 13453
rect 1857 13413 1869 13447
rect 1903 13444 1915 13447
rect 5074 13444 5080 13456
rect 1903 13416 5080 13444
rect 1903 13413 1915 13416
rect 1857 13407 1915 13413
rect 5074 13404 5080 13416
rect 5132 13404 5138 13456
rect 5537 13447 5595 13453
rect 5537 13413 5549 13447
rect 5583 13444 5595 13447
rect 6270 13444 6276 13456
rect 5583 13416 6276 13444
rect 5583 13413 5595 13416
rect 5537 13407 5595 13413
rect 6270 13404 6276 13416
rect 6328 13404 6334 13456
rect 7282 13404 7288 13456
rect 7340 13444 7346 13456
rect 7834 13444 7840 13456
rect 7340 13416 7840 13444
rect 7340 13404 7346 13416
rect 7834 13404 7840 13416
rect 7892 13404 7898 13456
rect 8297 13447 8355 13453
rect 8297 13413 8309 13447
rect 8343 13444 8355 13447
rect 9858 13444 9864 13456
rect 8343 13416 9864 13444
rect 8343 13413 8355 13416
rect 8297 13407 8355 13413
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 10137 13447 10195 13453
rect 10137 13413 10149 13447
rect 10183 13444 10195 13447
rect 10870 13444 10876 13456
rect 10183 13416 10876 13444
rect 10183 13413 10195 13416
rect 10137 13407 10195 13413
rect 10870 13404 10876 13416
rect 10928 13404 10934 13456
rect 10980 13444 11008 13484
rect 11054 13472 11060 13524
rect 11112 13512 11118 13524
rect 11241 13515 11299 13521
rect 11241 13512 11253 13515
rect 11112 13484 11253 13512
rect 11112 13472 11118 13484
rect 11241 13481 11253 13484
rect 11287 13481 11299 13515
rect 11241 13475 11299 13481
rect 11514 13472 11520 13524
rect 11572 13512 11578 13524
rect 11609 13515 11667 13521
rect 11609 13512 11621 13515
rect 11572 13484 11621 13512
rect 11572 13472 11578 13484
rect 11609 13481 11621 13484
rect 11655 13481 11667 13515
rect 11609 13475 11667 13481
rect 12066 13472 12072 13524
rect 12124 13512 12130 13524
rect 12529 13515 12587 13521
rect 12124 13484 12204 13512
rect 12124 13472 12130 13484
rect 11698 13444 11704 13456
rect 10980 13416 11704 13444
rect 11698 13404 11704 13416
rect 11756 13404 11762 13456
rect 1578 13376 1584 13388
rect 1539 13348 1584 13376
rect 1578 13336 1584 13348
rect 1636 13336 1642 13388
rect 2317 13379 2375 13385
rect 2317 13345 2329 13379
rect 2363 13376 2375 13379
rect 2406 13376 2412 13388
rect 2363 13348 2412 13376
rect 2363 13345 2375 13348
rect 2317 13339 2375 13345
rect 2406 13336 2412 13348
rect 2464 13336 2470 13388
rect 2590 13385 2596 13388
rect 2584 13376 2596 13385
rect 2503 13348 2596 13376
rect 2584 13339 2596 13348
rect 2648 13376 2654 13388
rect 4617 13379 4675 13385
rect 2648 13348 4108 13376
rect 2590 13336 2596 13339
rect 2648 13336 2654 13348
rect 4080 13320 4108 13348
rect 4617 13345 4629 13379
rect 4663 13376 4675 13379
rect 5442 13376 5448 13388
rect 4663 13348 5448 13376
rect 4663 13345 4675 13348
rect 4617 13339 4675 13345
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13345 6239 13379
rect 6181 13339 6239 13345
rect 7193 13379 7251 13385
rect 7193 13345 7205 13379
rect 7239 13376 7251 13379
rect 7742 13376 7748 13388
rect 7239 13348 7748 13376
rect 7239 13345 7251 13348
rect 7193 13339 7251 13345
rect 4062 13268 4068 13320
rect 4120 13308 4126 13320
rect 4709 13311 4767 13317
rect 4709 13308 4721 13311
rect 4120 13280 4721 13308
rect 4120 13268 4126 13280
rect 4709 13277 4721 13280
rect 4755 13277 4767 13311
rect 5626 13308 5632 13320
rect 5587 13280 5632 13308
rect 4709 13271 4767 13277
rect 5626 13268 5632 13280
rect 5684 13268 5690 13320
rect 5718 13268 5724 13320
rect 5776 13308 5782 13320
rect 5776 13280 5821 13308
rect 5776 13268 5782 13280
rect 6086 13240 6092 13252
rect 3528 13212 6092 13240
rect 1946 13132 1952 13184
rect 2004 13172 2010 13184
rect 3528 13172 3556 13212
rect 6086 13200 6092 13212
rect 6144 13200 6150 13252
rect 6196 13240 6224 13339
rect 7742 13336 7748 13348
rect 7800 13336 7806 13388
rect 8205 13379 8263 13385
rect 8205 13345 8217 13379
rect 8251 13376 8263 13379
rect 8754 13376 8760 13388
rect 8251 13348 8760 13376
rect 8251 13345 8263 13348
rect 8205 13339 8263 13345
rect 8754 13336 8760 13348
rect 8812 13336 8818 13388
rect 8849 13379 8907 13385
rect 8849 13345 8861 13379
rect 8895 13345 8907 13379
rect 8849 13339 8907 13345
rect 7282 13308 7288 13320
rect 7243 13280 7288 13308
rect 7282 13268 7288 13280
rect 7340 13268 7346 13320
rect 7469 13311 7527 13317
rect 7469 13277 7481 13311
rect 7515 13308 7527 13311
rect 8294 13308 8300 13320
rect 7515 13280 8300 13308
rect 7515 13277 7527 13280
rect 7469 13271 7527 13277
rect 8294 13268 8300 13280
rect 8352 13268 8358 13320
rect 8478 13308 8484 13320
rect 8439 13280 8484 13308
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 8864 13308 8892 13339
rect 9306 13336 9312 13388
rect 9364 13376 9370 13388
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 9364 13348 10057 13376
rect 9364 13336 9370 13348
rect 10045 13345 10057 13348
rect 10091 13345 10103 13379
rect 10689 13379 10747 13385
rect 10689 13376 10701 13379
rect 10045 13339 10103 13345
rect 10612 13348 10701 13376
rect 10612 13320 10640 13348
rect 10689 13345 10701 13348
rect 10735 13345 10747 13379
rect 10689 13339 10747 13345
rect 11422 13336 11428 13388
rect 11480 13376 11486 13388
rect 11790 13376 11796 13388
rect 11480 13348 11796 13376
rect 11480 13336 11486 13348
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 9490 13308 9496 13320
rect 8864 13280 9496 13308
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 10284 13280 10329 13308
rect 10284 13268 10290 13280
rect 10594 13268 10600 13320
rect 10652 13268 10658 13320
rect 11698 13308 11704 13320
rect 11659 13280 11704 13308
rect 11698 13268 11704 13280
rect 11756 13268 11762 13320
rect 11885 13311 11943 13317
rect 11885 13277 11897 13311
rect 11931 13308 11943 13311
rect 12176 13308 12204 13484
rect 12529 13481 12541 13515
rect 12575 13512 12587 13515
rect 15289 13515 15347 13521
rect 12575 13484 14228 13512
rect 12575 13481 12587 13484
rect 12529 13475 12587 13481
rect 12897 13447 12955 13453
rect 12897 13413 12909 13447
rect 12943 13444 12955 13447
rect 14090 13444 14096 13456
rect 12943 13416 14096 13444
rect 12943 13413 12955 13416
rect 12897 13407 12955 13413
rect 14090 13404 14096 13416
rect 14148 13404 14154 13456
rect 14200 13444 14228 13484
rect 15289 13481 15301 13515
rect 15335 13481 15347 13515
rect 15289 13475 15347 13481
rect 14550 13444 14556 13456
rect 14200 13416 14556 13444
rect 14550 13404 14556 13416
rect 14608 13404 14614 13456
rect 15304 13444 15332 13475
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 15749 13515 15807 13521
rect 15749 13512 15761 13515
rect 15528 13484 15761 13512
rect 15528 13472 15534 13484
rect 15749 13481 15761 13484
rect 15795 13481 15807 13515
rect 15749 13475 15807 13481
rect 16393 13515 16451 13521
rect 16393 13481 16405 13515
rect 16439 13512 16451 13515
rect 17126 13512 17132 13524
rect 16439 13484 17132 13512
rect 16439 13481 16451 13484
rect 16393 13475 16451 13481
rect 17126 13472 17132 13484
rect 17184 13472 17190 13524
rect 17402 13472 17408 13524
rect 17460 13512 17466 13524
rect 17773 13515 17831 13521
rect 17773 13512 17785 13515
rect 17460 13484 17785 13512
rect 17460 13472 17466 13484
rect 17773 13481 17785 13484
rect 17819 13481 17831 13515
rect 17773 13475 17831 13481
rect 17862 13472 17868 13524
rect 17920 13512 17926 13524
rect 19429 13515 19487 13521
rect 19429 13512 19441 13515
rect 17920 13484 19441 13512
rect 17920 13472 17926 13484
rect 19429 13481 19441 13484
rect 19475 13481 19487 13515
rect 19429 13475 19487 13481
rect 19702 13472 19708 13524
rect 19760 13512 19766 13524
rect 19797 13515 19855 13521
rect 19797 13512 19809 13515
rect 19760 13484 19809 13512
rect 19760 13472 19766 13484
rect 19797 13481 19809 13484
rect 19843 13481 19855 13515
rect 19797 13475 19855 13481
rect 16850 13444 16856 13456
rect 15304 13416 16856 13444
rect 16850 13404 16856 13416
rect 16908 13404 16914 13456
rect 17313 13447 17371 13453
rect 17313 13413 17325 13447
rect 17359 13444 17371 13447
rect 18690 13444 18696 13456
rect 17359 13416 18696 13444
rect 17359 13413 17371 13416
rect 17313 13407 17371 13413
rect 18690 13404 18696 13416
rect 18748 13404 18754 13456
rect 19058 13404 19064 13456
rect 19116 13444 19122 13456
rect 19889 13447 19947 13453
rect 19889 13444 19901 13447
rect 19116 13416 19901 13444
rect 19116 13404 19122 13416
rect 19889 13413 19901 13416
rect 19935 13413 19947 13447
rect 19889 13407 19947 13413
rect 13630 13376 13636 13388
rect 13188 13348 13636 13376
rect 12986 13308 12992 13320
rect 11931 13280 12204 13308
rect 12947 13280 12992 13308
rect 11931 13277 11943 13280
rect 11885 13271 11943 13277
rect 12986 13268 12992 13280
rect 13044 13268 13050 13320
rect 13188 13317 13216 13348
rect 13630 13336 13636 13348
rect 13688 13336 13694 13388
rect 13808 13379 13866 13385
rect 13808 13345 13820 13379
rect 13854 13376 13866 13379
rect 14274 13376 14280 13388
rect 13854 13348 14280 13376
rect 13854 13345 13866 13348
rect 13808 13339 13866 13345
rect 14274 13336 14280 13348
rect 14332 13336 14338 13388
rect 14642 13336 14648 13388
rect 14700 13376 14706 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 14700 13348 15669 13376
rect 14700 13336 14706 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 16574 13336 16580 13388
rect 16632 13376 16638 13388
rect 16761 13379 16819 13385
rect 16761 13376 16773 13379
rect 16632 13348 16773 13376
rect 16632 13336 16638 13348
rect 16761 13345 16773 13348
rect 16807 13345 16819 13379
rect 16761 13339 16819 13345
rect 17770 13336 17776 13388
rect 17828 13376 17834 13388
rect 17865 13379 17923 13385
rect 17865 13376 17877 13379
rect 17828 13348 17877 13376
rect 17828 13336 17834 13348
rect 17865 13345 17877 13348
rect 17911 13345 17923 13379
rect 17865 13339 17923 13345
rect 18046 13336 18052 13388
rect 18104 13376 18110 13388
rect 18785 13379 18843 13385
rect 18785 13376 18797 13379
rect 18104 13348 18797 13376
rect 18104 13336 18110 13348
rect 18785 13345 18797 13348
rect 18831 13376 18843 13379
rect 20346 13376 20352 13388
rect 18831 13348 20352 13376
rect 18831 13345 18843 13348
rect 18785 13339 18843 13345
rect 20346 13336 20352 13348
rect 20404 13336 20410 13388
rect 13173 13311 13231 13317
rect 13173 13277 13185 13311
rect 13219 13277 13231 13311
rect 13538 13308 13544 13320
rect 13499 13280 13544 13308
rect 13173 13271 13231 13277
rect 13538 13268 13544 13280
rect 13596 13268 13602 13320
rect 15013 13311 15071 13317
rect 15013 13277 15025 13311
rect 15059 13308 15071 13311
rect 15194 13308 15200 13320
rect 15059 13280 15200 13308
rect 15059 13277 15071 13280
rect 15013 13271 15071 13277
rect 15194 13268 15200 13280
rect 15252 13308 15258 13320
rect 15930 13308 15936 13320
rect 15252 13280 15936 13308
rect 15252 13268 15258 13280
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 16850 13308 16856 13320
rect 16811 13280 16856 13308
rect 16850 13268 16856 13280
rect 16908 13268 16914 13320
rect 16942 13268 16948 13320
rect 17000 13308 17006 13320
rect 17000 13280 17045 13308
rect 17000 13268 17006 13280
rect 17310 13268 17316 13320
rect 17368 13308 17374 13320
rect 17957 13311 18015 13317
rect 17957 13308 17969 13311
rect 17368 13280 17969 13308
rect 17368 13268 17374 13280
rect 17957 13277 17969 13280
rect 18003 13277 18015 13311
rect 17957 13271 18015 13277
rect 18230 13268 18236 13320
rect 18288 13308 18294 13320
rect 18877 13311 18935 13317
rect 18877 13308 18889 13311
rect 18288 13280 18889 13308
rect 18288 13268 18294 13280
rect 18877 13277 18889 13280
rect 18923 13277 18935 13311
rect 19058 13308 19064 13320
rect 19019 13280 19064 13308
rect 18877 13271 18935 13277
rect 19058 13268 19064 13280
rect 19116 13268 19122 13320
rect 19334 13268 19340 13320
rect 19392 13268 19398 13320
rect 19702 13268 19708 13320
rect 19760 13308 19766 13320
rect 19886 13308 19892 13320
rect 19760 13280 19892 13308
rect 19760 13268 19766 13280
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 19981 13311 20039 13317
rect 19981 13277 19993 13311
rect 20027 13277 20039 13311
rect 19981 13271 20039 13277
rect 10318 13240 10324 13252
rect 6196 13212 10324 13240
rect 10318 13200 10324 13212
rect 10376 13200 10382 13252
rect 10873 13243 10931 13249
rect 10873 13209 10885 13243
rect 10919 13240 10931 13243
rect 18782 13240 18788 13252
rect 10919 13212 13584 13240
rect 10919 13209 10931 13212
rect 10873 13203 10931 13209
rect 3694 13172 3700 13184
rect 2004 13144 3556 13172
rect 3655 13144 3700 13172
rect 2004 13132 2010 13144
rect 3694 13132 3700 13144
rect 3752 13132 3758 13184
rect 4154 13172 4160 13184
rect 4115 13144 4160 13172
rect 4154 13132 4160 13144
rect 4212 13132 4218 13184
rect 4982 13132 4988 13184
rect 5040 13172 5046 13184
rect 6365 13175 6423 13181
rect 6365 13172 6377 13175
rect 5040 13144 6377 13172
rect 5040 13132 5046 13144
rect 6365 13141 6377 13144
rect 6411 13141 6423 13175
rect 6365 13135 6423 13141
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 7837 13175 7895 13181
rect 7837 13172 7849 13175
rect 7708 13144 7849 13172
rect 7708 13132 7714 13144
rect 7837 13141 7849 13144
rect 7883 13141 7895 13175
rect 7837 13135 7895 13141
rect 9033 13175 9091 13181
rect 9033 13141 9045 13175
rect 9079 13172 9091 13175
rect 9398 13172 9404 13184
rect 9079 13144 9404 13172
rect 9079 13141 9091 13144
rect 9033 13135 9091 13141
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 9677 13175 9735 13181
rect 9677 13141 9689 13175
rect 9723 13172 9735 13175
rect 11054 13172 11060 13184
rect 9723 13144 11060 13172
rect 9723 13141 9735 13144
rect 9677 13135 9735 13141
rect 11054 13132 11060 13144
rect 11112 13132 11118 13184
rect 13556 13172 13584 13212
rect 14844 13212 18788 13240
rect 14844 13172 14872 13212
rect 18782 13200 18788 13212
rect 18840 13200 18846 13252
rect 19352 13240 19380 13268
rect 19996 13240 20024 13271
rect 19352 13212 20024 13240
rect 19904 13184 19932 13212
rect 13556 13144 14872 13172
rect 14921 13175 14979 13181
rect 14921 13141 14933 13175
rect 14967 13172 14979 13175
rect 15013 13175 15071 13181
rect 15013 13172 15025 13175
rect 14967 13144 15025 13172
rect 14967 13141 14979 13144
rect 14921 13135 14979 13141
rect 15013 13141 15025 13144
rect 15059 13141 15071 13175
rect 15013 13135 15071 13141
rect 15378 13132 15384 13184
rect 15436 13172 15442 13184
rect 15562 13172 15568 13184
rect 15436 13144 15568 13172
rect 15436 13132 15442 13144
rect 15562 13132 15568 13144
rect 15620 13132 15626 13184
rect 17313 13175 17371 13181
rect 17313 13141 17325 13175
rect 17359 13172 17371 13175
rect 17405 13175 17463 13181
rect 17405 13172 17417 13175
rect 17359 13144 17417 13172
rect 17359 13141 17371 13144
rect 17313 13135 17371 13141
rect 17405 13141 17417 13144
rect 17451 13141 17463 13175
rect 17405 13135 17463 13141
rect 18417 13175 18475 13181
rect 18417 13141 18429 13175
rect 18463 13172 18475 13175
rect 19334 13172 19340 13184
rect 18463 13144 19340 13172
rect 18463 13141 18475 13144
rect 18417 13135 18475 13141
rect 19334 13132 19340 13144
rect 19392 13132 19398 13184
rect 19886 13132 19892 13184
rect 19944 13132 19950 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 4154 12968 4160 12980
rect 2056 12940 4160 12968
rect 2056 12841 2084 12940
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 5442 12968 5448 12980
rect 5403 12940 5448 12968
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 6454 12968 6460 12980
rect 6415 12940 6460 12968
rect 6454 12928 6460 12940
rect 6512 12928 6518 12980
rect 6822 12928 6828 12980
rect 6880 12968 6886 12980
rect 7190 12968 7196 12980
rect 6880 12940 7196 12968
rect 6880 12928 6886 12940
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 7466 12928 7472 12980
rect 7524 12968 7530 12980
rect 7524 12940 8432 12968
rect 7524 12928 7530 12940
rect 3973 12903 4031 12909
rect 3973 12869 3985 12903
rect 4019 12900 4031 12903
rect 4062 12900 4068 12912
rect 4019 12872 4068 12900
rect 4019 12869 4031 12872
rect 3973 12863 4031 12869
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 6086 12860 6092 12912
rect 6144 12900 6150 12912
rect 6144 12872 6776 12900
rect 6144 12860 6150 12872
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12801 2099 12835
rect 2041 12795 2099 12801
rect 2225 12835 2283 12841
rect 2225 12801 2237 12835
rect 2271 12832 2283 12835
rect 4801 12835 4859 12841
rect 4801 12832 4813 12835
rect 2271 12804 2728 12832
rect 2271 12801 2283 12804
rect 2225 12795 2283 12801
rect 2406 12724 2412 12776
rect 2464 12764 2470 12776
rect 2593 12767 2651 12773
rect 2593 12764 2605 12767
rect 2464 12736 2605 12764
rect 2464 12724 2470 12736
rect 2593 12733 2605 12736
rect 2639 12733 2651 12767
rect 2700 12764 2728 12804
rect 4540 12804 4813 12832
rect 3694 12764 3700 12776
rect 2700 12736 3700 12764
rect 2593 12727 2651 12733
rect 3694 12724 3700 12736
rect 3752 12724 3758 12776
rect 2860 12699 2918 12705
rect 2860 12665 2872 12699
rect 2906 12696 2918 12699
rect 3602 12696 3608 12708
rect 2906 12668 3608 12696
rect 2906 12665 2918 12668
rect 2860 12659 2918 12665
rect 3602 12656 3608 12668
rect 3660 12696 3666 12708
rect 4540 12696 4568 12804
rect 4801 12801 4813 12804
rect 4847 12832 4859 12835
rect 5718 12832 5724 12844
rect 4847 12804 5724 12832
rect 4847 12801 4859 12804
rect 4801 12795 4859 12801
rect 5718 12792 5724 12804
rect 5776 12832 5782 12844
rect 5997 12835 6055 12841
rect 5997 12832 6009 12835
rect 5776 12804 6009 12832
rect 5776 12792 5782 12804
rect 5997 12801 6009 12804
rect 6043 12801 6055 12835
rect 6748 12832 6776 12872
rect 8404 12832 8432 12940
rect 8754 12928 8760 12980
rect 8812 12968 8818 12980
rect 9953 12971 10011 12977
rect 9953 12968 9965 12971
rect 8812 12940 9965 12968
rect 8812 12928 8818 12940
rect 9953 12937 9965 12940
rect 9999 12937 10011 12971
rect 9953 12931 10011 12937
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 10965 12971 11023 12977
rect 10560 12940 10640 12968
rect 10560 12928 10566 12940
rect 8478 12860 8484 12912
rect 8536 12900 8542 12912
rect 8665 12903 8723 12909
rect 8665 12900 8677 12903
rect 8536 12872 8677 12900
rect 8536 12860 8542 12872
rect 8665 12869 8677 12872
rect 8711 12900 8723 12903
rect 9030 12900 9036 12912
rect 8711 12872 9036 12900
rect 8711 12869 8723 12872
rect 8665 12863 8723 12869
rect 9030 12860 9036 12872
rect 9088 12860 9094 12912
rect 9493 12835 9551 12841
rect 9493 12832 9505 12835
rect 6748 12804 7420 12832
rect 8404 12804 9505 12832
rect 5997 12795 6055 12801
rect 4709 12767 4767 12773
rect 4709 12733 4721 12767
rect 4755 12764 4767 12767
rect 6546 12764 6552 12776
rect 4755 12736 6552 12764
rect 4755 12733 4767 12736
rect 4709 12727 4767 12733
rect 6546 12724 6552 12736
rect 6604 12724 6610 12776
rect 6641 12767 6699 12773
rect 6641 12733 6653 12767
rect 6687 12764 6699 12767
rect 7190 12764 7196 12776
rect 6687 12736 7196 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 7285 12767 7343 12773
rect 7285 12733 7297 12767
rect 7331 12733 7343 12767
rect 7392 12764 7420 12804
rect 9493 12801 9505 12804
rect 9539 12832 9551 12835
rect 10502 12832 10508 12844
rect 9539 12804 10508 12832
rect 9539 12801 9551 12804
rect 9493 12795 9551 12801
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 9309 12767 9367 12773
rect 7392 12736 8248 12764
rect 7285 12727 7343 12733
rect 3660 12668 4568 12696
rect 5813 12699 5871 12705
rect 3660 12656 3666 12668
rect 5813 12665 5825 12699
rect 5859 12696 5871 12699
rect 6362 12696 6368 12708
rect 5859 12668 6368 12696
rect 5859 12665 5871 12668
rect 5813 12659 5871 12665
rect 6362 12656 6368 12668
rect 6420 12656 6426 12708
rect 6822 12696 6828 12708
rect 6783 12668 6828 12696
rect 6822 12656 6828 12668
rect 6880 12656 6886 12708
rect 7300 12640 7328 12727
rect 7466 12656 7472 12708
rect 7524 12705 7530 12708
rect 7524 12699 7588 12705
rect 7524 12665 7542 12699
rect 7576 12665 7588 12699
rect 7524 12659 7588 12665
rect 7524 12656 7530 12659
rect 7834 12656 7840 12708
rect 7892 12656 7898 12708
rect 8220 12696 8248 12736
rect 9309 12733 9321 12767
rect 9355 12764 9367 12767
rect 9398 12764 9404 12776
rect 9355 12736 9404 12764
rect 9355 12733 9367 12736
rect 9309 12727 9367 12733
rect 9398 12724 9404 12736
rect 9456 12724 9462 12776
rect 10318 12764 10324 12776
rect 10279 12736 10324 12764
rect 10318 12724 10324 12736
rect 10376 12724 10382 12776
rect 10413 12767 10471 12773
rect 10413 12733 10425 12767
rect 10459 12764 10471 12767
rect 10612 12764 10640 12940
rect 10965 12937 10977 12971
rect 11011 12968 11023 12971
rect 11606 12968 11612 12980
rect 11011 12940 11612 12968
rect 11011 12937 11023 12940
rect 10965 12931 11023 12937
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 12066 12928 12072 12980
rect 12124 12968 12130 12980
rect 12250 12968 12256 12980
rect 12124 12940 12256 12968
rect 12124 12928 12130 12940
rect 12250 12928 12256 12940
rect 12308 12968 12314 12980
rect 14826 12968 14832 12980
rect 12308 12940 14832 12968
rect 12308 12928 12314 12940
rect 14826 12928 14832 12940
rect 14884 12928 14890 12980
rect 14918 12928 14924 12980
rect 14976 12968 14982 12980
rect 15749 12971 15807 12977
rect 14976 12940 15599 12968
rect 14976 12928 14982 12940
rect 11974 12900 11980 12912
rect 11624 12872 11980 12900
rect 11054 12792 11060 12844
rect 11112 12832 11118 12844
rect 11624 12841 11652 12872
rect 11974 12860 11980 12872
rect 12032 12860 12038 12912
rect 12710 12900 12716 12912
rect 12084 12872 12716 12900
rect 11425 12835 11483 12841
rect 11425 12832 11437 12835
rect 11112 12804 11437 12832
rect 11112 12792 11118 12804
rect 11425 12801 11437 12804
rect 11471 12801 11483 12835
rect 11425 12795 11483 12801
rect 11609 12835 11667 12841
rect 11609 12801 11621 12835
rect 11655 12801 11667 12835
rect 11882 12832 11888 12844
rect 11843 12804 11888 12832
rect 11609 12795 11667 12801
rect 11882 12792 11888 12804
rect 11940 12792 11946 12844
rect 10459 12736 10640 12764
rect 10459 12733 10471 12736
rect 10413 12727 10471 12733
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11333 12767 11391 12773
rect 11333 12764 11345 12767
rect 11204 12736 11345 12764
rect 11204 12724 11210 12736
rect 11333 12733 11345 12736
rect 11379 12733 11391 12767
rect 11333 12727 11391 12733
rect 8220 12668 9444 12696
rect 1946 12628 1952 12640
rect 1907 12600 1952 12628
rect 1946 12588 1952 12600
rect 2004 12588 2010 12640
rect 3418 12588 3424 12640
rect 3476 12628 3482 12640
rect 3694 12628 3700 12640
rect 3476 12600 3700 12628
rect 3476 12588 3482 12600
rect 3694 12588 3700 12600
rect 3752 12588 3758 12640
rect 4246 12628 4252 12640
rect 4207 12600 4252 12628
rect 4246 12588 4252 12600
rect 4304 12588 4310 12640
rect 4617 12631 4675 12637
rect 4617 12597 4629 12631
rect 4663 12628 4675 12631
rect 5258 12628 5264 12640
rect 4663 12600 5264 12628
rect 4663 12597 4675 12600
rect 4617 12591 4675 12597
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 5902 12588 5908 12640
rect 5960 12628 5966 12640
rect 5960 12600 6005 12628
rect 5960 12588 5966 12600
rect 6086 12588 6092 12640
rect 6144 12628 6150 12640
rect 6638 12628 6644 12640
rect 6144 12600 6644 12628
rect 6144 12588 6150 12600
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 7282 12628 7288 12640
rect 7195 12600 7288 12628
rect 7282 12588 7288 12600
rect 7340 12628 7346 12640
rect 7852 12628 7880 12656
rect 8294 12628 8300 12640
rect 7340 12600 8300 12628
rect 7340 12588 7346 12600
rect 8294 12588 8300 12600
rect 8352 12588 8358 12640
rect 8938 12628 8944 12640
rect 8899 12600 8944 12628
rect 8938 12588 8944 12600
rect 8996 12588 9002 12640
rect 9416 12637 9444 12668
rect 10870 12656 10876 12708
rect 10928 12696 10934 12708
rect 12084 12696 12112 12872
rect 12710 12860 12716 12872
rect 12768 12860 12774 12912
rect 14093 12903 14151 12909
rect 14093 12869 14105 12903
rect 14139 12900 14151 12903
rect 14182 12900 14188 12912
rect 14139 12872 14188 12900
rect 14139 12869 14151 12872
rect 14093 12863 14151 12869
rect 14182 12860 14188 12872
rect 14240 12860 14246 12912
rect 14369 12903 14427 12909
rect 14369 12869 14381 12903
rect 14415 12900 14427 12903
rect 15194 12900 15200 12912
rect 14415 12872 15200 12900
rect 14415 12869 14427 12872
rect 14369 12863 14427 12869
rect 15194 12860 15200 12872
rect 15252 12860 15258 12912
rect 15289 12903 15347 12909
rect 15289 12869 15301 12903
rect 15335 12900 15347 12903
rect 15470 12900 15476 12912
rect 15335 12872 15476 12900
rect 15335 12869 15347 12872
rect 15289 12863 15347 12869
rect 15470 12860 15476 12872
rect 15528 12860 15534 12912
rect 13814 12792 13820 12844
rect 13872 12832 13878 12844
rect 14967 12835 15025 12841
rect 14967 12832 14979 12835
rect 13872 12804 14979 12832
rect 13872 12792 13878 12804
rect 14967 12801 14979 12804
rect 15013 12801 15025 12835
rect 15571 12832 15599 12940
rect 15749 12937 15761 12971
rect 15795 12968 15807 12971
rect 16022 12968 16028 12980
rect 15795 12940 16028 12968
rect 15795 12937 15807 12940
rect 15749 12931 15807 12937
rect 16022 12928 16028 12940
rect 16080 12928 16086 12980
rect 16301 12971 16359 12977
rect 16301 12937 16313 12971
rect 16347 12968 16359 12971
rect 16482 12968 16488 12980
rect 16347 12940 16488 12968
rect 16347 12937 16359 12940
rect 16301 12931 16359 12937
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 19886 12968 19892 12980
rect 18984 12940 19892 12968
rect 15930 12860 15936 12912
rect 15988 12900 15994 12912
rect 15988 12872 16988 12900
rect 15988 12860 15994 12872
rect 16960 12844 16988 12872
rect 17310 12860 17316 12912
rect 17368 12900 17374 12912
rect 18984 12900 19012 12940
rect 19886 12928 19892 12940
rect 19944 12928 19950 12980
rect 17368 12872 19012 12900
rect 17368 12860 17374 12872
rect 19242 12860 19248 12912
rect 19300 12860 19306 12912
rect 19334 12860 19340 12912
rect 19392 12900 19398 12912
rect 19392 12872 19564 12900
rect 19392 12860 19398 12872
rect 16117 12835 16175 12841
rect 16117 12832 16129 12835
rect 15571 12804 16129 12832
rect 14967 12795 15025 12801
rect 16117 12801 16129 12804
rect 16163 12832 16175 12835
rect 16942 12832 16948 12844
rect 16163 12804 16712 12832
rect 16903 12804 16948 12832
rect 16163 12801 16175 12804
rect 16117 12795 16175 12801
rect 12158 12724 12164 12776
rect 12216 12764 12222 12776
rect 12434 12764 12440 12776
rect 12216 12736 12440 12764
rect 12216 12724 12222 12736
rect 12434 12724 12440 12736
rect 12492 12764 12498 12776
rect 12713 12767 12771 12773
rect 12713 12764 12725 12767
rect 12492 12736 12725 12764
rect 12492 12724 12498 12736
rect 12713 12733 12725 12736
rect 12759 12733 12771 12767
rect 13446 12764 13452 12776
rect 12713 12727 12771 12733
rect 12912 12736 13452 12764
rect 12912 12696 12940 12736
rect 13446 12724 13452 12736
rect 13504 12724 13510 12776
rect 14274 12724 14280 12776
rect 14332 12764 14338 12776
rect 15473 12767 15531 12773
rect 15473 12764 15485 12767
rect 14332 12736 15485 12764
rect 14332 12724 14338 12736
rect 15473 12733 15485 12736
rect 15519 12733 15531 12767
rect 15473 12727 15531 12733
rect 15565 12767 15623 12773
rect 15565 12733 15577 12767
rect 15611 12764 15623 12767
rect 16298 12764 16304 12776
rect 15611 12736 16304 12764
rect 15611 12733 15623 12736
rect 15565 12727 15623 12733
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 16684 12773 16712 12804
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 18598 12832 18604 12844
rect 18064 12804 18604 12832
rect 16669 12767 16727 12773
rect 16669 12733 16681 12767
rect 16715 12733 16727 12767
rect 16669 12727 16727 12733
rect 16758 12724 16764 12776
rect 16816 12764 16822 12776
rect 17405 12767 17463 12773
rect 17405 12764 17417 12767
rect 16816 12736 17417 12764
rect 16816 12724 16822 12736
rect 17405 12733 17417 12736
rect 17451 12733 17463 12767
rect 17405 12727 17463 12733
rect 10928 12668 12112 12696
rect 12728 12668 12940 12696
rect 12980 12699 13038 12705
rect 10928 12656 10934 12668
rect 9401 12631 9459 12637
rect 9401 12597 9413 12631
rect 9447 12628 9459 12631
rect 12728 12628 12756 12668
rect 12980 12665 12992 12699
rect 13026 12696 13038 12699
rect 13354 12696 13360 12708
rect 13026 12668 13360 12696
rect 13026 12665 13038 12668
rect 12980 12659 13038 12665
rect 13354 12656 13360 12668
rect 13412 12656 13418 12708
rect 13538 12656 13544 12708
rect 13596 12696 13602 12708
rect 13906 12696 13912 12708
rect 13596 12668 13912 12696
rect 13596 12656 13602 12668
rect 13906 12656 13912 12668
rect 13964 12656 13970 12708
rect 13998 12656 14004 12708
rect 14056 12696 14062 12708
rect 14918 12696 14924 12708
rect 14056 12668 14924 12696
rect 14056 12656 14062 12668
rect 14918 12656 14924 12668
rect 14976 12656 14982 12708
rect 18064 12696 18092 12804
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 18782 12792 18788 12844
rect 18840 12792 18846 12844
rect 18141 12767 18199 12773
rect 18141 12733 18153 12767
rect 18187 12764 18199 12767
rect 18800 12764 18828 12792
rect 18187 12736 18828 12764
rect 18187 12733 18199 12736
rect 18141 12727 18199 12733
rect 18874 12724 18880 12776
rect 18932 12764 18938 12776
rect 19058 12764 19064 12776
rect 18932 12736 19064 12764
rect 18932 12724 18938 12736
rect 19058 12724 19064 12736
rect 19116 12724 19122 12776
rect 19260 12773 19288 12860
rect 19429 12835 19487 12841
rect 19429 12801 19441 12835
rect 19475 12801 19487 12835
rect 19429 12795 19487 12801
rect 19245 12767 19303 12773
rect 19245 12733 19257 12767
rect 19291 12733 19303 12767
rect 19245 12727 19303 12733
rect 19334 12724 19340 12776
rect 19392 12764 19398 12776
rect 19444 12764 19472 12795
rect 19392 12736 19472 12764
rect 19536 12764 19564 12872
rect 20438 12832 20444 12844
rect 20399 12804 20444 12832
rect 20438 12792 20444 12804
rect 20496 12792 20502 12844
rect 20349 12767 20407 12773
rect 20349 12764 20361 12767
rect 19536 12736 20361 12764
rect 19392 12724 19398 12736
rect 20349 12733 20361 12736
rect 20395 12733 20407 12767
rect 20349 12727 20407 12733
rect 18414 12696 18420 12708
rect 15028 12668 15976 12696
rect 9447 12600 12756 12628
rect 9447 12597 9459 12600
rect 9401 12591 9459 12597
rect 13262 12588 13268 12640
rect 13320 12628 13326 12640
rect 13630 12628 13636 12640
rect 13320 12600 13636 12628
rect 13320 12588 13326 12600
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 14550 12588 14556 12640
rect 14608 12628 14614 12640
rect 14737 12631 14795 12637
rect 14737 12628 14749 12631
rect 14608 12600 14749 12628
rect 14608 12588 14614 12600
rect 14737 12597 14749 12600
rect 14783 12597 14795 12631
rect 14737 12591 14795 12597
rect 14829 12631 14887 12637
rect 14829 12597 14841 12631
rect 14875 12628 14887 12631
rect 15028 12628 15056 12668
rect 14875 12600 15056 12628
rect 15948 12628 15976 12668
rect 16776 12668 18092 12696
rect 18375 12668 18420 12696
rect 16574 12628 16580 12640
rect 15948 12600 16580 12628
rect 14875 12597 14887 12600
rect 14829 12591 14887 12597
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 16776 12637 16804 12668
rect 18414 12656 18420 12668
rect 18472 12656 18478 12708
rect 20257 12699 20315 12705
rect 20257 12696 20269 12699
rect 18892 12668 20269 12696
rect 16761 12631 16819 12637
rect 16761 12597 16773 12631
rect 16807 12597 16819 12631
rect 16761 12591 16819 12597
rect 17589 12631 17647 12637
rect 17589 12597 17601 12631
rect 17635 12628 17647 12631
rect 17954 12628 17960 12640
rect 17635 12600 17960 12628
rect 17635 12597 17647 12600
rect 17589 12591 17647 12597
rect 17954 12588 17960 12600
rect 18012 12588 18018 12640
rect 18892 12637 18920 12668
rect 20257 12665 20269 12668
rect 20303 12665 20315 12699
rect 20257 12659 20315 12665
rect 18877 12631 18935 12637
rect 18877 12597 18889 12631
rect 18923 12597 18935 12631
rect 18877 12591 18935 12597
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 19889 12631 19947 12637
rect 19392 12600 19437 12628
rect 19392 12588 19398 12600
rect 19889 12597 19901 12631
rect 19935 12628 19947 12631
rect 20806 12628 20812 12640
rect 19935 12600 20812 12628
rect 19935 12597 19947 12600
rect 19889 12591 19947 12597
rect 20806 12588 20812 12600
rect 20864 12588 20870 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 1118 12384 1124 12436
rect 1176 12424 1182 12436
rect 1581 12427 1639 12433
rect 1581 12424 1593 12427
rect 1176 12396 1593 12424
rect 1176 12384 1182 12396
rect 1581 12393 1593 12396
rect 1627 12393 1639 12427
rect 1946 12424 1952 12436
rect 1907 12396 1952 12424
rect 1581 12387 1639 12393
rect 1946 12384 1952 12396
rect 2004 12384 2010 12436
rect 2317 12427 2375 12433
rect 2317 12393 2329 12427
rect 2363 12424 2375 12427
rect 2961 12427 3019 12433
rect 2961 12424 2973 12427
rect 2363 12396 2973 12424
rect 2363 12393 2375 12396
rect 2317 12387 2375 12393
rect 2961 12393 2973 12396
rect 3007 12393 3019 12427
rect 2961 12387 3019 12393
rect 3160 12396 3740 12424
rect 2409 12359 2467 12365
rect 2409 12325 2421 12359
rect 2455 12356 2467 12359
rect 3160 12356 3188 12396
rect 2455 12328 3188 12356
rect 2455 12325 2467 12328
rect 2409 12319 2467 12325
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1486 12288 1492 12300
rect 1443 12260 1492 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1486 12248 1492 12260
rect 1544 12248 1550 12300
rect 3329 12291 3387 12297
rect 3329 12257 3341 12291
rect 3375 12288 3387 12291
rect 3510 12288 3516 12300
rect 3375 12260 3516 12288
rect 3375 12257 3387 12260
rect 3329 12251 3387 12257
rect 3510 12248 3516 12260
rect 3568 12248 3574 12300
rect 2590 12220 2596 12232
rect 2551 12192 2596 12220
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 3418 12220 3424 12232
rect 3379 12192 3424 12220
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3602 12220 3608 12232
rect 3563 12192 3608 12220
rect 3602 12180 3608 12192
rect 3660 12180 3666 12232
rect 3712 12220 3740 12396
rect 3878 12384 3884 12436
rect 3936 12424 3942 12436
rect 4249 12427 4307 12433
rect 4249 12424 4261 12427
rect 3936 12396 4261 12424
rect 3936 12384 3942 12396
rect 4249 12393 4261 12396
rect 4295 12393 4307 12427
rect 4249 12387 4307 12393
rect 5718 12384 5724 12436
rect 5776 12424 5782 12436
rect 6089 12427 6147 12433
rect 6089 12424 6101 12427
rect 5776 12396 6101 12424
rect 5776 12384 5782 12396
rect 6089 12393 6101 12396
rect 6135 12393 6147 12427
rect 6089 12387 6147 12393
rect 6733 12427 6791 12433
rect 6733 12393 6745 12427
rect 6779 12424 6791 12427
rect 7098 12424 7104 12436
rect 6779 12396 7104 12424
rect 6779 12393 6791 12396
rect 6733 12387 6791 12393
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 7374 12424 7380 12436
rect 7335 12396 7380 12424
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 7650 12384 7656 12436
rect 7708 12384 7714 12436
rect 8849 12427 8907 12433
rect 8849 12393 8861 12427
rect 8895 12424 8907 12427
rect 8938 12424 8944 12436
rect 8895 12396 8944 12424
rect 8895 12393 8907 12396
rect 8849 12387 8907 12393
rect 8938 12384 8944 12396
rect 8996 12384 9002 12436
rect 10318 12384 10324 12436
rect 10376 12424 10382 12436
rect 10594 12424 10600 12436
rect 10376 12396 10600 12424
rect 10376 12384 10382 12396
rect 10594 12384 10600 12396
rect 10652 12384 10658 12436
rect 10870 12384 10876 12436
rect 10928 12424 10934 12436
rect 11974 12424 11980 12436
rect 10928 12396 11980 12424
rect 10928 12384 10934 12396
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 12986 12384 12992 12436
rect 13044 12424 13050 12436
rect 13081 12427 13139 12433
rect 13081 12424 13093 12427
rect 13044 12396 13093 12424
rect 13044 12384 13050 12396
rect 13081 12393 13093 12396
rect 13127 12393 13139 12427
rect 14090 12424 14096 12436
rect 14051 12396 14096 12424
rect 13081 12387 13139 12393
rect 14090 12384 14096 12396
rect 14148 12384 14154 12436
rect 14461 12427 14519 12433
rect 14461 12393 14473 12427
rect 14507 12424 14519 12427
rect 15746 12424 15752 12436
rect 14507 12396 15752 12424
rect 14507 12393 14519 12396
rect 14461 12387 14519 12393
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 15930 12384 15936 12436
rect 15988 12424 15994 12436
rect 16393 12427 16451 12433
rect 16393 12424 16405 12427
rect 15988 12396 16405 12424
rect 15988 12384 15994 12396
rect 16393 12393 16405 12396
rect 16439 12424 16451 12427
rect 17034 12424 17040 12436
rect 16439 12396 17040 12424
rect 16439 12393 16451 12396
rect 16393 12387 16451 12393
rect 17034 12384 17040 12396
rect 17092 12424 17098 12436
rect 17865 12427 17923 12433
rect 17092 12396 17724 12424
rect 17092 12384 17098 12396
rect 6546 12356 6552 12368
rect 4080 12328 6552 12356
rect 4080 12297 4108 12328
rect 6546 12316 6552 12328
rect 6604 12316 6610 12368
rect 7668 12356 7696 12384
rect 8110 12356 8116 12368
rect 7668 12328 8116 12356
rect 8110 12316 8116 12328
rect 8168 12316 8174 12368
rect 8294 12316 8300 12368
rect 8352 12356 8358 12368
rect 8352 12328 8892 12356
rect 8352 12316 8358 12328
rect 4065 12291 4123 12297
rect 4065 12257 4077 12291
rect 4111 12257 4123 12291
rect 4065 12251 4123 12257
rect 4798 12248 4804 12300
rect 4856 12288 4862 12300
rect 4965 12291 5023 12297
rect 4965 12288 4977 12291
rect 4856 12260 4977 12288
rect 4856 12248 4862 12260
rect 4965 12257 4977 12260
rect 5011 12257 5023 12291
rect 4965 12251 5023 12257
rect 6086 12248 6092 12300
rect 6144 12288 6150 12300
rect 6825 12291 6883 12297
rect 6825 12288 6837 12291
rect 6144 12260 6837 12288
rect 6144 12248 6150 12260
rect 6825 12257 6837 12260
rect 6871 12288 6883 12291
rect 7558 12288 7564 12300
rect 6871 12260 7564 12288
rect 6871 12257 6883 12260
rect 6825 12251 6883 12257
rect 7558 12248 7564 12260
rect 7616 12248 7622 12300
rect 7745 12291 7803 12297
rect 7745 12257 7757 12291
rect 7791 12288 7803 12291
rect 8662 12288 8668 12300
rect 7791 12260 8668 12288
rect 7791 12257 7803 12260
rect 7745 12251 7803 12257
rect 8662 12248 8668 12260
rect 8720 12248 8726 12300
rect 8757 12291 8815 12297
rect 8757 12257 8769 12291
rect 8803 12257 8815 12291
rect 8864 12288 8892 12328
rect 9490 12316 9496 12368
rect 9548 12356 9554 12368
rect 13538 12356 13544 12368
rect 9548 12328 13544 12356
rect 9548 12316 9554 12328
rect 13538 12316 13544 12328
rect 13596 12316 13602 12368
rect 14182 12316 14188 12368
rect 14240 12356 14246 12368
rect 15841 12359 15899 12365
rect 15841 12356 15853 12359
rect 14240 12328 15853 12356
rect 14240 12316 14246 12328
rect 15841 12325 15853 12328
rect 15887 12325 15899 12359
rect 17696 12356 17724 12396
rect 17865 12393 17877 12427
rect 17911 12424 17923 12427
rect 18874 12424 18880 12436
rect 17911 12396 18880 12424
rect 17911 12393 17923 12396
rect 17865 12387 17923 12393
rect 18874 12384 18880 12396
rect 18932 12384 18938 12436
rect 18966 12384 18972 12436
rect 19024 12424 19030 12436
rect 19334 12424 19340 12436
rect 19024 12396 19340 12424
rect 19024 12384 19030 12396
rect 19334 12384 19340 12396
rect 19392 12384 19398 12436
rect 17954 12356 17960 12368
rect 15841 12319 15899 12325
rect 15948 12328 17632 12356
rect 17696 12328 17960 12356
rect 9769 12291 9827 12297
rect 9769 12288 9781 12291
rect 8864 12260 9781 12288
rect 8757 12251 8815 12257
rect 9769 12257 9781 12260
rect 9815 12257 9827 12291
rect 9769 12251 9827 12257
rect 10036 12291 10094 12297
rect 10036 12257 10048 12291
rect 10082 12288 10094 12291
rect 11054 12288 11060 12300
rect 10082 12260 11060 12288
rect 10082 12257 10094 12260
rect 10036 12251 10094 12257
rect 4246 12220 4252 12232
rect 3712 12192 4252 12220
rect 4246 12180 4252 12192
rect 4304 12180 4310 12232
rect 4338 12180 4344 12232
rect 4396 12220 4402 12232
rect 4709 12223 4767 12229
rect 4709 12220 4721 12223
rect 4396 12192 4721 12220
rect 4396 12180 4402 12192
rect 4709 12189 4721 12192
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 6914 12180 6920 12232
rect 6972 12220 6978 12232
rect 7834 12220 7840 12232
rect 6972 12192 7017 12220
rect 7795 12192 7840 12220
rect 6972 12180 6978 12192
rect 7834 12180 7840 12192
rect 7892 12180 7898 12232
rect 7929 12223 7987 12229
rect 7929 12189 7941 12223
rect 7975 12189 7987 12223
rect 8772 12220 8800 12251
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 11692 12291 11750 12297
rect 11692 12288 11704 12291
rect 11348 12260 11704 12288
rect 8846 12220 8852 12232
rect 8772 12192 8852 12220
rect 7929 12183 7987 12189
rect 5902 12112 5908 12164
rect 5960 12152 5966 12164
rect 6365 12155 6423 12161
rect 6365 12152 6377 12155
rect 5960 12124 6377 12152
rect 5960 12112 5966 12124
rect 6365 12121 6377 12124
rect 6411 12121 6423 12155
rect 6365 12115 6423 12121
rect 7098 12112 7104 12164
rect 7156 12152 7162 12164
rect 7944 12152 7972 12183
rect 8846 12180 8852 12192
rect 8904 12180 8910 12232
rect 9030 12220 9036 12232
rect 8991 12192 9036 12220
rect 9030 12180 9036 12192
rect 9088 12180 9094 12232
rect 9766 12152 9772 12164
rect 7156 12124 7972 12152
rect 8016 12124 9772 12152
rect 7156 12112 7162 12124
rect 4706 12044 4712 12096
rect 4764 12084 4770 12096
rect 8016 12084 8044 12124
rect 9766 12112 9772 12124
rect 9824 12112 9830 12164
rect 11149 12155 11207 12161
rect 11149 12121 11161 12155
rect 11195 12152 11207 12155
rect 11348 12152 11376 12260
rect 11692 12257 11704 12260
rect 11738 12288 11750 12291
rect 12710 12288 12716 12300
rect 11738 12260 12716 12288
rect 11738 12257 11750 12260
rect 11692 12251 11750 12257
rect 12710 12248 12716 12260
rect 12768 12248 12774 12300
rect 13449 12291 13507 12297
rect 13449 12257 13461 12291
rect 13495 12288 13507 12291
rect 13814 12288 13820 12300
rect 13495 12260 13820 12288
rect 13495 12257 13507 12260
rect 13449 12251 13507 12257
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 13906 12248 13912 12300
rect 13964 12288 13970 12300
rect 15948 12288 15976 12328
rect 16752 12291 16810 12297
rect 16752 12288 16764 12291
rect 13964 12260 14688 12288
rect 13964 12248 13970 12260
rect 11425 12223 11483 12229
rect 11425 12189 11437 12223
rect 11471 12189 11483 12223
rect 13538 12220 13544 12232
rect 13499 12192 13544 12220
rect 11425 12183 11483 12189
rect 11195 12124 11376 12152
rect 11195 12121 11207 12124
rect 11149 12115 11207 12121
rect 4764 12056 8044 12084
rect 4764 12044 4770 12056
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 8389 12087 8447 12093
rect 8389 12084 8401 12087
rect 8260 12056 8401 12084
rect 8260 12044 8266 12056
rect 8389 12053 8401 12056
rect 8435 12053 8447 12087
rect 8389 12047 8447 12053
rect 8570 12044 8576 12096
rect 8628 12084 8634 12096
rect 10962 12084 10968 12096
rect 8628 12056 10968 12084
rect 8628 12044 8634 12056
rect 10962 12044 10968 12056
rect 11020 12044 11026 12096
rect 11440 12084 11468 12183
rect 13538 12180 13544 12192
rect 13596 12180 13602 12232
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12220 13783 12223
rect 13924 12220 13952 12248
rect 13771 12192 13952 12220
rect 13771 12189 13783 12192
rect 13725 12183 13783 12189
rect 14366 12180 14372 12232
rect 14424 12220 14430 12232
rect 14660 12229 14688 12260
rect 14752 12260 15976 12288
rect 16132 12260 16764 12288
rect 14553 12223 14611 12229
rect 14553 12220 14565 12223
rect 14424 12192 14565 12220
rect 14424 12180 14430 12192
rect 14553 12189 14565 12192
rect 14599 12189 14611 12223
rect 14553 12183 14611 12189
rect 14645 12223 14703 12229
rect 14645 12189 14657 12223
rect 14691 12189 14703 12223
rect 14645 12183 14703 12189
rect 13078 12112 13084 12164
rect 13136 12152 13142 12164
rect 13630 12152 13636 12164
rect 13136 12124 13636 12152
rect 13136 12112 13142 12124
rect 13630 12112 13636 12124
rect 13688 12112 13694 12164
rect 14182 12112 14188 12164
rect 14240 12152 14246 12164
rect 14752 12152 14780 12260
rect 14826 12180 14832 12232
rect 14884 12220 14890 12232
rect 15378 12220 15384 12232
rect 14884 12192 15384 12220
rect 14884 12180 14890 12192
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 16132 12229 16160 12260
rect 16752 12257 16764 12260
rect 16798 12288 16810 12291
rect 17494 12288 17500 12300
rect 16798 12260 17500 12288
rect 16798 12257 16810 12260
rect 16752 12251 16810 12257
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 17604 12288 17632 12328
rect 17954 12316 17960 12328
rect 18012 12356 18018 12368
rect 18012 12328 18276 12356
rect 18012 12316 18018 12328
rect 17770 12288 17776 12300
rect 17604 12260 17776 12288
rect 17770 12248 17776 12260
rect 17828 12248 17834 12300
rect 18248 12297 18276 12328
rect 19242 12316 19248 12368
rect 19300 12356 19306 12368
rect 19797 12359 19855 12365
rect 19797 12356 19809 12359
rect 19300 12328 19809 12356
rect 19300 12316 19306 12328
rect 19797 12325 19809 12328
rect 19843 12325 19855 12359
rect 19797 12319 19855 12325
rect 20165 12359 20223 12365
rect 20165 12325 20177 12359
rect 20211 12356 20223 12359
rect 20898 12356 20904 12368
rect 20211 12328 20904 12356
rect 20211 12325 20223 12328
rect 20165 12319 20223 12325
rect 20898 12316 20904 12328
rect 20956 12316 20962 12368
rect 18233 12291 18291 12297
rect 18233 12257 18245 12291
rect 18279 12257 18291 12291
rect 18233 12251 18291 12257
rect 18500 12291 18558 12297
rect 18500 12257 18512 12291
rect 18546 12288 18558 12291
rect 18966 12288 18972 12300
rect 18546 12260 18972 12288
rect 18546 12257 18558 12260
rect 18500 12251 18558 12257
rect 18966 12248 18972 12260
rect 19024 12288 19030 12300
rect 19889 12291 19947 12297
rect 19024 12260 19288 12288
rect 19024 12248 19030 12260
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 15764 12192 15945 12220
rect 14240 12124 14780 12152
rect 14240 12112 14246 12124
rect 14918 12112 14924 12164
rect 14976 12152 14982 12164
rect 15102 12152 15108 12164
rect 14976 12124 15108 12152
rect 14976 12112 14982 12124
rect 15102 12112 15108 12124
rect 15160 12112 15166 12164
rect 15562 12152 15568 12164
rect 15396 12124 15568 12152
rect 12434 12084 12440 12096
rect 11440 12056 12440 12084
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 12618 12044 12624 12096
rect 12676 12084 12682 12096
rect 12805 12087 12863 12093
rect 12805 12084 12817 12087
rect 12676 12056 12817 12084
rect 12676 12044 12682 12056
rect 12805 12053 12817 12056
rect 12851 12053 12863 12087
rect 12805 12047 12863 12053
rect 12986 12044 12992 12096
rect 13044 12084 13050 12096
rect 15396 12084 15424 12124
rect 15562 12112 15568 12124
rect 15620 12152 15626 12164
rect 15764 12152 15792 12192
rect 15933 12189 15945 12192
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 16117 12223 16175 12229
rect 16117 12189 16129 12223
rect 16163 12189 16175 12223
rect 16117 12183 16175 12189
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12220 16451 12223
rect 16485 12223 16543 12229
rect 16485 12220 16497 12223
rect 16439 12192 16497 12220
rect 16439 12189 16451 12192
rect 16393 12183 16451 12189
rect 16485 12189 16497 12192
rect 16531 12189 16543 12223
rect 19260 12220 19288 12260
rect 19889 12257 19901 12291
rect 19935 12288 19947 12291
rect 20530 12288 20536 12300
rect 19935 12260 20536 12288
rect 19935 12257 19947 12260
rect 19889 12251 19947 12257
rect 20530 12248 20536 12260
rect 20588 12248 20594 12300
rect 20438 12220 20444 12232
rect 19260 12192 20444 12220
rect 16485 12183 16543 12189
rect 20438 12180 20444 12192
rect 20496 12180 20502 12232
rect 20901 12223 20959 12229
rect 20901 12189 20913 12223
rect 20947 12189 20959 12223
rect 20901 12183 20959 12189
rect 15620 12124 15792 12152
rect 15620 12112 15626 12124
rect 15838 12112 15844 12164
rect 15896 12152 15902 12164
rect 19797 12155 19855 12161
rect 15896 12124 16528 12152
rect 15896 12112 15902 12124
rect 13044 12056 15424 12084
rect 15473 12087 15531 12093
rect 13044 12044 13050 12056
rect 15473 12053 15485 12087
rect 15519 12084 15531 12087
rect 16206 12084 16212 12096
rect 15519 12056 16212 12084
rect 15519 12053 15531 12056
rect 15473 12047 15531 12053
rect 16206 12044 16212 12056
rect 16264 12044 16270 12096
rect 16500 12084 16528 12124
rect 19168 12124 19748 12152
rect 19168 12084 19196 12124
rect 19720 12096 19748 12124
rect 19797 12121 19809 12155
rect 19843 12152 19855 12155
rect 20916 12152 20944 12183
rect 19843 12124 20944 12152
rect 19843 12121 19855 12124
rect 19797 12115 19855 12121
rect 16500 12056 19196 12084
rect 19242 12044 19248 12096
rect 19300 12084 19306 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 19300 12056 19625 12084
rect 19300 12044 19306 12056
rect 19613 12053 19625 12056
rect 19659 12053 19671 12087
rect 19613 12047 19671 12053
rect 19702 12044 19708 12096
rect 19760 12044 19766 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 3234 11840 3240 11892
rect 3292 11880 3298 11892
rect 3602 11880 3608 11892
rect 3292 11852 3608 11880
rect 3292 11840 3298 11852
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 4154 11840 4160 11892
rect 4212 11880 4218 11892
rect 5077 11883 5135 11889
rect 5077 11880 5089 11883
rect 4212 11852 5089 11880
rect 4212 11840 4218 11852
rect 5077 11849 5089 11852
rect 5123 11849 5135 11883
rect 5077 11843 5135 11849
rect 5537 11883 5595 11889
rect 5537 11849 5549 11883
rect 5583 11880 5595 11883
rect 5626 11880 5632 11892
rect 5583 11852 5632 11880
rect 5583 11849 5595 11852
rect 5537 11843 5595 11849
rect 5626 11840 5632 11852
rect 5684 11840 5690 11892
rect 6362 11840 6368 11892
rect 6420 11880 6426 11892
rect 6825 11883 6883 11889
rect 6825 11880 6837 11883
rect 6420 11852 6837 11880
rect 6420 11840 6426 11852
rect 6825 11849 6837 11852
rect 6871 11849 6883 11883
rect 6825 11843 6883 11849
rect 7374 11840 7380 11892
rect 7432 11840 7438 11892
rect 7834 11880 7840 11892
rect 7795 11852 7840 11880
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 8386 11840 8392 11892
rect 8444 11880 8450 11892
rect 8570 11880 8576 11892
rect 8444 11852 8576 11880
rect 8444 11840 8450 11852
rect 8570 11840 8576 11852
rect 8628 11840 8634 11892
rect 9030 11880 9036 11892
rect 8991 11852 9036 11880
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 9858 11880 9864 11892
rect 9819 11852 9864 11880
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 12250 11880 12256 11892
rect 9968 11852 12256 11880
rect 2133 11815 2191 11821
rect 2133 11781 2145 11815
rect 2179 11781 2191 11815
rect 2133 11775 2191 11781
rect 4617 11815 4675 11821
rect 4617 11781 4629 11815
rect 4663 11812 4675 11815
rect 4798 11812 4804 11824
rect 4663 11784 4804 11812
rect 4663 11781 4675 11784
rect 4617 11775 4675 11781
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 2148 11676 2176 11775
rect 4798 11772 4804 11784
rect 4856 11812 4862 11824
rect 7392 11812 7420 11840
rect 7926 11812 7932 11824
rect 4856 11784 6132 11812
rect 7392 11784 7932 11812
rect 4856 11772 4862 11784
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11744 2835 11747
rect 2823 11716 3372 11744
rect 2823 11713 2835 11716
rect 2777 11707 2835 11713
rect 3344 11688 3372 11716
rect 5350 11704 5356 11756
rect 5408 11744 5414 11756
rect 6104 11753 6132 11784
rect 7926 11772 7932 11784
rect 7984 11812 7990 11824
rect 7984 11784 9260 11812
rect 7984 11772 7990 11784
rect 6089 11747 6147 11753
rect 5408 11716 5948 11744
rect 5408 11704 5414 11716
rect 1443 11648 2176 11676
rect 3237 11679 3295 11685
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 3237 11645 3249 11679
rect 3283 11645 3295 11679
rect 3237 11639 3295 11645
rect 1670 11608 1676 11620
rect 1631 11580 1676 11608
rect 1670 11568 1676 11580
rect 1728 11568 1734 11620
rect 1854 11568 1860 11620
rect 1912 11608 1918 11620
rect 2406 11608 2412 11620
rect 1912 11580 2412 11608
rect 1912 11568 1918 11580
rect 2406 11568 2412 11580
rect 2464 11608 2470 11620
rect 3252 11608 3280 11639
rect 3326 11636 3332 11688
rect 3384 11676 3390 11688
rect 3493 11679 3551 11685
rect 3493 11676 3505 11679
rect 3384 11648 3505 11676
rect 3384 11636 3390 11648
rect 3493 11645 3505 11648
rect 3539 11645 3551 11679
rect 4890 11676 4896 11688
rect 4851 11648 4896 11676
rect 3493 11639 3551 11645
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 5920 11685 5948 11716
rect 6089 11713 6101 11747
rect 6135 11744 6147 11747
rect 6914 11744 6920 11756
rect 6135 11716 6920 11744
rect 6135 11713 6147 11716
rect 6089 11707 6147 11713
rect 6914 11704 6920 11716
rect 6972 11744 6978 11756
rect 7377 11747 7435 11753
rect 7377 11744 7389 11747
rect 6972 11716 7389 11744
rect 6972 11704 6978 11716
rect 7377 11713 7389 11716
rect 7423 11713 7435 11747
rect 7377 11707 7435 11713
rect 8110 11704 8116 11756
rect 8168 11744 8174 11756
rect 8297 11747 8355 11753
rect 8297 11744 8309 11747
rect 8168 11716 8309 11744
rect 8168 11704 8174 11716
rect 8297 11713 8309 11716
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 8386 11704 8392 11756
rect 8444 11744 8450 11756
rect 9232 11744 9260 11784
rect 9306 11772 9312 11824
rect 9364 11812 9370 11824
rect 9968 11812 9996 11852
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 12710 11840 12716 11892
rect 12768 11880 12774 11892
rect 15749 11883 15807 11889
rect 12768 11852 15332 11880
rect 12768 11840 12774 11852
rect 11517 11815 11575 11821
rect 9364 11784 9996 11812
rect 10060 11784 11376 11812
rect 9364 11772 9370 11784
rect 9585 11747 9643 11753
rect 9585 11744 9597 11747
rect 8444 11716 8489 11744
rect 9232 11716 9597 11744
rect 8444 11704 8450 11716
rect 9585 11713 9597 11716
rect 9631 11744 9643 11747
rect 10060 11744 10088 11784
rect 10502 11744 10508 11756
rect 9631 11716 10088 11744
rect 10463 11716 10508 11744
rect 9631 11713 9643 11716
rect 9585 11707 9643 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10962 11704 10968 11756
rect 11020 11704 11026 11756
rect 11241 11747 11299 11753
rect 11241 11713 11253 11747
rect 11287 11713 11299 11747
rect 11348 11744 11376 11784
rect 11517 11781 11529 11815
rect 11563 11812 11575 11815
rect 11974 11812 11980 11824
rect 11563 11784 11980 11812
rect 11563 11781 11575 11784
rect 11517 11775 11575 11781
rect 11974 11772 11980 11784
rect 12032 11772 12038 11824
rect 13817 11815 13875 11821
rect 13817 11781 13829 11815
rect 13863 11812 13875 11815
rect 13906 11812 13912 11824
rect 13863 11784 13912 11812
rect 13863 11781 13875 11784
rect 13817 11775 13875 11781
rect 13906 11772 13912 11784
rect 13964 11772 13970 11824
rect 14093 11815 14151 11821
rect 14093 11781 14105 11815
rect 14139 11812 14151 11815
rect 14274 11812 14280 11824
rect 14139 11784 14280 11812
rect 14139 11781 14151 11784
rect 14093 11775 14151 11781
rect 14274 11772 14280 11784
rect 14332 11772 14338 11824
rect 15304 11812 15332 11852
rect 15749 11849 15761 11883
rect 15795 11880 15807 11883
rect 15838 11880 15844 11892
rect 15795 11852 15844 11880
rect 15795 11849 15807 11852
rect 15749 11843 15807 11849
rect 15838 11840 15844 11852
rect 15896 11840 15902 11892
rect 15930 11840 15936 11892
rect 15988 11880 15994 11892
rect 16025 11883 16083 11889
rect 16025 11880 16037 11883
rect 15988 11852 16037 11880
rect 15988 11840 15994 11852
rect 16025 11849 16037 11852
rect 16071 11849 16083 11883
rect 16025 11843 16083 11849
rect 16206 11840 16212 11892
rect 16264 11880 16270 11892
rect 16301 11883 16359 11889
rect 16301 11880 16313 11883
rect 16264 11852 16313 11880
rect 16264 11840 16270 11852
rect 16301 11849 16313 11852
rect 16347 11849 16359 11883
rect 16301 11843 16359 11849
rect 16577 11883 16635 11889
rect 16577 11849 16589 11883
rect 16623 11880 16635 11883
rect 17678 11880 17684 11892
rect 16623 11852 17684 11880
rect 16623 11849 16635 11852
rect 16577 11843 16635 11849
rect 17678 11840 17684 11852
rect 17736 11840 17742 11892
rect 17770 11840 17776 11892
rect 17828 11880 17834 11892
rect 19429 11883 19487 11889
rect 17828 11852 19380 11880
rect 17828 11840 17834 11852
rect 17310 11812 17316 11824
rect 15304 11784 17316 11812
rect 17310 11772 17316 11784
rect 17368 11772 17374 11824
rect 19352 11812 19380 11852
rect 19429 11849 19441 11883
rect 19475 11880 19487 11883
rect 20438 11880 20444 11892
rect 19475 11852 20444 11880
rect 19475 11849 19487 11852
rect 19429 11843 19487 11849
rect 20438 11840 20444 11852
rect 20496 11840 20502 11892
rect 20901 11883 20959 11889
rect 20901 11849 20913 11883
rect 20947 11880 20959 11883
rect 21174 11880 21180 11892
rect 20947 11852 21180 11880
rect 20947 11849 20959 11852
rect 20901 11843 20959 11849
rect 21174 11840 21180 11852
rect 21232 11840 21238 11892
rect 19521 11815 19579 11821
rect 19521 11812 19533 11815
rect 19352 11784 19533 11812
rect 19521 11781 19533 11784
rect 19567 11781 19579 11815
rect 19702 11812 19708 11824
rect 19663 11784 19708 11812
rect 19521 11775 19579 11781
rect 19702 11772 19708 11784
rect 19760 11772 19766 11824
rect 20806 11812 20812 11824
rect 20364 11784 20812 11812
rect 11698 11744 11704 11756
rect 11348 11716 11704 11744
rect 11241 11707 11299 11713
rect 5905 11679 5963 11685
rect 5905 11645 5917 11679
rect 5951 11645 5963 11679
rect 5905 11639 5963 11645
rect 7193 11679 7251 11685
rect 7193 11645 7205 11679
rect 7239 11676 7251 11679
rect 7834 11676 7840 11688
rect 7239 11648 7840 11676
rect 7239 11645 7251 11648
rect 7193 11639 7251 11645
rect 7834 11636 7840 11648
rect 7892 11636 7898 11688
rect 8202 11676 8208 11688
rect 8163 11648 8208 11676
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 10321 11679 10379 11685
rect 10321 11645 10333 11679
rect 10367 11676 10379 11679
rect 10686 11676 10692 11688
rect 10367 11648 10692 11676
rect 10367 11645 10379 11648
rect 10321 11639 10379 11645
rect 10686 11636 10692 11648
rect 10744 11636 10750 11688
rect 4246 11608 4252 11620
rect 2464 11580 4252 11608
rect 2464 11568 2470 11580
rect 4246 11568 4252 11580
rect 4304 11608 4310 11620
rect 5718 11608 5724 11620
rect 4304 11580 5724 11608
rect 4304 11568 4310 11580
rect 5718 11568 5724 11580
rect 5776 11568 5782 11620
rect 9401 11611 9459 11617
rect 9401 11608 9413 11611
rect 6840 11580 9413 11608
rect 6840 11552 6868 11580
rect 9401 11577 9413 11580
rect 9447 11577 9459 11611
rect 9401 11571 9459 11577
rect 9493 11611 9551 11617
rect 9493 11577 9505 11611
rect 9539 11608 9551 11611
rect 10778 11608 10784 11620
rect 9539 11580 10784 11608
rect 9539 11577 9551 11580
rect 9493 11571 9551 11577
rect 10778 11568 10784 11580
rect 10836 11568 10842 11620
rect 10980 11608 11008 11704
rect 11057 11679 11115 11685
rect 11057 11645 11069 11679
rect 11103 11676 11115 11679
rect 11146 11676 11152 11688
rect 11103 11648 11152 11676
rect 11103 11645 11115 11648
rect 11057 11639 11115 11645
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 11256 11676 11284 11707
rect 11698 11704 11704 11716
rect 11756 11704 11762 11756
rect 11882 11744 11888 11756
rect 11808 11716 11888 11744
rect 11808 11676 11836 11716
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11744 12219 11747
rect 12207 11716 12388 11744
rect 12207 11713 12219 11716
rect 12161 11707 12219 11713
rect 11256 11648 11836 11676
rect 12360 11676 12388 11716
rect 12434 11704 12440 11756
rect 12492 11744 12498 11756
rect 14182 11744 14188 11756
rect 12492 11716 12537 11744
rect 13924 11716 14188 11744
rect 12492 11704 12498 11716
rect 12710 11685 12716 11688
rect 12704 11676 12716 11685
rect 12360 11648 12716 11676
rect 12704 11639 12716 11648
rect 12710 11636 12716 11639
rect 12768 11636 12774 11688
rect 12986 11636 12992 11688
rect 13044 11676 13050 11688
rect 13924 11676 13952 11716
rect 14182 11704 14188 11716
rect 14240 11704 14246 11756
rect 15378 11704 15384 11756
rect 15436 11744 15442 11756
rect 15838 11744 15844 11756
rect 15436 11716 15844 11744
rect 15436 11704 15442 11716
rect 15838 11704 15844 11716
rect 15896 11704 15902 11756
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 17405 11747 17463 11753
rect 17405 11744 17417 11747
rect 16347 11716 17417 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 17405 11713 17417 11716
rect 17451 11713 17463 11747
rect 17405 11707 17463 11713
rect 17589 11747 17647 11753
rect 17589 11713 17601 11747
rect 17635 11744 17647 11747
rect 17635 11716 18184 11744
rect 17635 11713 17647 11716
rect 17589 11707 17647 11713
rect 13044 11648 13952 11676
rect 14277 11679 14335 11685
rect 13044 11636 13050 11648
rect 14277 11645 14289 11679
rect 14323 11645 14335 11679
rect 14277 11639 14335 11645
rect 14369 11679 14427 11685
rect 14369 11645 14381 11679
rect 14415 11676 14427 11679
rect 15930 11676 15936 11688
rect 14415 11648 15936 11676
rect 14415 11645 14427 11648
rect 14369 11639 14427 11645
rect 13722 11608 13728 11620
rect 10980 11580 13728 11608
rect 1946 11500 1952 11552
rect 2004 11540 2010 11552
rect 2501 11543 2559 11549
rect 2501 11540 2513 11543
rect 2004 11512 2513 11540
rect 2004 11500 2010 11512
rect 2501 11509 2513 11512
rect 2547 11509 2559 11543
rect 2501 11503 2559 11509
rect 2593 11543 2651 11549
rect 2593 11509 2605 11543
rect 2639 11540 2651 11543
rect 4062 11540 4068 11552
rect 2639 11512 4068 11540
rect 2639 11509 2651 11512
rect 2593 11503 2651 11509
rect 4062 11500 4068 11512
rect 4120 11500 4126 11552
rect 5902 11500 5908 11552
rect 5960 11540 5966 11552
rect 5997 11543 6055 11549
rect 5997 11540 6009 11543
rect 5960 11512 6009 11540
rect 5960 11500 5966 11512
rect 5997 11509 6009 11512
rect 6043 11540 6055 11543
rect 6178 11540 6184 11552
rect 6043 11512 6184 11540
rect 6043 11509 6055 11512
rect 5997 11503 6055 11509
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 6822 11500 6828 11552
rect 6880 11500 6886 11552
rect 7285 11543 7343 11549
rect 7285 11509 7297 11543
rect 7331 11540 7343 11543
rect 9122 11540 9128 11552
rect 7331 11512 9128 11540
rect 7331 11509 7343 11512
rect 7285 11503 7343 11509
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 10042 11500 10048 11552
rect 10100 11540 10106 11552
rect 10229 11543 10287 11549
rect 10229 11540 10241 11543
rect 10100 11512 10241 11540
rect 10100 11500 10106 11512
rect 10229 11509 10241 11512
rect 10275 11509 10287 11543
rect 10229 11503 10287 11509
rect 10689 11543 10747 11549
rect 10689 11509 10701 11543
rect 10735 11540 10747 11543
rect 10870 11540 10876 11552
rect 10735 11512 10876 11540
rect 10735 11509 10747 11512
rect 10689 11503 10747 11509
rect 10870 11500 10876 11512
rect 10928 11500 10934 11552
rect 11164 11549 11192 11580
rect 13722 11568 13728 11580
rect 13780 11568 13786 11620
rect 14182 11568 14188 11620
rect 14240 11608 14246 11620
rect 14292 11608 14320 11639
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 16022 11636 16028 11688
rect 16080 11676 16086 11688
rect 16209 11679 16267 11685
rect 16209 11676 16221 11679
rect 16080 11648 16221 11676
rect 16080 11636 16086 11648
rect 16209 11645 16221 11648
rect 16255 11645 16267 11679
rect 16390 11676 16396 11688
rect 16351 11648 16396 11676
rect 16209 11639 16267 11645
rect 16390 11636 16396 11648
rect 16448 11636 16454 11688
rect 17218 11636 17224 11688
rect 17276 11676 17282 11688
rect 17604 11676 17632 11707
rect 17276 11648 17632 11676
rect 17276 11636 17282 11648
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 18012 11648 18061 11676
rect 18012 11636 18018 11648
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 18156 11676 18184 11716
rect 19242 11704 19248 11756
rect 19300 11744 19306 11756
rect 20257 11747 20315 11753
rect 20257 11744 20269 11747
rect 19300 11716 20269 11744
rect 19300 11704 19306 11716
rect 20257 11713 20269 11716
rect 20303 11713 20315 11747
rect 20257 11707 20315 11713
rect 18316 11679 18374 11685
rect 18316 11676 18328 11679
rect 18156 11648 18328 11676
rect 18049 11639 18107 11645
rect 18316 11645 18328 11648
rect 18362 11676 18374 11679
rect 18874 11676 18880 11688
rect 18362 11648 18880 11676
rect 18362 11645 18374 11648
rect 18316 11639 18374 11645
rect 18874 11636 18880 11648
rect 18932 11636 18938 11688
rect 20073 11679 20131 11685
rect 20073 11645 20085 11679
rect 20119 11676 20131 11679
rect 20364 11676 20392 11784
rect 20806 11772 20812 11784
rect 20864 11772 20870 11824
rect 20119 11648 20392 11676
rect 20717 11679 20775 11685
rect 20119 11645 20131 11648
rect 20073 11639 20131 11645
rect 20717 11645 20729 11679
rect 20763 11676 20775 11679
rect 20806 11676 20812 11688
rect 20763 11648 20812 11676
rect 20763 11645 20775 11648
rect 20717 11639 20775 11645
rect 20806 11636 20812 11648
rect 20864 11636 20870 11688
rect 14642 11617 14648 11620
rect 14240 11580 14320 11608
rect 14625 11611 14648 11617
rect 14240 11568 14246 11580
rect 14625 11577 14637 11611
rect 14625 11571 14648 11577
rect 14642 11568 14648 11571
rect 14700 11568 14706 11620
rect 14826 11568 14832 11620
rect 14884 11568 14890 11620
rect 18414 11568 18420 11620
rect 18472 11608 18478 11620
rect 20165 11611 20223 11617
rect 20165 11608 20177 11611
rect 18472 11580 20177 11608
rect 18472 11568 18478 11580
rect 20165 11577 20177 11580
rect 20211 11577 20223 11611
rect 20165 11571 20223 11577
rect 11149 11543 11207 11549
rect 11149 11509 11161 11543
rect 11195 11509 11207 11543
rect 11149 11503 11207 11509
rect 11790 11500 11796 11552
rect 11848 11540 11854 11552
rect 11885 11543 11943 11549
rect 11885 11540 11897 11543
rect 11848 11512 11897 11540
rect 11848 11500 11854 11512
rect 11885 11509 11897 11512
rect 11931 11509 11943 11543
rect 11885 11503 11943 11509
rect 11977 11543 12035 11549
rect 11977 11509 11989 11543
rect 12023 11540 12035 11543
rect 14844 11540 14872 11568
rect 12023 11512 14872 11540
rect 12023 11509 12035 11512
rect 11977 11503 12035 11509
rect 15102 11500 15108 11552
rect 15160 11540 15166 11552
rect 16758 11540 16764 11552
rect 15160 11512 16764 11540
rect 15160 11500 15166 11512
rect 16758 11500 16764 11512
rect 16816 11500 16822 11552
rect 16945 11543 17003 11549
rect 16945 11509 16957 11543
rect 16991 11540 17003 11543
rect 17126 11540 17132 11552
rect 16991 11512 17132 11540
rect 16991 11509 17003 11512
rect 16945 11503 17003 11509
rect 17126 11500 17132 11512
rect 17184 11500 17190 11552
rect 17310 11540 17316 11552
rect 17271 11512 17316 11540
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 17402 11500 17408 11552
rect 17460 11540 17466 11552
rect 19426 11540 19432 11552
rect 17460 11512 19432 11540
rect 17460 11500 17466 11512
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 19521 11543 19579 11549
rect 19521 11509 19533 11543
rect 19567 11540 19579 11543
rect 20530 11540 20536 11552
rect 19567 11512 20536 11540
rect 19567 11509 19579 11512
rect 19521 11503 19579 11509
rect 20530 11500 20536 11512
rect 20588 11500 20594 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 3237 11339 3295 11345
rect 3237 11305 3249 11339
rect 3283 11336 3295 11339
rect 3326 11336 3332 11348
rect 3283 11308 3332 11336
rect 3283 11305 3295 11308
rect 3237 11299 3295 11305
rect 3326 11296 3332 11308
rect 3384 11296 3390 11348
rect 3510 11336 3516 11348
rect 3471 11308 3516 11336
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 4062 11336 4068 11348
rect 4023 11308 4068 11336
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 4154 11296 4160 11348
rect 4212 11336 4218 11348
rect 5261 11339 5319 11345
rect 5261 11336 5273 11339
rect 4212 11308 5273 11336
rect 4212 11296 4218 11308
rect 5261 11305 5273 11308
rect 5307 11305 5319 11339
rect 8294 11336 8300 11348
rect 5261 11299 5319 11305
rect 5460 11308 8300 11336
rect 3878 11228 3884 11280
rect 3936 11268 3942 11280
rect 4706 11268 4712 11280
rect 3936 11240 4712 11268
rect 3936 11228 3942 11240
rect 4706 11228 4712 11240
rect 4764 11228 4770 11280
rect 1854 11200 1860 11212
rect 1815 11172 1860 11200
rect 1854 11160 1860 11172
rect 1912 11160 1918 11212
rect 2124 11203 2182 11209
rect 2124 11169 2136 11203
rect 2170 11200 2182 11203
rect 2682 11200 2688 11212
rect 2170 11172 2688 11200
rect 2170 11169 2182 11172
rect 2124 11163 2182 11169
rect 2682 11160 2688 11172
rect 2740 11200 2746 11212
rect 2740 11172 3280 11200
rect 2740 11160 2746 11172
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11101 1455 11135
rect 1397 11095 1455 11101
rect 1412 10996 1440 11095
rect 3252 11076 3280 11172
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4212 11172 4445 11200
rect 4212 11160 4218 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 5074 11200 5080 11212
rect 5035 11172 5080 11200
rect 4433 11163 4491 11169
rect 5074 11160 5080 11172
rect 5132 11160 5138 11212
rect 4246 11092 4252 11144
rect 4304 11132 4310 11144
rect 4525 11135 4583 11141
rect 4525 11132 4537 11135
rect 4304 11104 4537 11132
rect 4304 11092 4310 11104
rect 4525 11101 4537 11104
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 3234 11024 3240 11076
rect 3292 11064 3298 11076
rect 4632 11064 4660 11095
rect 3292 11036 4660 11064
rect 3292 11024 3298 11036
rect 5074 11024 5080 11076
rect 5132 11064 5138 11076
rect 5350 11064 5356 11076
rect 5132 11036 5356 11064
rect 5132 11024 5138 11036
rect 5350 11024 5356 11036
rect 5408 11024 5414 11076
rect 5460 10996 5488 11308
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 8757 11339 8815 11345
rect 8757 11305 8769 11339
rect 8803 11305 8815 11339
rect 8757 11299 8815 11305
rect 9401 11339 9459 11345
rect 9401 11305 9413 11339
rect 9447 11336 9459 11339
rect 9490 11336 9496 11348
rect 9447 11308 9496 11336
rect 9447 11305 9459 11308
rect 9401 11299 9459 11305
rect 5988 11271 6046 11277
rect 5988 11237 6000 11271
rect 6034 11268 6046 11271
rect 8386 11268 8392 11280
rect 6034 11240 8392 11268
rect 6034 11237 6046 11240
rect 5988 11231 6046 11237
rect 8386 11228 8392 11240
rect 8444 11268 8450 11280
rect 8772 11268 8800 11299
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 9766 11296 9772 11348
rect 9824 11336 9830 11348
rect 9861 11339 9919 11345
rect 9861 11336 9873 11339
rect 9824 11308 9873 11336
rect 9824 11296 9830 11308
rect 9861 11305 9873 11308
rect 9907 11305 9919 11339
rect 12618 11336 12624 11348
rect 9861 11299 9919 11305
rect 10428 11308 12624 11336
rect 9306 11268 9312 11280
rect 8444 11240 9312 11268
rect 8444 11228 8450 11240
rect 9306 11228 9312 11240
rect 9364 11228 9370 11280
rect 10428 11277 10456 11308
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 12802 11296 12808 11348
rect 12860 11336 12866 11348
rect 13170 11336 13176 11348
rect 12860 11308 13176 11336
rect 12860 11296 12866 11308
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 13538 11296 13544 11348
rect 13596 11336 13602 11348
rect 15654 11336 15660 11348
rect 13596 11308 14872 11336
rect 15615 11308 15660 11336
rect 13596 11296 13602 11308
rect 10413 11271 10471 11277
rect 10413 11237 10425 11271
rect 10459 11237 10471 11271
rect 10413 11231 10471 11237
rect 12161 11271 12219 11277
rect 12161 11237 12173 11271
rect 12207 11268 12219 11271
rect 14090 11268 14096 11280
rect 12207 11240 14096 11268
rect 12207 11237 12219 11240
rect 12161 11231 12219 11237
rect 5718 11200 5724 11212
rect 5679 11172 5724 11200
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 6362 11200 6368 11212
rect 5828 11172 6368 11200
rect 5534 11092 5540 11144
rect 5592 11132 5598 11144
rect 5828 11132 5856 11172
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 7282 11160 7288 11212
rect 7340 11200 7346 11212
rect 7377 11203 7435 11209
rect 7377 11200 7389 11203
rect 7340 11172 7389 11200
rect 7340 11160 7346 11172
rect 7377 11169 7389 11172
rect 7423 11169 7435 11203
rect 7633 11203 7691 11209
rect 7633 11200 7645 11203
rect 7377 11163 7435 11169
rect 7484 11172 7645 11200
rect 7484 11132 7512 11172
rect 7633 11169 7645 11172
rect 7679 11169 7691 11203
rect 7633 11163 7691 11169
rect 8478 11160 8484 11212
rect 8536 11200 8542 11212
rect 9217 11203 9275 11209
rect 9217 11200 9229 11203
rect 8536 11172 9229 11200
rect 8536 11160 8542 11172
rect 9217 11169 9229 11172
rect 9263 11169 9275 11203
rect 9217 11163 9275 11169
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11200 9735 11203
rect 11790 11200 11796 11212
rect 9723 11172 11796 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 11790 11160 11796 11172
rect 11848 11200 11854 11212
rect 12066 11200 12072 11212
rect 11848 11172 12072 11200
rect 11848 11160 11854 11172
rect 12066 11160 12072 11172
rect 12124 11160 12130 11212
rect 5592 11104 5856 11132
rect 7392 11104 7512 11132
rect 5592 11092 5598 11104
rect 7392 11076 7420 11104
rect 8386 11092 8392 11144
rect 8444 11132 8450 11144
rect 11146 11132 11152 11144
rect 8444 11104 11152 11132
rect 8444 11092 8450 11104
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 7098 11064 7104 11076
rect 7059 11036 7104 11064
rect 7098 11024 7104 11036
rect 7156 11024 7162 11076
rect 7374 11024 7380 11076
rect 7432 11024 7438 11076
rect 12176 11064 12204 11231
rect 14090 11228 14096 11240
rect 14148 11228 14154 11280
rect 14461 11271 14519 11277
rect 14461 11237 14473 11271
rect 14507 11268 14519 11271
rect 14734 11268 14740 11280
rect 14507 11240 14740 11268
rect 14507 11237 14519 11240
rect 14461 11231 14519 11237
rect 14734 11228 14740 11240
rect 14792 11228 14798 11280
rect 14844 11268 14872 11308
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 16577 11339 16635 11345
rect 16577 11305 16589 11339
rect 16623 11336 16635 11339
rect 17957 11339 18015 11345
rect 17957 11336 17969 11339
rect 16623 11308 17969 11336
rect 16623 11305 16635 11308
rect 16577 11299 16635 11305
rect 17957 11305 17969 11308
rect 18003 11305 18015 11339
rect 17957 11299 18015 11305
rect 18506 11296 18512 11348
rect 18564 11336 18570 11348
rect 18785 11339 18843 11345
rect 18785 11336 18797 11339
rect 18564 11308 18797 11336
rect 18564 11296 18570 11308
rect 18785 11305 18797 11308
rect 18831 11305 18843 11339
rect 18785 11299 18843 11305
rect 18966 11296 18972 11348
rect 19024 11336 19030 11348
rect 19061 11339 19119 11345
rect 19061 11336 19073 11339
rect 19024 11308 19073 11336
rect 19024 11296 19030 11308
rect 19061 11305 19073 11308
rect 19107 11305 19119 11339
rect 20530 11336 20536 11348
rect 20491 11308 20536 11336
rect 19061 11299 19119 11305
rect 20530 11296 20536 11308
rect 20588 11296 20594 11348
rect 15749 11271 15807 11277
rect 15749 11268 15761 11271
rect 14844 11240 15761 11268
rect 15749 11237 15761 11240
rect 15795 11237 15807 11271
rect 15749 11231 15807 11237
rect 15838 11228 15844 11280
rect 15896 11268 15902 11280
rect 15896 11240 17080 11268
rect 15896 11228 15902 11240
rect 12434 11200 12440 11212
rect 12395 11172 12440 11200
rect 12434 11160 12440 11172
rect 12492 11160 12498 11212
rect 12704 11203 12762 11209
rect 12704 11169 12716 11203
rect 12750 11200 12762 11203
rect 12750 11172 13492 11200
rect 12750 11169 12762 11172
rect 12704 11163 12762 11169
rect 13464 11132 13492 11172
rect 13630 11160 13636 11212
rect 13688 11200 13694 11212
rect 14366 11200 14372 11212
rect 13688 11172 14372 11200
rect 13688 11160 13694 11172
rect 14366 11160 14372 11172
rect 14424 11160 14430 11212
rect 14553 11203 14611 11209
rect 14553 11169 14565 11203
rect 14599 11200 14611 11203
rect 16945 11203 17003 11209
rect 16945 11200 16957 11203
rect 14599 11172 15056 11200
rect 14599 11169 14611 11172
rect 14553 11163 14611 11169
rect 13906 11132 13912 11144
rect 13464 11104 13912 11132
rect 13906 11092 13912 11104
rect 13964 11092 13970 11144
rect 13998 11092 14004 11144
rect 14056 11132 14062 11144
rect 14645 11135 14703 11141
rect 14645 11132 14657 11135
rect 14056 11104 14657 11132
rect 14056 11092 14062 11104
rect 14645 11101 14657 11104
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 8772 11036 12204 11064
rect 1412 10968 5488 10996
rect 7742 10956 7748 11008
rect 7800 10996 7806 11008
rect 8772 10996 8800 11036
rect 13630 11024 13636 11076
rect 13688 11064 13694 11076
rect 13817 11067 13875 11073
rect 13817 11064 13829 11067
rect 13688 11036 13829 11064
rect 13688 11024 13694 11036
rect 13817 11033 13829 11036
rect 13863 11033 13875 11067
rect 14090 11064 14096 11076
rect 14051 11036 14096 11064
rect 13817 11027 13875 11033
rect 14090 11024 14096 11036
rect 14148 11024 14154 11076
rect 15028 11064 15056 11172
rect 15672 11172 16957 11200
rect 15470 11092 15476 11144
rect 15528 11132 15534 11144
rect 15672 11132 15700 11172
rect 16945 11169 16957 11172
rect 16991 11169 17003 11203
rect 17052 11200 17080 11240
rect 17126 11228 17132 11280
rect 17184 11268 17190 11280
rect 18049 11271 18107 11277
rect 18049 11268 18061 11271
rect 17184 11240 18061 11268
rect 17184 11228 17190 11240
rect 18049 11237 18061 11240
rect 18095 11237 18107 11271
rect 18049 11231 18107 11237
rect 18138 11228 18144 11280
rect 18196 11268 18202 11280
rect 19702 11268 19708 11280
rect 18196 11240 19708 11268
rect 18196 11228 18202 11240
rect 19702 11228 19708 11240
rect 19760 11228 19766 11280
rect 17402 11200 17408 11212
rect 17052 11172 17408 11200
rect 16945 11163 17003 11169
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 17586 11160 17592 11212
rect 17644 11200 17650 11212
rect 18601 11203 18659 11209
rect 18601 11200 18613 11203
rect 17644 11172 18613 11200
rect 17644 11160 17650 11172
rect 18601 11169 18613 11172
rect 18647 11169 18659 11203
rect 18601 11163 18659 11169
rect 18966 11160 18972 11212
rect 19024 11200 19030 11212
rect 19153 11203 19211 11209
rect 19153 11200 19165 11203
rect 19024 11172 19165 11200
rect 19024 11160 19030 11172
rect 19153 11169 19165 11172
rect 19199 11169 19211 11203
rect 19153 11163 19211 11169
rect 19420 11203 19478 11209
rect 19420 11169 19432 11203
rect 19466 11200 19478 11203
rect 20622 11200 20628 11212
rect 19466 11172 20628 11200
rect 19466 11169 19478 11172
rect 19420 11163 19478 11169
rect 20622 11160 20628 11172
rect 20680 11160 20686 11212
rect 15838 11132 15844 11144
rect 15528 11104 15700 11132
rect 15799 11104 15844 11132
rect 15528 11092 15534 11104
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 17034 11132 17040 11144
rect 16995 11104 17040 11132
rect 17034 11092 17040 11104
rect 17092 11092 17098 11144
rect 17218 11132 17224 11144
rect 17179 11104 17224 11132
rect 17218 11092 17224 11104
rect 17276 11092 17282 11144
rect 17862 11132 17868 11144
rect 17512 11104 17868 11132
rect 17512 11064 17540 11104
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 18233 11135 18291 11141
rect 18233 11101 18245 11135
rect 18279 11132 18291 11135
rect 19061 11135 19119 11141
rect 19061 11132 19073 11135
rect 18279 11104 19073 11132
rect 18279 11101 18291 11104
rect 18233 11095 18291 11101
rect 19061 11101 19073 11104
rect 19107 11101 19119 11135
rect 19061 11095 19119 11101
rect 20530 11092 20536 11144
rect 20588 11132 20594 11144
rect 21542 11132 21548 11144
rect 20588 11104 21548 11132
rect 20588 11092 20594 11104
rect 21542 11092 21548 11104
rect 21600 11092 21606 11144
rect 15028 11036 17540 11064
rect 17589 11067 17647 11073
rect 17589 11033 17601 11067
rect 17635 11064 17647 11067
rect 18414 11064 18420 11076
rect 17635 11036 18420 11064
rect 17635 11033 17647 11036
rect 17589 11027 17647 11033
rect 18414 11024 18420 11036
rect 18472 11024 18478 11076
rect 7800 10968 8800 10996
rect 7800 10956 7806 10968
rect 8846 10956 8852 11008
rect 8904 10996 8910 11008
rect 12802 10996 12808 11008
rect 8904 10968 12808 10996
rect 8904 10956 8910 10968
rect 12802 10956 12808 10968
rect 12860 10956 12866 11008
rect 14550 10956 14556 11008
rect 14608 10996 14614 11008
rect 15194 10996 15200 11008
rect 14608 10968 15200 10996
rect 14608 10956 14614 10968
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 15289 10999 15347 11005
rect 15289 10965 15301 10999
rect 15335 10996 15347 10999
rect 15930 10996 15936 11008
rect 15335 10968 15936 10996
rect 15335 10965 15347 10968
rect 15289 10959 15347 10965
rect 15930 10956 15936 10968
rect 15988 10956 15994 11008
rect 17126 10956 17132 11008
rect 17184 10996 17190 11008
rect 20438 10996 20444 11008
rect 17184 10968 20444 10996
rect 17184 10956 17190 10968
rect 20438 10956 20444 10968
rect 20496 10956 20502 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 3234 10792 3240 10804
rect 1872 10764 3096 10792
rect 3195 10764 3240 10792
rect 1872 10665 1900 10764
rect 3068 10724 3096 10764
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 3694 10792 3700 10804
rect 3655 10764 3700 10792
rect 3694 10752 3700 10764
rect 3752 10752 3758 10804
rect 3973 10795 4031 10801
rect 3973 10761 3985 10795
rect 4019 10792 4031 10795
rect 4154 10792 4160 10804
rect 4019 10764 4160 10792
rect 4019 10761 4031 10764
rect 3973 10755 4031 10761
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 4706 10752 4712 10804
rect 4764 10792 4770 10804
rect 6365 10795 6423 10801
rect 6365 10792 6377 10795
rect 4764 10764 6377 10792
rect 4764 10752 4770 10764
rect 6365 10761 6377 10764
rect 6411 10761 6423 10795
rect 6365 10755 6423 10761
rect 7466 10752 7472 10804
rect 7524 10792 7530 10804
rect 7561 10795 7619 10801
rect 7561 10792 7573 10795
rect 7524 10764 7573 10792
rect 7524 10752 7530 10764
rect 7561 10761 7573 10764
rect 7607 10792 7619 10795
rect 7653 10795 7711 10801
rect 7653 10792 7665 10795
rect 7607 10764 7665 10792
rect 7607 10761 7619 10764
rect 7561 10755 7619 10761
rect 7653 10761 7665 10764
rect 7699 10761 7711 10795
rect 7653 10755 7711 10761
rect 7760 10764 8524 10792
rect 4062 10724 4068 10736
rect 3068 10696 4068 10724
rect 4062 10684 4068 10696
rect 4120 10684 4126 10736
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10625 1915 10659
rect 4522 10656 4528 10668
rect 1857 10619 1915 10625
rect 3712 10628 4528 10656
rect 3510 10588 3516 10600
rect 3471 10560 3516 10588
rect 3510 10548 3516 10560
rect 3568 10548 3574 10600
rect 2124 10523 2182 10529
rect 2124 10489 2136 10523
rect 2170 10520 2182 10523
rect 2590 10520 2596 10532
rect 2170 10492 2596 10520
rect 2170 10489 2182 10492
rect 2124 10483 2182 10489
rect 2590 10480 2596 10492
rect 2648 10520 2654 10532
rect 3712 10520 3740 10628
rect 4522 10616 4528 10628
rect 4580 10616 4586 10668
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 5721 10659 5779 10665
rect 5721 10656 5733 10659
rect 5500 10628 5733 10656
rect 5500 10616 5506 10628
rect 5721 10625 5733 10628
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 7282 10616 7288 10668
rect 7340 10656 7346 10668
rect 7760 10656 7788 10764
rect 7837 10727 7895 10733
rect 7837 10693 7849 10727
rect 7883 10693 7895 10727
rect 7837 10687 7895 10693
rect 7340 10628 7788 10656
rect 7340 10616 7346 10628
rect 4890 10548 4896 10600
rect 4948 10588 4954 10600
rect 5077 10591 5135 10597
rect 5077 10588 5089 10591
rect 4948 10560 5089 10588
rect 4948 10548 4954 10560
rect 5077 10557 5089 10560
rect 5123 10588 5135 10591
rect 5537 10591 5595 10597
rect 5123 10560 5488 10588
rect 5123 10557 5135 10560
rect 5077 10551 5135 10557
rect 2648 10492 3740 10520
rect 4433 10523 4491 10529
rect 2648 10480 2654 10492
rect 4433 10489 4445 10523
rect 4479 10520 4491 10523
rect 5460 10520 5488 10560
rect 5537 10557 5549 10591
rect 5583 10588 5595 10591
rect 5626 10588 5632 10600
rect 5583 10560 5632 10588
rect 5583 10557 5595 10560
rect 5537 10551 5595 10557
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 6178 10588 6184 10600
rect 6139 10560 6184 10588
rect 6178 10548 6184 10560
rect 6236 10548 6242 10600
rect 6914 10548 6920 10600
rect 6972 10588 6978 10600
rect 7852 10588 7880 10687
rect 8496 10665 8524 10764
rect 8662 10752 8668 10804
rect 8720 10792 8726 10804
rect 8849 10795 8907 10801
rect 8849 10792 8861 10795
rect 8720 10764 8861 10792
rect 8720 10752 8726 10764
rect 8849 10761 8861 10764
rect 8895 10761 8907 10795
rect 8849 10755 8907 10761
rect 9306 10752 9312 10804
rect 9364 10792 9370 10804
rect 10410 10792 10416 10804
rect 9364 10764 9536 10792
rect 9364 10752 9370 10764
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10625 8539 10659
rect 8481 10619 8539 10625
rect 9030 10616 9036 10668
rect 9088 10656 9094 10668
rect 9508 10665 9536 10764
rect 9600 10764 10416 10792
rect 9309 10659 9367 10665
rect 9309 10656 9321 10659
rect 9088 10628 9321 10656
rect 9088 10616 9094 10628
rect 9309 10625 9321 10628
rect 9355 10625 9367 10659
rect 9309 10619 9367 10625
rect 9493 10659 9551 10665
rect 9493 10625 9505 10659
rect 9539 10625 9551 10659
rect 9493 10619 9551 10625
rect 6972 10560 7880 10588
rect 6972 10548 6978 10560
rect 8846 10548 8852 10600
rect 8904 10588 8910 10600
rect 9600 10588 9628 10764
rect 10410 10752 10416 10764
rect 10468 10752 10474 10804
rect 10686 10752 10692 10804
rect 10744 10752 10750 10804
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 11149 10795 11207 10801
rect 11149 10792 11161 10795
rect 11112 10764 11161 10792
rect 11112 10752 11118 10764
rect 11149 10761 11161 10764
rect 11195 10761 11207 10795
rect 11149 10755 11207 10761
rect 11701 10795 11759 10801
rect 11701 10761 11713 10795
rect 11747 10792 11759 10795
rect 12069 10795 12127 10801
rect 11747 10764 12020 10792
rect 11747 10761 11759 10764
rect 11701 10755 11759 10761
rect 10704 10724 10732 10752
rect 11992 10724 12020 10764
rect 12069 10761 12081 10795
rect 12115 10792 12127 10795
rect 13446 10792 13452 10804
rect 12115 10764 13452 10792
rect 12115 10761 12127 10764
rect 12069 10755 12127 10761
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 14182 10792 14188 10804
rect 13832 10764 14188 10792
rect 12434 10724 12440 10736
rect 10704 10696 11928 10724
rect 11992 10696 12440 10724
rect 9766 10588 9772 10600
rect 8904 10560 9628 10588
rect 9727 10560 9772 10588
rect 8904 10548 8910 10560
rect 9766 10548 9772 10560
rect 9824 10548 9830 10600
rect 11900 10597 11928 10696
rect 12434 10684 12440 10696
rect 12492 10684 12498 10736
rect 13832 10724 13860 10764
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 14829 10795 14887 10801
rect 14829 10761 14841 10795
rect 14875 10792 14887 10795
rect 16945 10795 17003 10801
rect 14875 10764 16427 10792
rect 14875 10761 14887 10764
rect 14829 10755 14887 10761
rect 16399 10724 16427 10764
rect 16945 10761 16957 10795
rect 16991 10792 17003 10795
rect 17310 10792 17316 10804
rect 16991 10764 17316 10792
rect 16991 10761 17003 10764
rect 16945 10755 17003 10761
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 18064 10764 19012 10792
rect 18064 10724 18092 10764
rect 13096 10696 13860 10724
rect 13924 10696 15599 10724
rect 16399 10696 18092 10724
rect 18984 10724 19012 10764
rect 19058 10752 19064 10804
rect 19116 10792 19122 10804
rect 19705 10795 19763 10801
rect 19705 10792 19717 10795
rect 19116 10764 19717 10792
rect 19116 10752 19122 10764
rect 19705 10761 19717 10764
rect 19751 10761 19763 10795
rect 19705 10755 19763 10761
rect 19426 10724 19432 10736
rect 18984 10696 19432 10724
rect 13096 10665 13124 10696
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10625 13139 10659
rect 13081 10619 13139 10625
rect 13630 10616 13636 10668
rect 13688 10656 13694 10668
rect 13924 10656 13952 10696
rect 13688 10628 13952 10656
rect 13688 10616 13694 10628
rect 13998 10616 14004 10668
rect 14056 10656 14062 10668
rect 14056 10628 14101 10656
rect 14056 10616 14062 10628
rect 15194 10616 15200 10668
rect 15252 10656 15258 10668
rect 15289 10659 15347 10665
rect 15289 10656 15301 10659
rect 15252 10628 15301 10656
rect 15252 10616 15258 10628
rect 15289 10625 15301 10628
rect 15335 10625 15347 10659
rect 15289 10619 15347 10625
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10625 15531 10659
rect 15571 10656 15599 10696
rect 19426 10684 19432 10696
rect 19484 10684 19490 10736
rect 16393 10659 16451 10665
rect 16393 10656 16405 10659
rect 15571 10628 16405 10656
rect 15473 10619 15531 10625
rect 16393 10625 16405 10628
rect 16439 10656 16451 10659
rect 17126 10656 17132 10668
rect 16439 10628 17132 10656
rect 16439 10625 16451 10628
rect 16393 10619 16451 10625
rect 11517 10591 11575 10597
rect 9968 10560 11284 10588
rect 6086 10520 6092 10532
rect 4479 10492 5212 10520
rect 5460 10492 6092 10520
rect 4479 10489 4491 10492
rect 4433 10483 4491 10489
rect 1397 10455 1455 10461
rect 1397 10421 1409 10455
rect 1443 10452 1455 10455
rect 2222 10452 2228 10464
rect 1443 10424 2228 10452
rect 1443 10421 1455 10424
rect 1397 10415 1455 10421
rect 2222 10412 2228 10424
rect 2280 10412 2286 10464
rect 4341 10455 4399 10461
rect 4341 10421 4353 10455
rect 4387 10452 4399 10455
rect 4706 10452 4712 10464
rect 4387 10424 4712 10452
rect 4387 10421 4399 10424
rect 4341 10415 4399 10421
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 5184 10461 5212 10492
rect 5644 10461 5672 10492
rect 6086 10480 6092 10492
rect 6144 10480 6150 10532
rect 9968 10520 9996 10560
rect 7484 10492 9996 10520
rect 10036 10523 10094 10529
rect 5169 10455 5227 10461
rect 5169 10421 5181 10455
rect 5215 10421 5227 10455
rect 5169 10415 5227 10421
rect 5629 10455 5687 10461
rect 5629 10421 5641 10455
rect 5675 10421 5687 10455
rect 5629 10415 5687 10421
rect 5902 10412 5908 10464
rect 5960 10452 5966 10464
rect 7484 10452 7512 10492
rect 10036 10489 10048 10523
rect 10082 10520 10094 10523
rect 10134 10520 10140 10532
rect 10082 10492 10140 10520
rect 10082 10489 10094 10492
rect 10036 10483 10094 10489
rect 10134 10480 10140 10492
rect 10192 10480 10198 10532
rect 5960 10424 7512 10452
rect 7561 10455 7619 10461
rect 5960 10412 5966 10424
rect 7561 10421 7573 10455
rect 7607 10452 7619 10455
rect 8205 10455 8263 10461
rect 8205 10452 8217 10455
rect 7607 10424 8217 10452
rect 7607 10421 7619 10424
rect 7561 10415 7619 10421
rect 8205 10421 8217 10424
rect 8251 10421 8263 10455
rect 8205 10415 8263 10421
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 9217 10455 9275 10461
rect 8352 10424 8397 10452
rect 8352 10412 8358 10424
rect 9217 10421 9229 10455
rect 9263 10452 9275 10455
rect 10686 10452 10692 10464
rect 9263 10424 10692 10452
rect 9263 10421 9275 10424
rect 9217 10415 9275 10421
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 11256 10452 11284 10560
rect 11517 10557 11529 10591
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 11885 10591 11943 10597
rect 11885 10557 11897 10591
rect 11931 10588 11943 10591
rect 13446 10588 13452 10600
rect 11931 10560 13452 10588
rect 11931 10557 11943 10560
rect 11885 10551 11943 10557
rect 11330 10480 11336 10532
rect 11388 10520 11394 10532
rect 11532 10520 11560 10551
rect 13446 10548 13452 10560
rect 13504 10588 13510 10600
rect 13814 10588 13820 10600
rect 13504 10560 13820 10588
rect 13504 10548 13510 10560
rect 13814 10548 13820 10560
rect 13872 10548 13878 10600
rect 15378 10588 15384 10600
rect 14752 10560 15384 10588
rect 12066 10520 12072 10532
rect 11388 10492 12072 10520
rect 11388 10480 11394 10492
rect 12066 10480 12072 10492
rect 12124 10480 12130 10532
rect 14752 10520 14780 10560
rect 15378 10548 15384 10560
rect 15436 10548 15442 10600
rect 15488 10588 15516 10619
rect 17126 10616 17132 10628
rect 17184 10616 17190 10668
rect 17494 10656 17500 10668
rect 17455 10628 17500 10656
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 15838 10588 15844 10600
rect 15488 10560 15844 10588
rect 15838 10548 15844 10560
rect 15896 10588 15902 10600
rect 18049 10591 18107 10597
rect 15896 10560 17540 10588
rect 15896 10548 15902 10560
rect 17144 10532 17172 10560
rect 12452 10492 14780 10520
rect 12158 10452 12164 10464
rect 11256 10424 12164 10452
rect 12158 10412 12164 10424
rect 12216 10412 12222 10464
rect 12452 10461 12480 10492
rect 14826 10480 14832 10532
rect 14884 10520 14890 10532
rect 16298 10520 16304 10532
rect 14884 10492 15884 10520
rect 16259 10492 16304 10520
rect 14884 10480 14890 10492
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10421 12495 10455
rect 12802 10452 12808 10464
rect 12763 10424 12808 10452
rect 12437 10415 12495 10421
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 13449 10455 13507 10461
rect 13449 10452 13461 10455
rect 12943 10424 13461 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 13449 10421 13461 10424
rect 13495 10421 13507 10455
rect 13814 10452 13820 10464
rect 13775 10424 13820 10452
rect 13449 10415 13507 10421
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 13909 10455 13967 10461
rect 13909 10421 13921 10455
rect 13955 10452 13967 10455
rect 14366 10452 14372 10464
rect 13955 10424 14372 10452
rect 13955 10421 13967 10424
rect 13909 10415 13967 10421
rect 14366 10412 14372 10424
rect 14424 10452 14430 10464
rect 15102 10452 15108 10464
rect 14424 10424 15108 10452
rect 14424 10412 14430 10424
rect 15102 10412 15108 10424
rect 15160 10412 15166 10464
rect 15197 10455 15255 10461
rect 15197 10421 15209 10455
rect 15243 10452 15255 10455
rect 15654 10452 15660 10464
rect 15243 10424 15660 10452
rect 15243 10421 15255 10424
rect 15197 10415 15255 10421
rect 15654 10412 15660 10424
rect 15712 10412 15718 10464
rect 15856 10461 15884 10492
rect 16298 10480 16304 10492
rect 16356 10480 16362 10532
rect 17126 10480 17132 10532
rect 17184 10480 17190 10532
rect 17310 10520 17316 10532
rect 17271 10492 17316 10520
rect 17310 10480 17316 10492
rect 17368 10480 17374 10532
rect 15841 10455 15899 10461
rect 15841 10421 15853 10455
rect 15887 10421 15899 10455
rect 16206 10452 16212 10464
rect 16167 10424 16212 10452
rect 15841 10415 15899 10421
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 16574 10412 16580 10464
rect 16632 10452 16638 10464
rect 17402 10452 17408 10464
rect 16632 10424 17408 10452
rect 16632 10412 16638 10424
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 17512 10452 17540 10560
rect 18049 10557 18061 10591
rect 18095 10588 18107 10591
rect 18138 10588 18144 10600
rect 18095 10560 18144 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 18316 10591 18374 10597
rect 18316 10557 18328 10591
rect 18362 10588 18374 10591
rect 19242 10588 19248 10600
rect 18362 10560 19248 10588
rect 18362 10557 18374 10560
rect 18316 10551 18374 10557
rect 19242 10548 19248 10560
rect 19300 10548 19306 10600
rect 19720 10588 19748 10755
rect 19886 10616 19892 10668
rect 19944 10656 19950 10668
rect 20533 10659 20591 10665
rect 19944 10628 20392 10656
rect 19944 10616 19950 10628
rect 20364 10597 20392 10628
rect 20533 10625 20545 10659
rect 20579 10625 20591 10659
rect 20533 10619 20591 10625
rect 20257 10591 20315 10597
rect 20257 10588 20269 10591
rect 19720 10560 20269 10588
rect 20257 10557 20269 10560
rect 20303 10557 20315 10591
rect 20257 10551 20315 10557
rect 20349 10591 20407 10597
rect 20349 10557 20361 10591
rect 20395 10557 20407 10591
rect 20349 10551 20407 10557
rect 20438 10548 20444 10600
rect 20496 10588 20502 10600
rect 20548 10588 20576 10619
rect 20496 10560 20576 10588
rect 20496 10548 20502 10560
rect 17862 10480 17868 10532
rect 17920 10520 17926 10532
rect 17920 10492 19932 10520
rect 17920 10480 17926 10492
rect 18874 10452 18880 10464
rect 17512 10424 18880 10452
rect 18874 10412 18880 10424
rect 18932 10452 18938 10464
rect 19904 10461 19932 10492
rect 19429 10455 19487 10461
rect 19429 10452 19441 10455
rect 18932 10424 19441 10452
rect 18932 10412 18938 10424
rect 19429 10421 19441 10424
rect 19475 10421 19487 10455
rect 19429 10415 19487 10421
rect 19889 10455 19947 10461
rect 19889 10421 19901 10455
rect 19935 10421 19947 10455
rect 19889 10415 19947 10421
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 1673 10251 1731 10257
rect 1673 10217 1685 10251
rect 1719 10248 1731 10251
rect 1762 10248 1768 10260
rect 1719 10220 1768 10248
rect 1719 10217 1731 10220
rect 1673 10211 1731 10217
rect 1762 10208 1768 10220
rect 1820 10208 1826 10260
rect 1854 10208 1860 10260
rect 1912 10248 1918 10260
rect 2038 10248 2044 10260
rect 1912 10220 2044 10248
rect 1912 10208 1918 10220
rect 2038 10208 2044 10220
rect 2096 10208 2102 10260
rect 2866 10208 2872 10260
rect 2924 10248 2930 10260
rect 3237 10251 3295 10257
rect 3237 10248 3249 10251
rect 2924 10220 3249 10248
rect 2924 10208 2930 10220
rect 3237 10217 3249 10220
rect 3283 10217 3295 10251
rect 3237 10211 3295 10217
rect 4522 10208 4528 10260
rect 4580 10248 4586 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 4580 10220 5457 10248
rect 4580 10208 4586 10220
rect 5445 10217 5457 10220
rect 5491 10217 5503 10251
rect 5445 10211 5503 10217
rect 5626 10208 5632 10260
rect 5684 10248 5690 10260
rect 6178 10248 6184 10260
rect 5684 10220 6184 10248
rect 5684 10208 5690 10220
rect 6178 10208 6184 10220
rect 6236 10208 6242 10260
rect 6638 10248 6644 10260
rect 6288 10220 6644 10248
rect 2409 10183 2467 10189
rect 2409 10149 2421 10183
rect 2455 10180 2467 10183
rect 2774 10180 2780 10192
rect 2455 10152 2780 10180
rect 2455 10149 2467 10152
rect 2409 10143 2467 10149
rect 2774 10140 2780 10152
rect 2832 10140 2838 10192
rect 6288 10180 6316 10220
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 7745 10251 7803 10257
rect 7745 10248 7757 10251
rect 7248 10220 7757 10248
rect 7248 10208 7254 10220
rect 7745 10217 7757 10220
rect 7791 10217 7803 10251
rect 8202 10248 8208 10260
rect 8163 10220 8208 10248
rect 7745 10211 7803 10217
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 8294 10208 8300 10260
rect 8352 10248 8358 10260
rect 9030 10248 9036 10260
rect 8352 10220 9036 10248
rect 8352 10208 8358 10220
rect 9030 10208 9036 10220
rect 9088 10248 9094 10260
rect 10502 10248 10508 10260
rect 9088 10220 10508 10248
rect 9088 10208 9094 10220
rect 10502 10208 10508 10220
rect 10560 10208 10566 10260
rect 10686 10248 10692 10260
rect 10647 10220 10692 10248
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 11054 10208 11060 10260
rect 11112 10248 11118 10260
rect 12618 10248 12624 10260
rect 11112 10220 12624 10248
rect 11112 10208 11118 10220
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 12805 10251 12863 10257
rect 12805 10217 12817 10251
rect 12851 10248 12863 10251
rect 14458 10248 14464 10260
rect 12851 10220 14464 10248
rect 12851 10217 12863 10220
rect 12805 10211 12863 10217
rect 14458 10208 14464 10220
rect 14516 10208 14522 10260
rect 14829 10251 14887 10257
rect 14829 10217 14841 10251
rect 14875 10248 14887 10251
rect 16114 10248 16120 10260
rect 14875 10220 16120 10248
rect 14875 10217 14887 10220
rect 14829 10211 14887 10217
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 16206 10208 16212 10260
rect 16264 10248 16270 10260
rect 16761 10251 16819 10257
rect 16761 10248 16773 10251
rect 16264 10220 16773 10248
rect 16264 10208 16270 10220
rect 16761 10217 16773 10220
rect 16807 10217 16819 10251
rect 16761 10211 16819 10217
rect 17034 10208 17040 10260
rect 17092 10248 17098 10260
rect 17405 10251 17463 10257
rect 17405 10248 17417 10251
rect 17092 10220 17417 10248
rect 17092 10208 17098 10220
rect 17405 10217 17417 10220
rect 17451 10217 17463 10251
rect 17405 10211 17463 10217
rect 17494 10208 17500 10260
rect 17552 10248 17558 10260
rect 17773 10251 17831 10257
rect 17773 10248 17785 10251
rect 17552 10220 17785 10248
rect 17552 10208 17558 10220
rect 17773 10217 17785 10220
rect 17819 10217 17831 10251
rect 17773 10211 17831 10217
rect 18230 10208 18236 10260
rect 18288 10248 18294 10260
rect 20162 10248 20168 10260
rect 18288 10220 20168 10248
rect 18288 10208 18294 10220
rect 20162 10208 20168 10220
rect 20220 10208 20226 10260
rect 20441 10251 20499 10257
rect 20441 10217 20453 10251
rect 20487 10248 20499 10251
rect 20622 10248 20628 10260
rect 20487 10220 20628 10248
rect 20487 10217 20499 10220
rect 20441 10211 20499 10217
rect 20622 10208 20628 10220
rect 20680 10208 20686 10260
rect 3068 10152 6316 10180
rect 6457 10183 6515 10189
rect 1489 10115 1547 10121
rect 1489 10081 1501 10115
rect 1535 10112 1547 10115
rect 2314 10112 2320 10124
rect 1535 10084 2320 10112
rect 1535 10081 1547 10084
rect 1489 10075 1547 10081
rect 2314 10072 2320 10084
rect 2372 10072 2378 10124
rect 2498 10112 2504 10124
rect 2459 10084 2504 10112
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 3068 10121 3096 10152
rect 6457 10149 6469 10183
rect 6503 10180 6515 10183
rect 12526 10180 12532 10192
rect 6503 10152 12532 10180
rect 6503 10149 6515 10152
rect 6457 10143 6515 10149
rect 12526 10140 12532 10152
rect 12584 10140 12590 10192
rect 12897 10183 12955 10189
rect 12897 10149 12909 10183
rect 12943 10180 12955 10183
rect 19328 10183 19386 10189
rect 12943 10152 14964 10180
rect 12943 10149 12955 10152
rect 12897 10143 12955 10149
rect 3053 10115 3111 10121
rect 3053 10081 3065 10115
rect 3099 10081 3111 10115
rect 4062 10112 4068 10124
rect 4023 10084 4068 10112
rect 3053 10075 3111 10081
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 4154 10072 4160 10124
rect 4212 10112 4218 10124
rect 4321 10115 4379 10121
rect 4321 10112 4333 10115
rect 4212 10084 4333 10112
rect 4212 10072 4218 10084
rect 4321 10081 4333 10084
rect 4367 10081 4379 10115
rect 4321 10075 4379 10081
rect 4706 10072 4712 10124
rect 4764 10112 4770 10124
rect 4890 10112 4896 10124
rect 4764 10084 4896 10112
rect 4764 10072 4770 10084
rect 4890 10072 4896 10084
rect 4948 10072 4954 10124
rect 6365 10115 6423 10121
rect 6365 10081 6377 10115
rect 6411 10112 6423 10115
rect 7006 10112 7012 10124
rect 6411 10084 7012 10112
rect 6411 10081 6423 10084
rect 6365 10075 6423 10081
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 7193 10115 7251 10121
rect 7193 10081 7205 10115
rect 7239 10081 7251 10115
rect 7193 10075 7251 10081
rect 7285 10115 7343 10121
rect 7285 10081 7297 10115
rect 7331 10112 7343 10115
rect 7331 10084 7696 10112
rect 7331 10081 7343 10084
rect 7285 10075 7343 10081
rect 2332 9976 2360 10072
rect 2590 10044 2596 10056
rect 2551 10016 2596 10044
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 6086 10004 6092 10056
rect 6144 10044 6150 10056
rect 6549 10047 6607 10053
rect 6549 10044 6561 10047
rect 6144 10016 6561 10044
rect 6144 10004 6150 10016
rect 6549 10013 6561 10016
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 6638 10004 6644 10056
rect 6696 10044 6702 10056
rect 7208 10044 7236 10075
rect 6696 10016 7236 10044
rect 7377 10047 7435 10053
rect 6696 10004 6702 10016
rect 7377 10013 7389 10047
rect 7423 10013 7435 10047
rect 7668 10044 7696 10084
rect 7742 10072 7748 10124
rect 7800 10112 7806 10124
rect 7929 10115 7987 10121
rect 7929 10112 7941 10115
rect 7800 10084 7941 10112
rect 7800 10072 7806 10084
rect 7929 10081 7941 10084
rect 7975 10081 7987 10115
rect 7929 10075 7987 10081
rect 8018 10072 8024 10124
rect 8076 10112 8082 10124
rect 8076 10084 8121 10112
rect 8076 10072 8082 10084
rect 8294 10072 8300 10124
rect 8352 10112 8358 10124
rect 8662 10112 8668 10124
rect 8352 10084 8668 10112
rect 8352 10072 8358 10084
rect 8662 10072 8668 10084
rect 8720 10112 8726 10124
rect 8941 10115 8999 10121
rect 8941 10112 8953 10115
rect 8720 10084 8953 10112
rect 8720 10072 8726 10084
rect 8941 10081 8953 10084
rect 8987 10081 8999 10115
rect 8941 10075 8999 10081
rect 9493 10115 9551 10121
rect 9493 10081 9505 10115
rect 9539 10112 9551 10115
rect 9858 10112 9864 10124
rect 9539 10084 9864 10112
rect 9539 10081 9551 10084
rect 9493 10075 9551 10081
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 10045 10115 10103 10121
rect 10045 10081 10057 10115
rect 10091 10112 10103 10115
rect 10091 10084 10463 10112
rect 10091 10081 10103 10084
rect 10045 10075 10103 10081
rect 8754 10044 8760 10056
rect 7668 10016 8760 10044
rect 7377 10007 7435 10013
rect 3878 9976 3884 9988
rect 2332 9948 3884 9976
rect 3878 9936 3884 9948
rect 3936 9936 3942 9988
rect 5000 9948 6960 9976
rect 2041 9911 2099 9917
rect 2041 9877 2053 9911
rect 2087 9908 2099 9911
rect 2314 9908 2320 9920
rect 2087 9880 2320 9908
rect 2087 9877 2099 9880
rect 2041 9871 2099 9877
rect 2314 9868 2320 9880
rect 2372 9868 2378 9920
rect 3510 9868 3516 9920
rect 3568 9908 3574 9920
rect 5000 9908 5028 9948
rect 5994 9908 6000 9920
rect 3568 9880 5028 9908
rect 5955 9880 6000 9908
rect 3568 9868 3574 9880
rect 5994 9868 6000 9880
rect 6052 9868 6058 9920
rect 6822 9908 6828 9920
rect 6783 9880 6828 9908
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 6932 9908 6960 9948
rect 7282 9936 7288 9988
rect 7340 9976 7346 9988
rect 7392 9976 7420 10007
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 8846 10004 8852 10056
rect 8904 10044 8910 10056
rect 9030 10044 9036 10056
rect 8904 10016 9036 10044
rect 8904 10004 8910 10016
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 9122 10004 9128 10056
rect 9180 10044 9186 10056
rect 9950 10044 9956 10056
rect 9180 10016 9225 10044
rect 9784 10016 9956 10044
rect 9180 10004 9186 10016
rect 7340 9948 7420 9976
rect 7340 9936 7346 9948
rect 7466 9936 7472 9988
rect 7524 9976 7530 9988
rect 7834 9976 7840 9988
rect 7524 9948 7840 9976
rect 7524 9936 7530 9948
rect 7834 9936 7840 9948
rect 7892 9936 7898 9988
rect 8110 9936 8116 9988
rect 8168 9976 8174 9988
rect 8386 9976 8392 9988
rect 8168 9948 8392 9976
rect 8168 9936 8174 9948
rect 8386 9936 8392 9948
rect 8444 9936 8450 9988
rect 8573 9979 8631 9985
rect 8573 9945 8585 9979
rect 8619 9976 8631 9979
rect 9784 9976 9812 10016
rect 9950 10004 9956 10016
rect 10008 10004 10014 10056
rect 10137 10047 10195 10053
rect 10137 10013 10149 10047
rect 10183 10013 10195 10047
rect 10318 10044 10324 10056
rect 10279 10016 10324 10044
rect 10137 10007 10195 10013
rect 8619 9948 9812 9976
rect 10152 9976 10180 10007
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 10435 10044 10463 10084
rect 10502 10072 10508 10124
rect 10560 10112 10566 10124
rect 11054 10112 11060 10124
rect 10560 10084 10723 10112
rect 11015 10084 11060 10112
rect 10560 10072 10566 10084
rect 10594 10044 10600 10056
rect 10435 10016 10600 10044
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 10695 10044 10723 10084
rect 11054 10072 11060 10084
rect 11112 10072 11118 10124
rect 11790 10072 11796 10124
rect 11848 10112 11854 10124
rect 11885 10115 11943 10121
rect 11885 10112 11897 10115
rect 11848 10084 11897 10112
rect 11848 10072 11854 10084
rect 11885 10081 11897 10084
rect 11931 10081 11943 10115
rect 11885 10075 11943 10081
rect 13446 10072 13452 10124
rect 13504 10112 13510 10124
rect 13817 10115 13875 10121
rect 13817 10112 13829 10115
rect 13504 10084 13829 10112
rect 13504 10072 13510 10084
rect 13817 10081 13829 10084
rect 13863 10081 13875 10115
rect 13817 10075 13875 10081
rect 14550 10072 14556 10124
rect 14608 10112 14614 10124
rect 14645 10115 14703 10121
rect 14645 10112 14657 10115
rect 14608 10084 14657 10112
rect 14608 10072 14614 10084
rect 14645 10081 14657 10084
rect 14691 10081 14703 10115
rect 14936 10112 14964 10152
rect 15396 10152 19196 10180
rect 15396 10112 15424 10152
rect 14936 10084 15424 10112
rect 15556 10115 15614 10121
rect 14645 10075 14703 10081
rect 15556 10081 15568 10115
rect 15602 10112 15614 10115
rect 17126 10112 17132 10124
rect 15602 10084 17132 10112
rect 15602 10081 15614 10084
rect 15556 10075 15614 10081
rect 17126 10072 17132 10084
rect 17184 10072 17190 10124
rect 17865 10115 17923 10121
rect 17865 10081 17877 10115
rect 17911 10112 17923 10115
rect 18230 10112 18236 10124
rect 17911 10084 18236 10112
rect 17911 10081 17923 10084
rect 17865 10075 17923 10081
rect 18230 10072 18236 10084
rect 18288 10072 18294 10124
rect 18414 10072 18420 10124
rect 18472 10112 18478 10124
rect 18509 10115 18567 10121
rect 18509 10112 18521 10115
rect 18472 10084 18521 10112
rect 18472 10072 18478 10084
rect 18509 10081 18521 10084
rect 18555 10081 18567 10115
rect 19058 10112 19064 10124
rect 19019 10084 19064 10112
rect 18509 10075 18567 10081
rect 19058 10072 19064 10084
rect 19116 10072 19122 10124
rect 19168 10112 19196 10152
rect 19328 10149 19340 10183
rect 19374 10180 19386 10183
rect 19610 10180 19616 10192
rect 19374 10152 19616 10180
rect 19374 10149 19386 10152
rect 19328 10143 19386 10149
rect 19610 10140 19616 10152
rect 19668 10140 19674 10192
rect 19886 10112 19892 10124
rect 19168 10084 19892 10112
rect 19886 10072 19892 10084
rect 19944 10072 19950 10124
rect 11149 10047 11207 10053
rect 10695 10016 11100 10044
rect 11072 9988 11100 10016
rect 11149 10013 11161 10047
rect 11195 10013 11207 10047
rect 11149 10007 11207 10013
rect 11333 10047 11391 10053
rect 11333 10013 11345 10047
rect 11379 10044 11391 10047
rect 11698 10044 11704 10056
rect 11379 10016 11704 10044
rect 11379 10013 11391 10016
rect 11333 10007 11391 10013
rect 10502 9976 10508 9988
rect 10152 9948 10508 9976
rect 8619 9945 8631 9948
rect 8573 9939 8631 9945
rect 10502 9936 10508 9948
rect 10560 9936 10566 9988
rect 11054 9936 11060 9988
rect 11112 9936 11118 9988
rect 9493 9911 9551 9917
rect 9493 9908 9505 9911
rect 6932 9880 9505 9908
rect 9493 9877 9505 9880
rect 9539 9877 9551 9911
rect 9674 9908 9680 9920
rect 9635 9880 9680 9908
rect 9493 9871 9551 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 9858 9868 9864 9920
rect 9916 9908 9922 9920
rect 11164 9908 11192 10007
rect 11698 10004 11704 10016
rect 11756 10004 11762 10056
rect 12986 10044 12992 10056
rect 12947 10016 12992 10044
rect 12986 10004 12992 10016
rect 13044 10004 13050 10056
rect 13909 10047 13967 10053
rect 13909 10013 13921 10047
rect 13955 10013 13967 10047
rect 13909 10007 13967 10013
rect 14093 10047 14151 10053
rect 14093 10013 14105 10047
rect 14139 10044 14151 10047
rect 14182 10044 14188 10056
rect 14139 10016 14188 10044
rect 14139 10013 14151 10016
rect 14093 10007 14151 10013
rect 11606 9936 11612 9988
rect 11664 9976 11670 9988
rect 12158 9976 12164 9988
rect 11664 9948 12164 9976
rect 11664 9936 11670 9948
rect 12158 9936 12164 9948
rect 12216 9936 12222 9988
rect 12066 9908 12072 9920
rect 9916 9880 11192 9908
rect 12027 9880 12072 9908
rect 9916 9868 9922 9880
rect 12066 9868 12072 9880
rect 12124 9868 12130 9920
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 13446 9908 13452 9920
rect 12492 9880 12537 9908
rect 13407 9880 13452 9908
rect 12492 9868 12498 9880
rect 13446 9868 13452 9880
rect 13504 9868 13510 9920
rect 13538 9868 13544 9920
rect 13596 9908 13602 9920
rect 13924 9908 13952 10007
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 14918 10004 14924 10056
rect 14976 10044 14982 10056
rect 15289 10047 15347 10053
rect 15289 10044 15301 10047
rect 14976 10016 15301 10044
rect 14976 10004 14982 10016
rect 15289 10013 15301 10016
rect 15335 10013 15347 10047
rect 17218 10044 17224 10056
rect 17179 10016 17224 10044
rect 15289 10007 15347 10013
rect 17218 10004 17224 10016
rect 17276 10044 17282 10056
rect 17494 10044 17500 10056
rect 17276 10016 17500 10044
rect 17276 10004 17282 10016
rect 17494 10004 17500 10016
rect 17552 10004 17558 10056
rect 17586 10004 17592 10056
rect 17644 10044 17650 10056
rect 17957 10047 18015 10053
rect 17957 10044 17969 10047
rect 17644 10016 17969 10044
rect 17644 10004 17650 10016
rect 17957 10013 17969 10016
rect 18003 10013 18015 10047
rect 17957 10007 18015 10013
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 19076 10044 19104 10072
rect 18380 10016 19104 10044
rect 18380 10004 18386 10016
rect 18693 9979 18751 9985
rect 16224 9948 18644 9976
rect 13596 9880 13952 9908
rect 13596 9868 13602 9880
rect 14458 9868 14464 9920
rect 14516 9908 14522 9920
rect 16224 9908 16252 9948
rect 14516 9880 16252 9908
rect 16669 9911 16727 9917
rect 14516 9868 14522 9880
rect 16669 9877 16681 9911
rect 16715 9908 16727 9911
rect 17034 9908 17040 9920
rect 16715 9880 17040 9908
rect 16715 9877 16727 9880
rect 16669 9871 16727 9877
rect 17034 9868 17040 9880
rect 17092 9868 17098 9920
rect 18616 9908 18644 9948
rect 18693 9945 18705 9979
rect 18739 9976 18751 9979
rect 18782 9976 18788 9988
rect 18739 9948 18788 9976
rect 18739 9945 18751 9948
rect 18693 9939 18751 9945
rect 18782 9936 18788 9948
rect 18840 9936 18846 9988
rect 19058 9908 19064 9920
rect 18616 9880 19064 9908
rect 19058 9868 19064 9880
rect 19116 9868 19122 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 2498 9664 2504 9716
rect 2556 9704 2562 9716
rect 3145 9707 3203 9713
rect 3145 9704 3157 9707
rect 2556 9676 3157 9704
rect 2556 9664 2562 9676
rect 3145 9673 3157 9676
rect 3191 9673 3203 9707
rect 3145 9667 3203 9673
rect 3878 9664 3884 9716
rect 3936 9704 3942 9716
rect 8662 9704 8668 9716
rect 3936 9676 8668 9704
rect 3936 9664 3942 9676
rect 1765 9639 1823 9645
rect 1765 9605 1777 9639
rect 1811 9636 1823 9639
rect 4065 9639 4123 9645
rect 1811 9608 3188 9636
rect 1811 9605 1823 9608
rect 1765 9599 1823 9605
rect 3160 9580 3188 9608
rect 4065 9605 4077 9639
rect 4111 9636 4123 9639
rect 4246 9636 4252 9648
rect 4111 9608 4252 9636
rect 4111 9605 4123 9608
rect 4065 9599 4123 9605
rect 4246 9596 4252 9608
rect 4304 9596 4310 9648
rect 5721 9639 5779 9645
rect 5721 9636 5733 9639
rect 4816 9608 5733 9636
rect 2590 9528 2596 9580
rect 2648 9568 2654 9580
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 2648 9540 2697 9568
rect 2648 9528 2654 9540
rect 2685 9537 2697 9540
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9500 1639 9503
rect 1762 9500 1768 9512
rect 1627 9472 1768 9500
rect 1627 9469 1639 9472
rect 1581 9463 1639 9469
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 2406 9432 2412 9444
rect 2148 9404 2412 9432
rect 2148 9373 2176 9404
rect 2406 9392 2412 9404
rect 2464 9392 2470 9444
rect 2700 9432 2728 9531
rect 3142 9528 3148 9580
rect 3200 9528 3206 9580
rect 3326 9528 3332 9580
rect 3384 9568 3390 9580
rect 3602 9568 3608 9580
rect 3384 9540 3608 9568
rect 3384 9528 3390 9540
rect 3602 9528 3608 9540
rect 3660 9528 3666 9580
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9568 3847 9571
rect 4154 9568 4160 9580
rect 3835 9540 4160 9568
rect 3835 9537 3847 9540
rect 3789 9531 3847 9537
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 4617 9571 4675 9577
rect 4617 9568 4629 9571
rect 4336 9540 4629 9568
rect 3510 9500 3516 9512
rect 3471 9472 3516 9500
rect 3510 9460 3516 9472
rect 3568 9460 3574 9512
rect 4336 9432 4364 9540
rect 4617 9537 4629 9540
rect 4663 9537 4675 9571
rect 4617 9531 4675 9537
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9500 4491 9503
rect 4816 9500 4844 9608
rect 5721 9605 5733 9608
rect 5767 9605 5779 9639
rect 5721 9599 5779 9605
rect 5442 9568 5448 9580
rect 4479 9472 4844 9500
rect 4908 9540 5448 9568
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 4908 9432 4936 9540
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 6104 9568 6132 9676
rect 8662 9664 8668 9676
rect 8720 9664 8726 9716
rect 9122 9704 9128 9716
rect 8772 9676 9128 9704
rect 8772 9636 8800 9676
rect 9122 9664 9128 9676
rect 9180 9704 9186 9716
rect 10134 9704 10140 9716
rect 9180 9676 9720 9704
rect 10047 9676 10140 9704
rect 9180 9664 9186 9676
rect 8312 9608 8800 9636
rect 9692 9636 9720 9676
rect 10134 9664 10140 9676
rect 10192 9704 10198 9716
rect 11882 9704 11888 9716
rect 10192 9676 11888 9704
rect 10192 9664 10198 9676
rect 11882 9664 11888 9676
rect 11940 9664 11946 9716
rect 13078 9664 13084 9716
rect 13136 9704 13142 9716
rect 13817 9707 13875 9713
rect 13817 9704 13829 9707
rect 13136 9676 13829 9704
rect 13136 9664 13142 9676
rect 13817 9673 13829 9676
rect 13863 9673 13875 9707
rect 13817 9667 13875 9673
rect 15102 9664 15108 9716
rect 15160 9704 15166 9716
rect 16574 9704 16580 9716
rect 15160 9676 16580 9704
rect 15160 9664 15166 9676
rect 16574 9664 16580 9676
rect 16632 9664 16638 9716
rect 16758 9664 16764 9716
rect 16816 9704 16822 9716
rect 16816 9676 18184 9704
rect 16816 9664 16822 9676
rect 18156 9648 18184 9676
rect 11974 9636 11980 9648
rect 9692 9608 11100 9636
rect 11935 9608 11980 9636
rect 6181 9571 6239 9577
rect 6181 9568 6193 9571
rect 6104 9540 6193 9568
rect 6181 9537 6193 9540
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 6273 9571 6331 9577
rect 6273 9537 6285 9571
rect 6319 9537 6331 9571
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 6273 9531 6331 9537
rect 6656 9540 7113 9568
rect 5460 9500 5488 9528
rect 6288 9500 6316 9531
rect 6656 9512 6684 9540
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 6454 9500 6460 9512
rect 5460 9472 6460 9500
rect 6454 9460 6460 9472
rect 6512 9460 6518 9512
rect 6638 9460 6644 9512
rect 6696 9460 6702 9512
rect 7009 9503 7067 9509
rect 7009 9469 7021 9503
rect 7055 9469 7067 9503
rect 7009 9463 7067 9469
rect 7368 9503 7426 9509
rect 7368 9469 7380 9503
rect 7414 9500 7426 9503
rect 8312 9500 8340 9608
rect 9766 9528 9772 9580
rect 9824 9528 9830 9580
rect 11072 9577 11100 9608
rect 11974 9596 11980 9608
rect 12032 9596 12038 9648
rect 14369 9639 14427 9645
rect 14369 9605 14381 9639
rect 14415 9636 14427 9639
rect 15654 9636 15660 9648
rect 14415 9608 15660 9636
rect 14415 9605 14427 9608
rect 14369 9599 14427 9605
rect 15654 9596 15660 9608
rect 15712 9596 15718 9648
rect 16850 9596 16856 9648
rect 16908 9636 16914 9648
rect 17221 9639 17279 9645
rect 17221 9636 17233 9639
rect 16908 9608 17233 9636
rect 16908 9596 16914 9608
rect 17221 9605 17233 9608
rect 17267 9605 17279 9639
rect 17221 9599 17279 9605
rect 17494 9596 17500 9648
rect 17552 9636 17558 9648
rect 18049 9639 18107 9645
rect 18049 9636 18061 9639
rect 17552 9608 18061 9636
rect 17552 9596 17558 9608
rect 18049 9605 18061 9608
rect 18095 9605 18107 9639
rect 18049 9599 18107 9605
rect 18138 9596 18144 9648
rect 18196 9596 18202 9648
rect 19061 9639 19119 9645
rect 19061 9605 19073 9639
rect 19107 9636 19119 9639
rect 19150 9636 19156 9648
rect 19107 9608 19156 9636
rect 19107 9605 19119 9608
rect 19061 9599 19119 9605
rect 19150 9596 19156 9608
rect 19208 9596 19214 9648
rect 19886 9596 19892 9648
rect 19944 9636 19950 9648
rect 20073 9639 20131 9645
rect 20073 9636 20085 9639
rect 19944 9608 20085 9636
rect 19944 9596 19950 9608
rect 20073 9605 20085 9608
rect 20119 9605 20131 9639
rect 20073 9599 20131 9605
rect 11057 9571 11115 9577
rect 11057 9537 11069 9571
rect 11103 9568 11115 9571
rect 11146 9568 11152 9580
rect 11103 9540 11152 9568
rect 11103 9537 11115 9540
rect 11057 9531 11115 9537
rect 11146 9528 11152 9540
rect 11204 9528 11210 9580
rect 12250 9528 12256 9580
rect 12308 9568 12314 9580
rect 12437 9571 12495 9577
rect 12437 9568 12449 9571
rect 12308 9540 12449 9568
rect 12308 9528 12314 9540
rect 12437 9537 12449 9540
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 14182 9528 14188 9580
rect 14240 9568 14246 9580
rect 14921 9571 14979 9577
rect 14921 9568 14933 9571
rect 14240 9540 14933 9568
rect 14240 9528 14246 9540
rect 14921 9537 14933 9540
rect 14967 9537 14979 9571
rect 14921 9531 14979 9537
rect 15286 9528 15292 9580
rect 15344 9568 15350 9580
rect 15381 9571 15439 9577
rect 15381 9568 15393 9571
rect 15344 9540 15393 9568
rect 15344 9528 15350 9540
rect 15381 9537 15393 9540
rect 15427 9537 15439 9571
rect 15746 9568 15752 9580
rect 15381 9531 15439 9537
rect 15672 9540 15752 9568
rect 7414 9472 8340 9500
rect 8757 9503 8815 9509
rect 7414 9469 7426 9472
rect 7368 9463 7426 9469
rect 8757 9469 8769 9503
rect 8803 9500 8815 9503
rect 9306 9500 9312 9512
rect 8803 9472 9312 9500
rect 8803 9469 8815 9472
rect 8757 9463 8815 9469
rect 5074 9432 5080 9444
rect 2700 9404 4364 9432
rect 4632 9404 5080 9432
rect 4632 9376 4660 9404
rect 5074 9392 5080 9404
rect 5132 9392 5138 9444
rect 6089 9435 6147 9441
rect 6089 9401 6101 9435
rect 6135 9432 6147 9435
rect 6362 9432 6368 9444
rect 6135 9404 6368 9432
rect 6135 9401 6147 9404
rect 6089 9395 6147 9401
rect 6362 9392 6368 9404
rect 6420 9392 6426 9444
rect 7024 9432 7052 9463
rect 9306 9460 9312 9472
rect 9364 9500 9370 9512
rect 9784 9500 9812 9528
rect 9364 9472 9812 9500
rect 9364 9460 9370 9472
rect 9858 9460 9864 9512
rect 9916 9500 9922 9512
rect 10594 9500 10600 9512
rect 9916 9472 10600 9500
rect 9916 9460 9922 9472
rect 10594 9460 10600 9472
rect 10652 9500 10658 9512
rect 10873 9503 10931 9509
rect 10873 9500 10885 9503
rect 10652 9472 10885 9500
rect 10652 9460 10658 9472
rect 10873 9469 10885 9472
rect 10919 9469 10931 9503
rect 10873 9463 10931 9469
rect 11793 9503 11851 9509
rect 11793 9469 11805 9503
rect 11839 9500 11851 9503
rect 12342 9500 12348 9512
rect 11839 9472 12348 9500
rect 11839 9469 11851 9472
rect 11793 9463 11851 9469
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 12704 9503 12762 9509
rect 12704 9469 12716 9503
rect 12750 9500 12762 9503
rect 13630 9500 13636 9512
rect 12750 9472 13636 9500
rect 12750 9469 12762 9472
rect 12704 9463 12762 9469
rect 13630 9460 13636 9472
rect 13688 9460 13694 9512
rect 14274 9500 14280 9512
rect 14235 9472 14280 9500
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 14737 9503 14795 9509
rect 14737 9469 14749 9503
rect 14783 9500 14795 9503
rect 15672 9500 15700 9540
rect 15746 9528 15752 9540
rect 15804 9528 15810 9580
rect 15838 9528 15844 9580
rect 15896 9568 15902 9580
rect 15896 9540 15941 9568
rect 15896 9528 15902 9540
rect 17034 9528 17040 9580
rect 17092 9568 17098 9580
rect 18693 9571 18751 9577
rect 17092 9540 18644 9568
rect 17092 9528 17098 9540
rect 17586 9500 17592 9512
rect 14783 9472 15700 9500
rect 15764 9472 17592 9500
rect 14783 9469 14795 9472
rect 14737 9463 14795 9469
rect 7190 9432 7196 9444
rect 7024 9404 7196 9432
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 7282 9392 7288 9444
rect 7340 9432 7346 9444
rect 8846 9432 8852 9444
rect 7340 9404 7788 9432
rect 7340 9392 7346 9404
rect 2133 9367 2191 9373
rect 2133 9333 2145 9367
rect 2179 9333 2191 9367
rect 2498 9364 2504 9376
rect 2459 9336 2504 9364
rect 2133 9327 2191 9333
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 2593 9367 2651 9373
rect 2593 9333 2605 9367
rect 2639 9364 2651 9367
rect 3418 9364 3424 9376
rect 2639 9336 3424 9364
rect 2639 9333 2651 9336
rect 2593 9327 2651 9333
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 4522 9364 4528 9376
rect 3660 9336 3705 9364
rect 4483 9336 4528 9364
rect 3660 9324 3666 9336
rect 4522 9324 4528 9336
rect 4580 9324 4586 9376
rect 4614 9324 4620 9376
rect 4672 9324 4678 9376
rect 4890 9364 4896 9376
rect 4851 9336 4896 9364
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 5258 9364 5264 9376
rect 5219 9336 5264 9364
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5350 9324 5356 9376
rect 5408 9364 5414 9376
rect 5408 9336 5453 9364
rect 5408 9324 5414 9336
rect 6270 9324 6276 9376
rect 6328 9364 6334 9376
rect 6825 9367 6883 9373
rect 6825 9364 6837 9367
rect 6328 9336 6837 9364
rect 6328 9324 6334 9336
rect 6825 9333 6837 9336
rect 6871 9333 6883 9367
rect 7760 9364 7788 9404
rect 8496 9404 8852 9432
rect 8386 9364 8392 9376
rect 7760 9336 8392 9364
rect 6825 9327 6883 9333
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 8496 9373 8524 9404
rect 8846 9392 8852 9404
rect 8904 9392 8910 9444
rect 9024 9435 9082 9441
rect 9024 9401 9036 9435
rect 9070 9432 9082 9435
rect 9214 9432 9220 9444
rect 9070 9404 9220 9432
rect 9070 9401 9082 9404
rect 9024 9395 9082 9401
rect 9214 9392 9220 9404
rect 9272 9392 9278 9444
rect 9766 9392 9772 9444
rect 9824 9432 9830 9444
rect 10781 9435 10839 9441
rect 10781 9432 10793 9435
rect 9824 9404 10793 9432
rect 9824 9392 9830 9404
rect 10781 9401 10793 9404
rect 10827 9401 10839 9435
rect 10781 9395 10839 9401
rect 11054 9392 11060 9444
rect 11112 9432 11118 9444
rect 11974 9432 11980 9444
rect 11112 9404 11980 9432
rect 11112 9392 11118 9404
rect 11974 9392 11980 9404
rect 12032 9392 12038 9444
rect 12158 9392 12164 9444
rect 12216 9432 12222 9444
rect 15764 9432 15792 9472
rect 17586 9460 17592 9472
rect 17644 9460 17650 9512
rect 18138 9460 18144 9512
rect 18196 9500 18202 9512
rect 18509 9503 18567 9509
rect 18509 9500 18521 9503
rect 18196 9472 18521 9500
rect 18196 9460 18202 9472
rect 18509 9469 18521 9472
rect 18555 9469 18567 9503
rect 18616 9500 18644 9540
rect 18693 9537 18705 9571
rect 18739 9568 18751 9571
rect 18782 9568 18788 9580
rect 18739 9540 18788 9568
rect 18739 9537 18751 9540
rect 18693 9531 18751 9537
rect 18782 9528 18788 9540
rect 18840 9528 18846 9580
rect 19426 9528 19432 9580
rect 19484 9568 19490 9580
rect 19521 9571 19579 9577
rect 19521 9568 19533 9571
rect 19484 9540 19533 9568
rect 19484 9528 19490 9540
rect 19521 9537 19533 9540
rect 19567 9537 19579 9571
rect 19521 9531 19579 9537
rect 19613 9571 19671 9577
rect 19613 9537 19625 9571
rect 19659 9537 19671 9571
rect 19613 9531 19671 9537
rect 19628 9500 19656 9531
rect 20438 9528 20444 9580
rect 20496 9568 20502 9580
rect 20625 9571 20683 9577
rect 20625 9568 20637 9571
rect 20496 9540 20637 9568
rect 20496 9528 20502 9540
rect 20625 9537 20637 9540
rect 20671 9537 20683 9571
rect 20625 9531 20683 9537
rect 18616 9472 19656 9500
rect 18509 9463 18567 9469
rect 20162 9460 20168 9512
rect 20220 9500 20226 9512
rect 20530 9500 20536 9512
rect 20220 9472 20536 9500
rect 20220 9460 20226 9472
rect 20530 9460 20536 9472
rect 20588 9460 20594 9512
rect 12216 9404 15792 9432
rect 16108 9435 16166 9441
rect 12216 9392 12222 9404
rect 16108 9401 16120 9435
rect 16154 9432 16166 9435
rect 16298 9432 16304 9444
rect 16154 9404 16304 9432
rect 16154 9401 16166 9404
rect 16108 9395 16166 9401
rect 16298 9392 16304 9404
rect 16356 9392 16362 9444
rect 17497 9435 17555 9441
rect 17497 9401 17509 9435
rect 17543 9432 17555 9435
rect 18417 9435 18475 9441
rect 18417 9432 18429 9435
rect 17543 9404 18429 9432
rect 17543 9401 17555 9404
rect 17497 9395 17555 9401
rect 18417 9401 18429 9404
rect 18463 9401 18475 9435
rect 18417 9395 18475 9401
rect 8481 9367 8539 9373
rect 8481 9333 8493 9367
rect 8527 9333 8539 9367
rect 8481 9327 8539 9333
rect 10410 9324 10416 9376
rect 10468 9364 10474 9376
rect 10468 9336 10513 9364
rect 10468 9324 10474 9336
rect 10594 9324 10600 9376
rect 10652 9364 10658 9376
rect 13078 9364 13084 9376
rect 10652 9336 13084 9364
rect 10652 9324 10658 9336
rect 13078 9324 13084 9336
rect 13136 9324 13142 9376
rect 14093 9367 14151 9373
rect 14093 9333 14105 9367
rect 14139 9364 14151 9367
rect 14550 9364 14556 9376
rect 14139 9336 14556 9364
rect 14139 9333 14151 9336
rect 14093 9327 14151 9333
rect 14550 9324 14556 9336
rect 14608 9324 14614 9376
rect 14829 9367 14887 9373
rect 14829 9333 14841 9367
rect 14875 9364 14887 9367
rect 17862 9364 17868 9376
rect 14875 9336 17868 9364
rect 14875 9333 14887 9336
rect 14829 9327 14887 9333
rect 17862 9324 17868 9336
rect 17920 9324 17926 9376
rect 19426 9364 19432 9376
rect 19387 9336 19432 9364
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 20438 9364 20444 9376
rect 20399 9336 20444 9364
rect 20438 9324 20444 9336
rect 20496 9324 20502 9376
rect 20530 9324 20536 9376
rect 20588 9364 20594 9376
rect 20588 9336 20633 9364
rect 20588 9324 20594 9336
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 2406 9160 2412 9172
rect 2367 9132 2412 9160
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 2961 9163 3019 9169
rect 2961 9160 2973 9163
rect 2832 9132 2973 9160
rect 2832 9120 2838 9132
rect 2961 9129 2973 9132
rect 3007 9129 3019 9163
rect 2961 9123 3019 9129
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 3476 9132 4077 9160
rect 3476 9120 3482 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 4522 9120 4528 9172
rect 4580 9160 4586 9172
rect 5166 9160 5172 9172
rect 4580 9132 5172 9160
rect 4580 9120 4586 9132
rect 5166 9120 5172 9132
rect 5224 9120 5230 9172
rect 6178 9160 6184 9172
rect 5276 9132 6184 9160
rect 2314 9092 2320 9104
rect 2275 9064 2320 9092
rect 2314 9052 2320 9064
rect 2372 9052 2378 9104
rect 3329 9095 3387 9101
rect 3329 9061 3341 9095
rect 3375 9092 3387 9095
rect 3786 9092 3792 9104
rect 3375 9064 3792 9092
rect 3375 9061 3387 9064
rect 3329 9055 3387 9061
rect 3786 9052 3792 9064
rect 3844 9052 3850 9104
rect 3878 9052 3884 9104
rect 3936 9092 3942 9104
rect 4433 9095 4491 9101
rect 4433 9092 4445 9095
rect 3936 9064 4445 9092
rect 3936 9052 3942 9064
rect 4433 9061 4445 9064
rect 4479 9092 4491 9095
rect 5276 9092 5304 9132
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 6454 9160 6460 9172
rect 6415 9132 6460 9160
rect 6454 9120 6460 9132
rect 6512 9120 6518 9172
rect 7193 9163 7251 9169
rect 7193 9129 7205 9163
rect 7239 9160 7251 9163
rect 7466 9160 7472 9172
rect 7239 9132 7472 9160
rect 7239 9129 7251 9132
rect 7193 9123 7251 9129
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 7742 9120 7748 9172
rect 7800 9120 7806 9172
rect 9214 9160 9220 9172
rect 7852 9132 8975 9160
rect 9175 9132 9220 9160
rect 4479 9064 5304 9092
rect 5344 9095 5402 9101
rect 4479 9061 4491 9064
rect 4433 9055 4491 9061
rect 5344 9061 5356 9095
rect 5390 9092 5402 9095
rect 5442 9092 5448 9104
rect 5390 9064 5448 9092
rect 5390 9061 5402 9064
rect 5344 9055 5402 9061
rect 5442 9052 5448 9064
rect 5500 9092 5506 9104
rect 5500 9064 6316 9092
rect 5500 9052 5506 9064
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 1670 9024 1676 9036
rect 1443 8996 1676 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 4525 9027 4583 9033
rect 4525 8993 4537 9027
rect 4571 9024 4583 9027
rect 4571 8996 4752 9024
rect 4571 8993 4583 8996
rect 4525 8987 4583 8993
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8956 2651 8959
rect 2682 8956 2688 8968
rect 2639 8928 2688 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 3418 8956 3424 8968
rect 3379 8928 3424 8956
rect 3418 8916 3424 8928
rect 3476 8916 3482 8968
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8956 3571 8959
rect 4154 8956 4160 8968
rect 3559 8928 4160 8956
rect 3559 8925 3571 8928
rect 3513 8919 3571 8925
rect 1581 8891 1639 8897
rect 1581 8857 1593 8891
rect 1627 8888 1639 8891
rect 3050 8888 3056 8900
rect 1627 8860 3056 8888
rect 1627 8857 1639 8860
rect 1581 8851 1639 8857
rect 3050 8848 3056 8860
rect 3108 8848 3114 8900
rect 3234 8848 3240 8900
rect 3292 8888 3298 8900
rect 3528 8888 3556 8919
rect 4154 8916 4160 8928
rect 4212 8956 4218 8968
rect 4614 8956 4620 8968
rect 4212 8928 4620 8956
rect 4212 8916 4218 8928
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 3292 8860 3556 8888
rect 3292 8848 3298 8860
rect 4724 8820 4752 8996
rect 4890 8984 4896 9036
rect 4948 9024 4954 9036
rect 5077 9027 5135 9033
rect 5077 9024 5089 9027
rect 4948 8996 5089 9024
rect 4948 8984 4954 8996
rect 5077 8993 5089 8996
rect 5123 9024 5135 9027
rect 6178 9024 6184 9036
rect 5123 8996 6184 9024
rect 5123 8993 5135 8996
rect 5077 8987 5135 8993
rect 6178 8984 6184 8996
rect 6236 8984 6242 9036
rect 6288 8956 6316 9064
rect 6362 9052 6368 9104
rect 6420 9092 6426 9104
rect 7760 9092 7788 9120
rect 6420 9064 7788 9092
rect 6420 9052 6426 9064
rect 7101 9027 7159 9033
rect 7101 8993 7113 9027
rect 7147 9024 7159 9027
rect 7147 8996 7696 9024
rect 7147 8993 7159 8996
rect 7101 8987 7159 8993
rect 7285 8959 7343 8965
rect 7285 8956 7297 8959
rect 6288 8928 7297 8956
rect 7285 8925 7297 8928
rect 7331 8925 7343 8959
rect 7668 8956 7696 8996
rect 7742 8984 7748 9036
rect 7800 9024 7806 9036
rect 7852 9033 7880 9132
rect 8104 9095 8162 9101
rect 8104 9061 8116 9095
rect 8150 9092 8162 9095
rect 8846 9092 8852 9104
rect 8150 9064 8852 9092
rect 8150 9061 8162 9064
rect 8104 9055 8162 9061
rect 8846 9052 8852 9064
rect 8904 9052 8910 9104
rect 8947 9092 8975 9132
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 10045 9163 10103 9169
rect 10045 9129 10057 9163
rect 10091 9160 10103 9163
rect 10410 9160 10416 9172
rect 10091 9132 10416 9160
rect 10091 9129 10103 9132
rect 10045 9123 10103 9129
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 10686 9120 10692 9172
rect 10744 9160 10750 9172
rect 11790 9160 11796 9172
rect 10744 9132 11796 9160
rect 10744 9120 10750 9132
rect 11790 9120 11796 9132
rect 11848 9120 11854 9172
rect 12434 9120 12440 9172
rect 12492 9160 12498 9172
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 12492 9132 13001 9160
rect 12492 9120 12498 9132
rect 12989 9129 13001 9132
rect 13035 9129 13047 9163
rect 14090 9160 14096 9172
rect 12989 9123 13047 9129
rect 13464 9132 14096 9160
rect 9306 9092 9312 9104
rect 8947 9064 9312 9092
rect 9306 9052 9312 9064
rect 9364 9052 9370 9104
rect 9950 9052 9956 9104
rect 10008 9092 10014 9104
rect 10137 9095 10195 9101
rect 10137 9092 10149 9095
rect 10008 9064 10149 9092
rect 10008 9052 10014 9064
rect 10137 9061 10149 9064
rect 10183 9061 10195 9095
rect 12342 9092 12348 9104
rect 10137 9055 10195 9061
rect 10888 9064 12348 9092
rect 7837 9027 7895 9033
rect 7837 9024 7849 9027
rect 7800 8996 7849 9024
rect 7800 8984 7806 8996
rect 7837 8993 7849 8996
rect 7883 8993 7895 9027
rect 8386 9024 8392 9036
rect 7837 8987 7895 8993
rect 7944 8996 8392 9024
rect 7944 8956 7972 8996
rect 8386 8984 8392 8996
rect 8444 9024 8450 9036
rect 9858 9024 9864 9036
rect 8444 8996 9864 9024
rect 8444 8984 8450 8996
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 10594 8984 10600 9036
rect 10652 9024 10658 9036
rect 10888 9033 10916 9064
rect 12342 9052 12348 9064
rect 12400 9052 12406 9104
rect 12897 9095 12955 9101
rect 12897 9061 12909 9095
rect 12943 9092 12955 9095
rect 13464 9092 13492 9132
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 14829 9163 14887 9169
rect 14829 9129 14841 9163
rect 14875 9160 14887 9163
rect 15194 9160 15200 9172
rect 14875 9132 15200 9160
rect 14875 9129 14887 9132
rect 14829 9123 14887 9129
rect 15194 9120 15200 9132
rect 15252 9120 15258 9172
rect 15838 9120 15844 9172
rect 15896 9160 15902 9172
rect 16301 9163 16359 9169
rect 16301 9160 16313 9163
rect 15896 9132 16313 9160
rect 15896 9120 15902 9132
rect 16301 9129 16313 9132
rect 16347 9129 16359 9163
rect 16301 9123 16359 9129
rect 16482 9120 16488 9172
rect 16540 9160 16546 9172
rect 18138 9160 18144 9172
rect 16540 9132 18144 9160
rect 16540 9120 16546 9132
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 19610 9160 19616 9172
rect 18432 9132 18736 9160
rect 19571 9132 19616 9160
rect 12943 9064 13492 9092
rect 14001 9095 14059 9101
rect 12943 9061 12955 9064
rect 12897 9055 12955 9061
rect 14001 9061 14013 9095
rect 14047 9092 14059 9095
rect 15286 9092 15292 9104
rect 14047 9064 15292 9092
rect 14047 9061 14059 9064
rect 14001 9055 14059 9061
rect 15286 9052 15292 9064
rect 15344 9052 15350 9104
rect 15562 9052 15568 9104
rect 15620 9092 15626 9104
rect 15749 9095 15807 9101
rect 15749 9092 15761 9095
rect 15620 9064 15761 9092
rect 15620 9052 15626 9064
rect 15749 9061 15761 9064
rect 15795 9061 15807 9095
rect 15749 9055 15807 9061
rect 16117 9095 16175 9101
rect 16117 9061 16129 9095
rect 16163 9092 16175 9095
rect 18432 9092 18460 9132
rect 16163 9064 18460 9092
rect 18500 9095 18558 9101
rect 16163 9061 16175 9064
rect 16117 9055 16175 9061
rect 18500 9061 18512 9095
rect 18546 9092 18558 9095
rect 18598 9092 18604 9104
rect 18546 9064 18604 9092
rect 18546 9061 18558 9064
rect 18500 9055 18558 9061
rect 18598 9052 18604 9064
rect 18656 9052 18662 9104
rect 18708 9092 18736 9132
rect 19610 9120 19616 9132
rect 19668 9120 19674 9172
rect 20898 9092 20904 9104
rect 18708 9064 20904 9092
rect 20898 9052 20904 9064
rect 20956 9052 20962 9104
rect 10873 9027 10931 9033
rect 10873 9024 10885 9027
rect 10652 8996 10885 9024
rect 10652 8984 10658 8996
rect 10873 8993 10885 8996
rect 10919 8993 10931 9027
rect 10873 8987 10931 8993
rect 11140 9027 11198 9033
rect 11140 8993 11152 9027
rect 11186 9024 11198 9027
rect 12986 9024 12992 9036
rect 11186 8996 12992 9024
rect 11186 8993 11198 8996
rect 11140 8987 11198 8993
rect 12986 8984 12992 8996
rect 13044 8984 13050 9036
rect 13909 9027 13967 9033
rect 13909 8993 13921 9027
rect 13955 9024 13967 9027
rect 14458 9024 14464 9036
rect 13955 8996 14464 9024
rect 13955 8993 13967 8996
rect 13909 8987 13967 8993
rect 14458 8984 14464 8996
rect 14516 8984 14522 9036
rect 14645 9027 14703 9033
rect 14645 8993 14657 9027
rect 14691 9024 14703 9027
rect 15010 9024 15016 9036
rect 14691 8996 15016 9024
rect 14691 8993 14703 8996
rect 14645 8987 14703 8993
rect 15010 8984 15016 8996
rect 15068 8984 15074 9036
rect 15105 9027 15163 9033
rect 15105 8993 15117 9027
rect 15151 9024 15163 9027
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 15151 8996 15669 9024
rect 15151 8993 15163 8996
rect 15105 8987 15163 8993
rect 15657 8993 15669 8996
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 16574 8984 16580 9036
rect 16632 9024 16638 9036
rect 16669 9027 16727 9033
rect 16669 9024 16681 9027
rect 16632 8996 16681 9024
rect 16632 8984 16638 8996
rect 16669 8993 16681 8996
rect 16715 8993 16727 9027
rect 16669 8987 16727 8993
rect 16761 9027 16819 9033
rect 16761 8993 16773 9027
rect 16807 9024 16819 9027
rect 16942 9024 16948 9036
rect 16807 8996 16948 9024
rect 16807 8993 16819 8996
rect 16761 8987 16819 8993
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 17494 9024 17500 9036
rect 17455 8996 17500 9024
rect 17494 8984 17500 8996
rect 17552 8984 17558 9036
rect 17954 9024 17960 9036
rect 17880 8996 17960 9024
rect 7668 8928 7972 8956
rect 7285 8919 7343 8925
rect 8846 8916 8852 8968
rect 8904 8956 8910 8968
rect 10134 8956 10140 8968
rect 8904 8928 10140 8956
rect 8904 8916 8910 8928
rect 10134 8916 10140 8928
rect 10192 8956 10198 8968
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 10192 8928 10241 8956
rect 10192 8916 10198 8928
rect 10229 8925 10241 8928
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8956 12495 8959
rect 13081 8959 13139 8965
rect 13081 8956 13093 8959
rect 12483 8928 13093 8956
rect 12483 8925 12495 8928
rect 12437 8919 12495 8925
rect 13081 8925 13093 8928
rect 13127 8925 13139 8959
rect 13081 8919 13139 8925
rect 13998 8916 14004 8968
rect 14056 8956 14062 8968
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 14056 8928 14105 8956
rect 14056 8916 14062 8928
rect 14093 8925 14105 8928
rect 14139 8925 14151 8959
rect 14093 8919 14151 8925
rect 14274 8916 14280 8968
rect 14332 8956 14338 8968
rect 15841 8959 15899 8965
rect 15841 8956 15853 8959
rect 14332 8928 15853 8956
rect 14332 8916 14338 8928
rect 15841 8925 15853 8928
rect 15887 8956 15899 8959
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 15887 8928 16865 8956
rect 15887 8925 15899 8928
rect 15841 8919 15899 8925
rect 16853 8925 16865 8928
rect 16899 8956 16911 8959
rect 17126 8956 17132 8968
rect 16899 8928 17132 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 17681 8959 17739 8965
rect 17681 8925 17693 8959
rect 17727 8925 17739 8959
rect 17681 8919 17739 8925
rect 6362 8848 6368 8900
rect 6420 8888 6426 8900
rect 6420 8860 6868 8888
rect 6420 8848 6426 8860
rect 4982 8820 4988 8832
rect 4724 8792 4988 8820
rect 4982 8780 4988 8792
rect 5040 8820 5046 8832
rect 5350 8820 5356 8832
rect 5040 8792 5356 8820
rect 5040 8780 5046 8792
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 6638 8780 6644 8832
rect 6696 8820 6702 8832
rect 6733 8823 6791 8829
rect 6733 8820 6745 8823
rect 6696 8792 6745 8820
rect 6696 8780 6702 8792
rect 6733 8789 6745 8792
rect 6779 8789 6791 8823
rect 6840 8820 6868 8860
rect 8938 8848 8944 8900
rect 8996 8888 9002 8900
rect 9214 8888 9220 8900
rect 8996 8860 9220 8888
rect 8996 8848 9002 8860
rect 9214 8848 9220 8860
rect 9272 8848 9278 8900
rect 13906 8888 13912 8900
rect 11808 8860 13912 8888
rect 8570 8820 8576 8832
rect 6840 8792 8576 8820
rect 6733 8783 6791 8789
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 8846 8780 8852 8832
rect 8904 8820 8910 8832
rect 9677 8823 9735 8829
rect 9677 8820 9689 8823
rect 8904 8792 9689 8820
rect 8904 8780 8910 8792
rect 9677 8789 9689 8792
rect 9723 8789 9735 8823
rect 9677 8783 9735 8789
rect 9858 8780 9864 8832
rect 9916 8820 9922 8832
rect 11808 8820 11836 8860
rect 13906 8848 13912 8860
rect 13964 8848 13970 8900
rect 15289 8891 15347 8897
rect 15289 8888 15301 8891
rect 14752 8860 15301 8888
rect 9916 8792 11836 8820
rect 9916 8780 9922 8792
rect 12158 8780 12164 8832
rect 12216 8820 12222 8832
rect 12253 8823 12311 8829
rect 12253 8820 12265 8823
rect 12216 8792 12265 8820
rect 12216 8780 12222 8792
rect 12253 8789 12265 8792
rect 12299 8820 12311 8823
rect 12437 8823 12495 8829
rect 12437 8820 12449 8823
rect 12299 8792 12449 8820
rect 12299 8789 12311 8792
rect 12253 8783 12311 8789
rect 12437 8789 12449 8792
rect 12483 8789 12495 8823
rect 12437 8783 12495 8789
rect 12529 8823 12587 8829
rect 12529 8789 12541 8823
rect 12575 8820 12587 8823
rect 12618 8820 12624 8832
rect 12575 8792 12624 8820
rect 12575 8789 12587 8792
rect 12529 8783 12587 8789
rect 12618 8780 12624 8792
rect 12676 8780 12682 8832
rect 13446 8780 13452 8832
rect 13504 8820 13510 8832
rect 13541 8823 13599 8829
rect 13541 8820 13553 8823
rect 13504 8792 13553 8820
rect 13504 8780 13510 8792
rect 13541 8789 13553 8792
rect 13587 8789 13599 8823
rect 13541 8783 13599 8789
rect 13630 8780 13636 8832
rect 13688 8820 13694 8832
rect 14752 8820 14780 8860
rect 15289 8857 15301 8860
rect 15335 8857 15347 8891
rect 16117 8891 16175 8897
rect 16117 8888 16129 8891
rect 15289 8851 15347 8857
rect 15856 8860 16129 8888
rect 15856 8832 15884 8860
rect 16117 8857 16129 8860
rect 16163 8857 16175 8891
rect 16117 8851 16175 8857
rect 16298 8848 16304 8900
rect 16356 8888 16362 8900
rect 17696 8888 17724 8919
rect 16356 8860 17724 8888
rect 16356 8848 16362 8860
rect 13688 8792 14780 8820
rect 13688 8780 13694 8792
rect 14918 8780 14924 8832
rect 14976 8820 14982 8832
rect 15105 8823 15163 8829
rect 15105 8820 15117 8823
rect 14976 8792 15117 8820
rect 14976 8780 14982 8792
rect 15105 8789 15117 8792
rect 15151 8789 15163 8823
rect 15105 8783 15163 8789
rect 15838 8780 15844 8832
rect 15896 8780 15902 8832
rect 16022 8780 16028 8832
rect 16080 8820 16086 8832
rect 17880 8820 17908 8996
rect 17954 8984 17960 8996
rect 18012 8984 18018 9036
rect 18233 9027 18291 9033
rect 18233 8993 18245 9027
rect 18279 9024 18291 9027
rect 18322 9024 18328 9036
rect 18279 8996 18328 9024
rect 18279 8993 18291 8996
rect 18233 8987 18291 8993
rect 18322 8984 18328 8996
rect 18380 8984 18386 9036
rect 19889 9027 19947 9033
rect 19889 8993 19901 9027
rect 19935 9024 19947 9027
rect 19978 9024 19984 9036
rect 19935 8996 19984 9024
rect 19935 8993 19947 8996
rect 19889 8987 19947 8993
rect 19978 8984 19984 8996
rect 20036 8984 20042 9036
rect 19334 8916 19340 8968
rect 19392 8956 19398 8968
rect 20073 8959 20131 8965
rect 20073 8956 20085 8959
rect 19392 8928 20085 8956
rect 19392 8916 19398 8928
rect 20073 8925 20085 8928
rect 20119 8925 20131 8959
rect 20073 8919 20131 8925
rect 18138 8848 18144 8900
rect 18196 8848 18202 8900
rect 16080 8792 17908 8820
rect 18156 8820 18184 8848
rect 19150 8820 19156 8832
rect 18156 8792 19156 8820
rect 16080 8780 16086 8792
rect 19150 8780 19156 8792
rect 19208 8780 19214 8832
rect 19886 8780 19892 8832
rect 19944 8820 19950 8832
rect 20714 8820 20720 8832
rect 19944 8792 20720 8820
rect 19944 8780 19950 8792
rect 20714 8780 20720 8792
rect 20772 8780 20778 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 2409 8619 2467 8625
rect 2409 8585 2421 8619
rect 2455 8616 2467 8619
rect 2498 8616 2504 8628
rect 2455 8588 2504 8616
rect 2455 8585 2467 8588
rect 2409 8579 2467 8585
rect 2498 8576 2504 8588
rect 2556 8576 2562 8628
rect 3605 8619 3663 8625
rect 3605 8585 3617 8619
rect 3651 8616 3663 8619
rect 3970 8616 3976 8628
rect 3651 8588 3976 8616
rect 3651 8585 3663 8588
rect 3605 8579 3663 8585
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 5166 8576 5172 8628
rect 5224 8616 5230 8628
rect 5721 8619 5779 8625
rect 5721 8616 5733 8619
rect 5224 8588 5733 8616
rect 5224 8576 5230 8588
rect 5721 8585 5733 8588
rect 5767 8585 5779 8619
rect 5721 8579 5779 8585
rect 6178 8576 6184 8628
rect 6236 8616 6242 8628
rect 6546 8616 6552 8628
rect 6236 8588 6552 8616
rect 6236 8576 6242 8588
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 6638 8576 6644 8628
rect 6696 8576 6702 8628
rect 7742 8616 7748 8628
rect 6840 8588 7748 8616
rect 3418 8548 3424 8560
rect 1872 8520 3424 8548
rect 1872 8489 1900 8520
rect 3418 8508 3424 8520
rect 3476 8548 3482 8560
rect 3786 8548 3792 8560
rect 3476 8520 3792 8548
rect 3476 8508 3482 8520
rect 3786 8508 3792 8520
rect 3844 8508 3850 8560
rect 5442 8548 5448 8560
rect 5403 8520 5448 8548
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 6656 8548 6684 8576
rect 6196 8520 6684 8548
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8449 1915 8483
rect 2038 8480 2044 8492
rect 1999 8452 2044 8480
rect 1857 8443 1915 8449
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8480 3019 8483
rect 3234 8480 3240 8492
rect 3007 8452 3240 8480
rect 3007 8449 3019 8452
rect 2961 8443 3019 8449
rect 3234 8440 3240 8452
rect 3292 8440 3298 8492
rect 6196 8489 6224 8520
rect 6840 8489 6868 8588
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 8202 8576 8208 8628
rect 8260 8616 8266 8628
rect 12253 8619 12311 8625
rect 12253 8616 12265 8619
rect 8260 8588 12265 8616
rect 8260 8576 8266 8588
rect 12253 8585 12265 8588
rect 12299 8585 12311 8619
rect 12253 8579 12311 8585
rect 12437 8619 12495 8625
rect 12437 8585 12449 8619
rect 12483 8616 12495 8619
rect 12526 8616 12532 8628
rect 12483 8588 12532 8616
rect 12483 8585 12495 8588
rect 12437 8579 12495 8585
rect 12526 8576 12532 8588
rect 12584 8576 12590 8628
rect 13630 8616 13636 8628
rect 12728 8588 13636 8616
rect 7834 8508 7840 8560
rect 7892 8548 7898 8560
rect 9858 8548 9864 8560
rect 7892 8520 9864 8548
rect 7892 8508 7898 8520
rect 8220 8492 8248 8520
rect 9858 8508 9864 8520
rect 9916 8508 9922 8560
rect 10029 8520 11928 8548
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8449 6239 8483
rect 6181 8443 6239 8449
rect 6273 8483 6331 8489
rect 6273 8449 6285 8483
rect 6319 8449 6331 8483
rect 6273 8443 6331 8449
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8449 6883 8483
rect 6825 8443 6883 8449
rect 1394 8372 1400 8424
rect 1452 8412 1458 8424
rect 1765 8415 1823 8421
rect 1765 8412 1777 8415
rect 1452 8384 1777 8412
rect 1452 8372 1458 8384
rect 1765 8381 1777 8384
rect 1811 8381 1823 8415
rect 1765 8375 1823 8381
rect 2777 8415 2835 8421
rect 2777 8381 2789 8415
rect 2823 8412 2835 8415
rect 3050 8412 3056 8424
rect 2823 8384 3056 8412
rect 2823 8381 2835 8384
rect 2777 8375 2835 8381
rect 3050 8372 3056 8384
rect 3108 8412 3114 8424
rect 3326 8412 3332 8424
rect 3108 8384 3332 8412
rect 3108 8372 3114 8384
rect 3326 8372 3332 8384
rect 3384 8372 3390 8424
rect 3421 8415 3479 8421
rect 3421 8381 3433 8415
rect 3467 8412 3479 8415
rect 3694 8412 3700 8424
rect 3467 8384 3700 8412
rect 3467 8381 3479 8384
rect 3421 8375 3479 8381
rect 3694 8372 3700 8384
rect 3752 8372 3758 8424
rect 4062 8412 4068 8424
rect 3975 8384 4068 8412
rect 4062 8372 4068 8384
rect 4120 8412 4126 8424
rect 4890 8412 4896 8424
rect 4120 8384 4896 8412
rect 4120 8372 4126 8384
rect 4890 8372 4896 8384
rect 4948 8372 4954 8424
rect 5074 8372 5080 8424
rect 5132 8412 5138 8424
rect 6288 8412 6316 8443
rect 8202 8440 8208 8492
rect 8260 8440 8266 8492
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 8570 8480 8576 8492
rect 8444 8452 8576 8480
rect 8444 8440 8450 8452
rect 8570 8440 8576 8452
rect 8628 8440 8634 8492
rect 9030 8480 9036 8492
rect 8991 8452 9036 8480
rect 9030 8440 9036 8452
rect 9088 8440 9094 8492
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8480 9459 8483
rect 10029 8480 10057 8520
rect 10134 8480 10140 8492
rect 9447 8452 10057 8480
rect 10095 8452 10140 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 10134 8440 10140 8452
rect 10192 8440 10198 8492
rect 11054 8480 11060 8492
rect 11015 8452 11060 8480
rect 11054 8440 11060 8452
rect 11112 8440 11118 8492
rect 11900 8480 11928 8520
rect 11974 8508 11980 8560
rect 12032 8548 12038 8560
rect 12032 8520 12077 8548
rect 12032 8508 12038 8520
rect 12728 8480 12756 8588
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 13906 8576 13912 8628
rect 13964 8616 13970 8628
rect 18506 8616 18512 8628
rect 13964 8588 18512 8616
rect 13964 8576 13970 8588
rect 18506 8576 18512 8588
rect 18564 8576 18570 8628
rect 19058 8616 19064 8628
rect 19019 8588 19064 8616
rect 19058 8576 19064 8588
rect 19116 8576 19122 8628
rect 19702 8576 19708 8628
rect 19760 8576 19766 8628
rect 20073 8619 20131 8625
rect 20073 8585 20085 8619
rect 20119 8616 20131 8619
rect 20438 8616 20444 8628
rect 20119 8588 20444 8616
rect 20119 8585 20131 8588
rect 20073 8579 20131 8585
rect 20438 8576 20444 8588
rect 20496 8576 20502 8628
rect 12802 8508 12808 8560
rect 12860 8548 12866 8560
rect 13449 8551 13507 8557
rect 13449 8548 13461 8551
rect 12860 8520 13461 8548
rect 12860 8508 12866 8520
rect 13449 8517 13461 8520
rect 13495 8517 13507 8551
rect 14458 8548 14464 8560
rect 14419 8520 14464 8548
rect 13449 8511 13507 8517
rect 14458 8508 14464 8520
rect 14516 8508 14522 8560
rect 17126 8508 17132 8560
rect 17184 8548 17190 8560
rect 17497 8551 17555 8557
rect 17497 8548 17509 8551
rect 17184 8520 17509 8548
rect 17184 8508 17190 8520
rect 17497 8517 17509 8520
rect 17543 8517 17555 8551
rect 17497 8511 17555 8517
rect 18049 8551 18107 8557
rect 18049 8517 18061 8551
rect 18095 8548 18107 8551
rect 19426 8548 19432 8560
rect 18095 8520 19432 8548
rect 18095 8517 18107 8520
rect 18049 8511 18107 8517
rect 12897 8483 12955 8489
rect 12897 8480 12909 8483
rect 11900 8452 12909 8480
rect 12897 8449 12909 8452
rect 12943 8449 12955 8483
rect 13078 8480 13084 8492
rect 13039 8452 13084 8480
rect 12897 8443 12955 8449
rect 13078 8440 13084 8452
rect 13136 8480 13142 8492
rect 13538 8480 13544 8492
rect 13136 8452 13544 8480
rect 13136 8440 13142 8452
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 14090 8480 14096 8492
rect 14051 8452 14096 8480
rect 14090 8440 14096 8452
rect 14148 8480 14154 8492
rect 14274 8480 14280 8492
rect 14148 8452 14280 8480
rect 14148 8440 14154 8452
rect 14274 8440 14280 8452
rect 14332 8440 14338 8492
rect 14366 8440 14372 8492
rect 14424 8480 14430 8492
rect 14921 8483 14979 8489
rect 14921 8480 14933 8483
rect 14424 8452 14933 8480
rect 14424 8440 14430 8452
rect 14921 8449 14933 8452
rect 14967 8449 14979 8483
rect 14921 8443 14979 8449
rect 15010 8440 15016 8492
rect 15068 8480 15074 8492
rect 15068 8452 15113 8480
rect 15068 8440 15074 8452
rect 15746 8440 15752 8492
rect 15804 8480 15810 8492
rect 17512 8480 17540 8511
rect 19426 8508 19432 8520
rect 19484 8508 19490 8560
rect 19720 8548 19748 8576
rect 19720 8520 20668 8548
rect 18414 8480 18420 8492
rect 15804 8452 16252 8480
rect 17512 8452 18420 8480
rect 15804 8440 15810 8452
rect 5132 8384 6316 8412
rect 5132 8372 5138 8384
rect 6454 8372 6460 8424
rect 6512 8412 6518 8424
rect 8846 8412 8852 8424
rect 6512 8384 8708 8412
rect 8807 8384 8852 8412
rect 6512 8372 6518 8384
rect 2869 8347 2927 8353
rect 2869 8313 2881 8347
rect 2915 8344 2927 8347
rect 4154 8344 4160 8356
rect 2915 8316 4160 8344
rect 2915 8313 2927 8316
rect 2869 8307 2927 8313
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 4338 8353 4344 8356
rect 4332 8344 4344 8353
rect 4299 8316 4344 8344
rect 4332 8307 4344 8316
rect 4338 8304 4344 8307
rect 4396 8304 4402 8356
rect 7098 8353 7104 8356
rect 7092 8307 7104 8353
rect 7156 8344 7162 8356
rect 8680 8344 8708 8384
rect 8846 8372 8852 8384
rect 8904 8372 8910 8424
rect 9122 8372 9128 8424
rect 9180 8412 9186 8424
rect 11072 8412 11100 8440
rect 11790 8412 11796 8424
rect 9180 8384 11100 8412
rect 11751 8384 11796 8412
rect 9180 8372 9186 8384
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8412 12311 8415
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 12299 8384 12817 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12805 8381 12817 8384
rect 12851 8412 12863 8415
rect 13722 8412 13728 8424
rect 12851 8384 13728 8412
rect 12851 8381 12863 8384
rect 12805 8375 12863 8381
rect 13722 8372 13728 8384
rect 13780 8372 13786 8424
rect 13906 8372 13912 8424
rect 13964 8412 13970 8424
rect 15102 8412 15108 8424
rect 13964 8384 15108 8412
rect 13964 8372 13970 8384
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 15562 8412 15568 8424
rect 15523 8384 15568 8412
rect 15562 8372 15568 8384
rect 15620 8372 15626 8424
rect 16022 8372 16028 8424
rect 16080 8412 16086 8424
rect 16117 8415 16175 8421
rect 16117 8412 16129 8415
rect 16080 8384 16129 8412
rect 16080 8372 16086 8384
rect 16117 8381 16129 8384
rect 16163 8381 16175 8415
rect 16224 8412 16252 8452
rect 18414 8440 18420 8452
rect 18472 8440 18478 8492
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8480 18659 8483
rect 18782 8480 18788 8492
rect 18647 8452 18788 8480
rect 18647 8449 18659 8452
rect 18601 8443 18659 8449
rect 18782 8440 18788 8452
rect 18840 8440 18846 8492
rect 18874 8440 18880 8492
rect 18932 8480 18938 8492
rect 19521 8483 19579 8489
rect 19521 8480 19533 8483
rect 18932 8452 19533 8480
rect 18932 8440 18938 8452
rect 19521 8449 19533 8452
rect 19567 8449 19579 8483
rect 19521 8443 19579 8449
rect 19705 8483 19763 8489
rect 19705 8449 19717 8483
rect 19751 8480 19763 8483
rect 20346 8480 20352 8492
rect 19751 8452 20352 8480
rect 19751 8449 19763 8452
rect 19705 8443 19763 8449
rect 20346 8440 20352 8452
rect 20404 8440 20410 8492
rect 20640 8489 20668 8520
rect 20625 8483 20683 8489
rect 20625 8449 20637 8483
rect 20671 8449 20683 8483
rect 20625 8443 20683 8449
rect 16384 8415 16442 8421
rect 16224 8384 16344 8412
rect 16117 8375 16175 8381
rect 9401 8347 9459 8353
rect 9401 8344 9413 8347
rect 7156 8316 7192 8344
rect 8680 8316 9413 8344
rect 7098 8304 7104 8307
rect 7156 8304 7162 8316
rect 9401 8313 9413 8316
rect 9447 8313 9459 8347
rect 9401 8307 9459 8313
rect 9861 8347 9919 8353
rect 9861 8313 9873 8347
rect 9907 8344 9919 8347
rect 9907 8316 10548 8344
rect 9907 8313 9919 8316
rect 9861 8307 9919 8313
rect 1394 8276 1400 8288
rect 1355 8248 1400 8276
rect 1394 8236 1400 8248
rect 1452 8236 1458 8288
rect 3970 8236 3976 8288
rect 4028 8276 4034 8288
rect 5626 8276 5632 8288
rect 4028 8248 5632 8276
rect 4028 8236 4034 8248
rect 5626 8236 5632 8248
rect 5684 8236 5690 8288
rect 6089 8279 6147 8285
rect 6089 8245 6101 8279
rect 6135 8276 6147 8279
rect 6362 8276 6368 8288
rect 6135 8248 6368 8276
rect 6135 8245 6147 8248
rect 6089 8239 6147 8245
rect 6362 8236 6368 8248
rect 6420 8236 6426 8288
rect 6546 8236 6552 8288
rect 6604 8276 6610 8288
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 6604 8248 8217 8276
rect 6604 8236 6610 8248
rect 8205 8245 8217 8248
rect 8251 8245 8263 8279
rect 8478 8276 8484 8288
rect 8439 8248 8484 8276
rect 8205 8239 8263 8245
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 8662 8236 8668 8288
rect 8720 8276 8726 8288
rect 8846 8276 8852 8288
rect 8720 8248 8852 8276
rect 8720 8236 8726 8248
rect 8846 8236 8852 8248
rect 8904 8236 8910 8288
rect 8941 8279 8999 8285
rect 8941 8245 8953 8279
rect 8987 8276 8999 8279
rect 9493 8279 9551 8285
rect 9493 8276 9505 8279
rect 8987 8248 9505 8276
rect 8987 8245 8999 8248
rect 8941 8239 8999 8245
rect 9493 8245 9505 8248
rect 9539 8245 9551 8279
rect 9950 8276 9956 8288
rect 9911 8248 9956 8276
rect 9493 8239 9551 8245
rect 9950 8236 9956 8248
rect 10008 8236 10014 8288
rect 10520 8285 10548 8316
rect 10686 8304 10692 8356
rect 10744 8344 10750 8356
rect 10873 8347 10931 8353
rect 10873 8344 10885 8347
rect 10744 8316 10885 8344
rect 10744 8304 10750 8316
rect 10873 8313 10885 8316
rect 10919 8344 10931 8347
rect 14829 8347 14887 8353
rect 10919 8316 12112 8344
rect 10919 8313 10931 8316
rect 10873 8307 10931 8313
rect 10505 8279 10563 8285
rect 10505 8245 10517 8279
rect 10551 8245 10563 8279
rect 10505 8239 10563 8245
rect 10965 8279 11023 8285
rect 10965 8245 10977 8279
rect 11011 8276 11023 8279
rect 11974 8276 11980 8288
rect 11011 8248 11980 8276
rect 11011 8245 11023 8248
rect 10965 8239 11023 8245
rect 11974 8236 11980 8248
rect 12032 8236 12038 8288
rect 12084 8276 12112 8316
rect 14829 8313 14841 8347
rect 14875 8344 14887 8347
rect 16206 8344 16212 8356
rect 14875 8316 16212 8344
rect 14875 8313 14887 8316
rect 14829 8307 14887 8313
rect 16206 8304 16212 8316
rect 16264 8304 16270 8356
rect 16316 8344 16344 8384
rect 16384 8381 16396 8415
rect 16430 8412 16442 8415
rect 16850 8412 16856 8424
rect 16430 8384 16856 8412
rect 16430 8381 16442 8384
rect 16384 8375 16442 8381
rect 16850 8372 16856 8384
rect 16908 8372 16914 8424
rect 18509 8415 18567 8421
rect 18509 8381 18521 8415
rect 18555 8412 18567 8415
rect 18690 8412 18696 8424
rect 18555 8384 18696 8412
rect 18555 8381 18567 8384
rect 18509 8375 18567 8381
rect 18690 8372 18696 8384
rect 18748 8372 18754 8424
rect 19150 8372 19156 8424
rect 19208 8412 19214 8424
rect 20441 8415 20499 8421
rect 20441 8412 20453 8415
rect 19208 8384 20453 8412
rect 19208 8372 19214 8384
rect 20441 8381 20453 8384
rect 20487 8381 20499 8415
rect 20441 8375 20499 8381
rect 20533 8415 20591 8421
rect 20533 8381 20545 8415
rect 20579 8412 20591 8415
rect 20714 8412 20720 8424
rect 20579 8384 20720 8412
rect 20579 8381 20591 8384
rect 20533 8375 20591 8381
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 19429 8347 19487 8353
rect 19429 8344 19441 8347
rect 16316 8316 19441 8344
rect 19429 8313 19441 8316
rect 19475 8313 19487 8347
rect 20254 8344 20260 8356
rect 19429 8307 19487 8313
rect 19536 8316 20260 8344
rect 13817 8279 13875 8285
rect 13817 8276 13829 8279
rect 12084 8248 13829 8276
rect 13817 8245 13829 8248
rect 13863 8245 13875 8279
rect 13817 8239 13875 8245
rect 14458 8236 14464 8288
rect 14516 8276 14522 8288
rect 15194 8276 15200 8288
rect 14516 8248 15200 8276
rect 14516 8236 14522 8248
rect 15194 8236 15200 8248
rect 15252 8236 15258 8288
rect 15749 8279 15807 8285
rect 15749 8245 15761 8279
rect 15795 8276 15807 8279
rect 15838 8276 15844 8288
rect 15795 8248 15844 8276
rect 15795 8245 15807 8248
rect 15749 8239 15807 8245
rect 15838 8236 15844 8248
rect 15896 8236 15902 8288
rect 16390 8236 16396 8288
rect 16448 8276 16454 8288
rect 17586 8276 17592 8288
rect 16448 8248 17592 8276
rect 16448 8236 16454 8248
rect 17586 8236 17592 8248
rect 17644 8236 17650 8288
rect 18417 8279 18475 8285
rect 18417 8245 18429 8279
rect 18463 8276 18475 8279
rect 19536 8276 19564 8316
rect 20254 8304 20260 8316
rect 20312 8304 20318 8356
rect 21358 8276 21364 8288
rect 18463 8248 21364 8276
rect 18463 8245 18475 8248
rect 18417 8239 18475 8245
rect 21358 8236 21364 8248
rect 21416 8236 21422 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 2133 8075 2191 8081
rect 2133 8041 2145 8075
rect 2179 8072 2191 8075
rect 3970 8072 3976 8084
rect 2179 8044 3976 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 3970 8032 3976 8044
rect 4028 8032 4034 8084
rect 4065 8075 4123 8081
rect 4065 8041 4077 8075
rect 4111 8041 4123 8075
rect 4065 8035 4123 8041
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 4571 8044 5089 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 5077 8041 5089 8044
rect 5123 8041 5135 8075
rect 5077 8035 5135 8041
rect 5537 8075 5595 8081
rect 5537 8041 5549 8075
rect 5583 8072 5595 8075
rect 5994 8072 6000 8084
rect 5583 8044 6000 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 4080 8004 4108 8035
rect 5994 8032 6000 8044
rect 6052 8032 6058 8084
rect 6089 8075 6147 8081
rect 6089 8041 6101 8075
rect 6135 8072 6147 8075
rect 6178 8072 6184 8084
rect 6135 8044 6184 8072
rect 6135 8041 6147 8044
rect 6089 8035 6147 8041
rect 6178 8032 6184 8044
rect 6236 8032 6242 8084
rect 6454 8032 6460 8084
rect 6512 8072 6518 8084
rect 6549 8075 6607 8081
rect 6549 8072 6561 8075
rect 6512 8044 6561 8072
rect 6512 8032 6518 8044
rect 6549 8041 6561 8044
rect 6595 8041 6607 8075
rect 6549 8035 6607 8041
rect 6917 8075 6975 8081
rect 6917 8041 6929 8075
rect 6963 8072 6975 8075
rect 8294 8072 8300 8084
rect 6963 8044 8300 8072
rect 6963 8041 6975 8044
rect 6917 8035 6975 8041
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 8496 8044 8892 8072
rect 4893 8007 4951 8013
rect 4893 8004 4905 8007
rect 1596 7976 4108 8004
rect 4172 7976 4905 8004
rect 1596 7945 1624 7976
rect 2590 7945 2596 7948
rect 1581 7939 1639 7945
rect 1581 7905 1593 7939
rect 1627 7905 1639 7939
rect 1581 7899 1639 7905
rect 1857 7939 1915 7945
rect 1857 7905 1869 7939
rect 1903 7936 1915 7939
rect 2133 7939 2191 7945
rect 2133 7936 2145 7939
rect 1903 7908 2145 7936
rect 1903 7905 1915 7908
rect 1857 7899 1915 7905
rect 2133 7905 2145 7908
rect 2179 7905 2191 7939
rect 2584 7936 2596 7945
rect 2503 7908 2596 7936
rect 2133 7899 2191 7905
rect 2584 7899 2596 7908
rect 2648 7936 2654 7948
rect 4172 7936 4200 7976
rect 4893 7973 4905 7976
rect 4939 7973 4951 8007
rect 7285 8007 7343 8013
rect 4893 7967 4951 7973
rect 5276 7976 7236 8004
rect 2648 7908 4200 7936
rect 2590 7896 2596 7899
rect 2648 7896 2654 7908
rect 4246 7896 4252 7948
rect 4304 7936 4310 7948
rect 4433 7939 4491 7945
rect 4433 7936 4445 7939
rect 4304 7908 4445 7936
rect 4304 7896 4310 7908
rect 4433 7905 4445 7908
rect 4479 7905 4491 7939
rect 5276 7936 5304 7976
rect 5442 7936 5448 7948
rect 4433 7899 4491 7905
rect 4540 7908 5304 7936
rect 5403 7908 5448 7936
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 1762 7692 1768 7744
rect 1820 7732 1826 7744
rect 2332 7732 2360 7831
rect 3970 7828 3976 7880
rect 4028 7868 4034 7880
rect 4540 7868 4568 7908
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 6270 7936 6276 7948
rect 6231 7908 6276 7936
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 6365 7939 6423 7945
rect 6365 7905 6377 7939
rect 6411 7905 6423 7939
rect 7208 7936 7236 7976
rect 7285 7973 7297 8007
rect 7331 8004 7343 8007
rect 8496 8004 8524 8044
rect 7331 7976 8524 8004
rect 8864 8004 8892 8044
rect 9122 8032 9128 8084
rect 9180 8072 9186 8084
rect 9309 8075 9367 8081
rect 9309 8072 9321 8075
rect 9180 8044 9321 8072
rect 9180 8032 9186 8044
rect 9309 8041 9321 8044
rect 9355 8041 9367 8075
rect 9309 8035 9367 8041
rect 9401 8075 9459 8081
rect 9401 8041 9413 8075
rect 9447 8072 9459 8075
rect 9950 8072 9956 8084
rect 9447 8044 9956 8072
rect 9447 8041 9459 8044
rect 9401 8035 9459 8041
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 10100 8044 12296 8072
rect 10100 8032 10106 8044
rect 9674 8004 9680 8016
rect 8864 7976 9680 8004
rect 7331 7973 7343 7976
rect 7285 7967 7343 7973
rect 9674 7964 9680 7976
rect 9732 7964 9738 8016
rect 10318 8004 10324 8016
rect 9784 7976 10324 8004
rect 7466 7936 7472 7948
rect 7208 7908 7472 7936
rect 6365 7899 6423 7905
rect 4028 7840 4568 7868
rect 4617 7871 4675 7877
rect 4028 7828 4034 7840
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7868 4951 7871
rect 5629 7871 5687 7877
rect 5629 7868 5641 7871
rect 4939 7840 5641 7868
rect 4939 7837 4951 7840
rect 4893 7831 4951 7837
rect 5629 7837 5641 7840
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 3697 7803 3755 7809
rect 3697 7769 3709 7803
rect 3743 7800 3755 7803
rect 4338 7800 4344 7812
rect 3743 7772 4344 7800
rect 3743 7769 3755 7772
rect 3697 7763 3755 7769
rect 4338 7760 4344 7772
rect 4396 7800 4402 7812
rect 4632 7800 4660 7831
rect 4396 7772 4660 7800
rect 4396 7760 4402 7772
rect 4798 7760 4804 7812
rect 4856 7800 4862 7812
rect 6380 7800 6408 7899
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 7650 7896 7656 7948
rect 7708 7936 7714 7948
rect 7834 7936 7840 7948
rect 7708 7908 7840 7936
rect 7708 7896 7714 7908
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 8202 7945 8208 7948
rect 8196 7936 8208 7945
rect 8115 7908 8208 7936
rect 8196 7899 8208 7908
rect 8260 7936 8266 7948
rect 9784 7936 9812 7976
rect 10318 7964 10324 7976
rect 10376 8004 10382 8016
rect 10864 8007 10922 8013
rect 10376 7976 10723 8004
rect 10376 7964 10382 7976
rect 9950 7936 9956 7948
rect 8260 7908 9812 7936
rect 9911 7908 9956 7936
rect 8202 7896 8208 7899
rect 8260 7896 8266 7908
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 10594 7936 10600 7948
rect 10555 7908 10600 7936
rect 10594 7896 10600 7908
rect 10652 7896 10658 7948
rect 10695 7936 10723 7976
rect 10864 7973 10876 8007
rect 10910 8004 10922 8007
rect 12158 8004 12164 8016
rect 10910 7976 12164 8004
rect 10910 7973 10922 7976
rect 10864 7967 10922 7973
rect 12158 7964 12164 7976
rect 12216 7964 12222 8016
rect 12268 8004 12296 8044
rect 12342 8032 12348 8084
rect 12400 8072 12406 8084
rect 12713 8075 12771 8081
rect 12713 8072 12725 8075
rect 12400 8044 12725 8072
rect 12400 8032 12406 8044
rect 12713 8041 12725 8044
rect 12759 8041 12771 8075
rect 13814 8072 13820 8084
rect 12713 8035 12771 8041
rect 12995 8044 13820 8072
rect 12621 8007 12679 8013
rect 12621 8004 12633 8007
rect 12268 7976 12633 8004
rect 12621 7973 12633 7976
rect 12667 8004 12679 8007
rect 12995 8004 13023 8044
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 14366 8032 14372 8084
rect 14424 8072 14430 8084
rect 15010 8072 15016 8084
rect 14424 8044 15016 8072
rect 14424 8032 14430 8044
rect 15010 8032 15016 8044
rect 15068 8032 15074 8084
rect 15286 8072 15292 8084
rect 15247 8044 15292 8072
rect 15286 8032 15292 8044
rect 15344 8032 15350 8084
rect 15654 8032 15660 8084
rect 15712 8072 15718 8084
rect 15749 8075 15807 8081
rect 15749 8072 15761 8075
rect 15712 8044 15761 8072
rect 15712 8032 15718 8044
rect 15749 8041 15761 8044
rect 15795 8041 15807 8075
rect 15749 8035 15807 8041
rect 16669 8075 16727 8081
rect 16669 8041 16681 8075
rect 16715 8072 16727 8075
rect 17678 8072 17684 8084
rect 16715 8044 17684 8072
rect 16715 8041 16727 8044
rect 16669 8035 16727 8041
rect 17678 8032 17684 8044
rect 17736 8032 17742 8084
rect 18693 8075 18751 8081
rect 18693 8041 18705 8075
rect 18739 8072 18751 8075
rect 18874 8072 18880 8084
rect 18739 8044 18880 8072
rect 18739 8041 18751 8044
rect 18693 8035 18751 8041
rect 18874 8032 18880 8044
rect 18932 8032 18938 8084
rect 19705 8075 19763 8081
rect 19705 8041 19717 8075
rect 19751 8072 19763 8075
rect 20070 8072 20076 8084
rect 19751 8044 20076 8072
rect 19751 8041 19763 8044
rect 19705 8035 19763 8041
rect 20070 8032 20076 8044
rect 20128 8032 20134 8084
rect 14642 8004 14648 8016
rect 12667 7976 13023 8004
rect 13464 7976 14648 8004
rect 12667 7973 12679 7976
rect 12621 7967 12679 7973
rect 10695 7908 11652 7936
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7837 7435 7871
rect 7377 7831 7435 7837
rect 7561 7871 7619 7877
rect 7561 7837 7573 7871
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 4856 7772 6408 7800
rect 4856 7760 4862 7772
rect 7392 7744 7420 7831
rect 4062 7732 4068 7744
rect 1820 7704 4068 7732
rect 1820 7692 1826 7704
rect 4062 7692 4068 7704
rect 4120 7692 4126 7744
rect 5994 7692 6000 7744
rect 6052 7732 6058 7744
rect 7282 7732 7288 7744
rect 6052 7704 7288 7732
rect 6052 7692 6058 7704
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 7374 7692 7380 7744
rect 7432 7692 7438 7744
rect 7576 7732 7604 7831
rect 7742 7828 7748 7880
rect 7800 7868 7806 7880
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 7800 7840 7941 7868
rect 7800 7828 7806 7840
rect 7929 7837 7941 7840
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 10502 7868 10508 7880
rect 9548 7840 10508 7868
rect 9548 7828 9554 7840
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 11624 7868 11652 7908
rect 11974 7896 11980 7948
rect 12032 7936 12038 7948
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 12032 7908 12081 7936
rect 12032 7896 12038 7908
rect 12069 7905 12081 7908
rect 12115 7905 12127 7939
rect 12069 7899 12127 7905
rect 12434 7896 12440 7948
rect 12492 7936 12498 7948
rect 13464 7945 13492 7976
rect 14642 7964 14648 7976
rect 14700 7964 14706 8016
rect 15102 7964 15108 8016
rect 15160 8004 15166 8016
rect 19061 8007 19119 8013
rect 19061 8004 19073 8007
rect 15160 7976 19073 8004
rect 15160 7964 15166 7976
rect 19061 7973 19073 7976
rect 19107 7973 19119 8007
rect 19061 7967 19119 7973
rect 13449 7939 13507 7945
rect 12492 7908 12931 7936
rect 12492 7896 12498 7908
rect 12805 7871 12863 7877
rect 12805 7868 12817 7871
rect 11624 7840 12817 7868
rect 12805 7837 12817 7840
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 9214 7760 9220 7812
rect 9272 7800 9278 7812
rect 10410 7800 10416 7812
rect 9272 7772 10416 7800
rect 9272 7760 9278 7772
rect 10410 7760 10416 7772
rect 10468 7760 10474 7812
rect 12903 7800 12931 7908
rect 13449 7905 13461 7939
rect 13495 7905 13507 7939
rect 13449 7899 13507 7905
rect 13808 7939 13866 7945
rect 13808 7905 13820 7939
rect 13854 7936 13866 7939
rect 14090 7936 14096 7948
rect 13854 7908 14096 7936
rect 13854 7905 13866 7908
rect 13808 7899 13866 7905
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 15470 7896 15476 7948
rect 15528 7936 15534 7948
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 15528 7908 15669 7936
rect 15528 7896 15534 7908
rect 15657 7905 15669 7908
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 16485 7939 16543 7945
rect 16485 7905 16497 7939
rect 16531 7936 16543 7939
rect 16853 7939 16911 7945
rect 16853 7936 16865 7939
rect 16531 7908 16865 7936
rect 16531 7905 16543 7908
rect 16485 7899 16543 7905
rect 16853 7905 16865 7908
rect 16899 7905 16911 7939
rect 16853 7899 16911 7905
rect 17304 7939 17362 7945
rect 17304 7905 17316 7939
rect 17350 7936 17362 7939
rect 17586 7936 17592 7948
rect 17350 7908 17592 7936
rect 17350 7905 17362 7908
rect 17304 7899 17362 7905
rect 17586 7896 17592 7908
rect 17644 7896 17650 7948
rect 18046 7896 18052 7948
rect 18104 7936 18110 7948
rect 19153 7939 19211 7945
rect 19153 7936 19165 7939
rect 18104 7908 19165 7936
rect 18104 7896 18110 7908
rect 19153 7905 19165 7908
rect 19199 7905 19211 7939
rect 20070 7936 20076 7948
rect 20031 7908 20076 7936
rect 19153 7899 19211 7905
rect 20070 7896 20076 7908
rect 20128 7896 20134 7948
rect 13541 7871 13599 7877
rect 13541 7868 13553 7871
rect 13280 7840 13553 7868
rect 13280 7809 13308 7840
rect 13541 7837 13553 7840
rect 13587 7837 13599 7871
rect 13541 7831 13599 7837
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 15841 7871 15899 7877
rect 15841 7868 15853 7871
rect 15068 7840 15853 7868
rect 15068 7828 15074 7840
rect 15841 7837 15853 7840
rect 15887 7837 15899 7871
rect 15841 7831 15899 7837
rect 16022 7828 16028 7880
rect 16080 7868 16086 7880
rect 17034 7868 17040 7880
rect 16080 7840 17040 7868
rect 16080 7828 16086 7840
rect 17034 7828 17040 7840
rect 17092 7828 17098 7880
rect 19337 7871 19395 7877
rect 19337 7837 19349 7871
rect 19383 7868 19395 7871
rect 19702 7868 19708 7880
rect 19383 7840 19708 7868
rect 19383 7837 19395 7840
rect 19337 7831 19395 7837
rect 19702 7828 19708 7840
rect 19760 7828 19766 7880
rect 20162 7868 20168 7880
rect 20123 7840 20168 7868
rect 20162 7828 20168 7840
rect 20220 7828 20226 7880
rect 20257 7871 20315 7877
rect 20257 7837 20269 7871
rect 20303 7837 20315 7871
rect 20257 7831 20315 7837
rect 13265 7803 13323 7809
rect 13265 7800 13277 7803
rect 11900 7772 12756 7800
rect 12903 7772 13277 7800
rect 9122 7732 9128 7744
rect 7576 7704 9128 7732
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 9306 7692 9312 7744
rect 9364 7732 9370 7744
rect 9401 7735 9459 7741
rect 9401 7732 9413 7735
rect 9364 7704 9413 7732
rect 9364 7692 9370 7704
rect 9401 7701 9413 7704
rect 9447 7701 9459 7735
rect 9401 7695 9459 7701
rect 10137 7735 10195 7741
rect 10137 7701 10149 7735
rect 10183 7732 10195 7735
rect 11900 7732 11928 7772
rect 12728 7744 12756 7772
rect 13265 7769 13277 7772
rect 13311 7769 13323 7803
rect 13265 7763 13323 7769
rect 16853 7803 16911 7809
rect 16853 7769 16865 7803
rect 16899 7800 16911 7803
rect 19058 7800 19064 7812
rect 16899 7772 17080 7800
rect 16899 7769 16911 7772
rect 16853 7763 16911 7769
rect 10183 7704 11928 7732
rect 10183 7701 10195 7704
rect 10137 7695 10195 7701
rect 11974 7692 11980 7744
rect 12032 7732 12038 7744
rect 12161 7735 12219 7741
rect 12032 7704 12077 7732
rect 12032 7692 12038 7704
rect 12161 7701 12173 7735
rect 12207 7732 12219 7735
rect 12253 7735 12311 7741
rect 12253 7732 12265 7735
rect 12207 7704 12265 7732
rect 12207 7701 12219 7704
rect 12161 7695 12219 7701
rect 12253 7701 12265 7704
rect 12299 7701 12311 7735
rect 12253 7695 12311 7701
rect 12710 7692 12716 7744
rect 12768 7692 12774 7744
rect 14182 7692 14188 7744
rect 14240 7732 14246 7744
rect 14918 7732 14924 7744
rect 14240 7704 14924 7732
rect 14240 7692 14246 7704
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 17052 7732 17080 7772
rect 18340 7772 19064 7800
rect 18340 7732 18368 7772
rect 19058 7760 19064 7772
rect 19116 7760 19122 7812
rect 19610 7760 19616 7812
rect 19668 7800 19674 7812
rect 20272 7800 20300 7831
rect 19668 7772 20300 7800
rect 19668 7760 19674 7772
rect 17052 7704 18368 7732
rect 18417 7735 18475 7741
rect 18417 7701 18429 7735
rect 18463 7732 18475 7735
rect 18598 7732 18604 7744
rect 18463 7704 18604 7732
rect 18463 7701 18475 7704
rect 18417 7695 18475 7701
rect 18598 7692 18604 7704
rect 18656 7692 18662 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 2740 7500 3157 7528
rect 2740 7488 2746 7500
rect 3145 7497 3157 7500
rect 3191 7497 3203 7531
rect 4062 7528 4068 7540
rect 3145 7491 3203 7497
rect 3804 7500 4068 7528
rect 1762 7392 1768 7404
rect 1723 7364 1768 7392
rect 1762 7352 1768 7364
rect 1820 7352 1826 7404
rect 3804 7401 3832 7500
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 5442 7528 5448 7540
rect 5403 7500 5448 7528
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 6454 7488 6460 7540
rect 6512 7528 6518 7540
rect 7834 7528 7840 7540
rect 6512 7500 7840 7528
rect 6512 7488 6518 7500
rect 7834 7488 7840 7500
rect 7892 7528 7898 7540
rect 7892 7500 8064 7528
rect 7892 7488 7898 7500
rect 5169 7463 5227 7469
rect 5169 7429 5181 7463
rect 5215 7429 5227 7463
rect 8036 7460 8064 7500
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 8481 7531 8539 7537
rect 8481 7528 8493 7531
rect 8260 7500 8493 7528
rect 8260 7488 8266 7500
rect 8481 7497 8493 7500
rect 8527 7528 8539 7531
rect 8662 7528 8668 7540
rect 8527 7500 8668 7528
rect 8527 7497 8539 7500
rect 8481 7491 8539 7497
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 8849 7531 8907 7537
rect 8849 7497 8861 7531
rect 8895 7528 8907 7531
rect 9214 7528 9220 7540
rect 8895 7500 9220 7528
rect 8895 7497 8907 7500
rect 8849 7491 8907 7497
rect 9214 7488 9220 7500
rect 9272 7488 9278 7540
rect 9490 7488 9496 7540
rect 9548 7488 9554 7540
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 11606 7528 11612 7540
rect 9640 7500 11612 7528
rect 9640 7488 9646 7500
rect 11606 7488 11612 7500
rect 11664 7488 11670 7540
rect 15105 7531 15163 7537
rect 11707 7500 14504 7528
rect 9508 7460 9536 7488
rect 8036 7432 9536 7460
rect 9677 7463 9735 7469
rect 5169 7423 5227 7429
rect 9677 7429 9689 7463
rect 9723 7460 9735 7463
rect 11707 7460 11735 7500
rect 9723 7432 11735 7460
rect 9723 7429 9735 7432
rect 9677 7423 9735 7429
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7361 3847 7395
rect 3789 7355 3847 7361
rect 5074 7352 5080 7404
rect 5132 7392 5138 7404
rect 5184 7392 5212 7423
rect 13722 7420 13728 7472
rect 13780 7460 13786 7472
rect 13817 7463 13875 7469
rect 13817 7460 13829 7463
rect 13780 7432 13829 7460
rect 13780 7420 13786 7432
rect 13817 7429 13829 7432
rect 13863 7429 13875 7463
rect 14090 7460 14096 7472
rect 14051 7432 14096 7460
rect 13817 7423 13875 7429
rect 6086 7392 6092 7404
rect 5132 7364 6092 7392
rect 5132 7352 5138 7364
rect 6086 7352 6092 7364
rect 6144 7352 6150 7404
rect 8202 7352 8208 7404
rect 8260 7352 8266 7404
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 9214 7392 9220 7404
rect 8352 7364 9220 7392
rect 8352 7352 8358 7364
rect 9214 7352 9220 7364
rect 9272 7352 9278 7404
rect 9398 7392 9404 7404
rect 9359 7364 9404 7392
rect 9398 7352 9404 7364
rect 9456 7352 9462 7404
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7392 10379 7395
rect 10410 7392 10416 7404
rect 10367 7364 10416 7392
rect 10367 7361 10379 7364
rect 10321 7355 10379 7361
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 10505 7395 10563 7401
rect 10505 7361 10517 7395
rect 10551 7392 10563 7395
rect 10962 7392 10968 7404
rect 10551 7364 10968 7392
rect 10551 7361 10563 7364
rect 10505 7355 10563 7361
rect 10962 7352 10968 7364
rect 11020 7392 11026 7404
rect 11425 7395 11483 7401
rect 11425 7392 11437 7395
rect 11020 7364 11437 7392
rect 11020 7352 11026 7364
rect 11425 7361 11437 7364
rect 11471 7361 11483 7395
rect 11606 7392 11612 7404
rect 11425 7355 11483 7361
rect 11532 7364 11612 7392
rect 5813 7327 5871 7333
rect 5813 7293 5825 7327
rect 5859 7324 5871 7327
rect 6822 7324 6828 7336
rect 5859 7296 6828 7324
rect 5859 7293 5871 7296
rect 5813 7287 5871 7293
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7324 7159 7327
rect 7190 7324 7196 7336
rect 7147 7296 7196 7324
rect 7147 7293 7159 7296
rect 7101 7287 7159 7293
rect 7190 7284 7196 7296
rect 7248 7324 7254 7336
rect 7742 7324 7748 7336
rect 7248 7296 7748 7324
rect 7248 7284 7254 7296
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 7834 7284 7840 7336
rect 7892 7324 7898 7336
rect 8110 7324 8116 7336
rect 7892 7296 8116 7324
rect 7892 7284 7898 7296
rect 8110 7284 8116 7296
rect 8168 7284 8174 7336
rect 2038 7265 2044 7268
rect 2032 7219 2044 7265
rect 2096 7256 2102 7268
rect 4062 7265 4068 7268
rect 4056 7256 4068 7265
rect 2096 7228 2180 7256
rect 3975 7228 4068 7256
rect 2038 7216 2044 7219
rect 2096 7216 2102 7228
rect 4056 7219 4068 7228
rect 4120 7256 4126 7268
rect 5905 7259 5963 7265
rect 4120 7228 5304 7256
rect 4062 7216 4068 7219
rect 4120 7216 4126 7228
rect 2047 7188 2075 7216
rect 5074 7188 5080 7200
rect 2047 7160 5080 7188
rect 5074 7148 5080 7160
rect 5132 7148 5138 7200
rect 5276 7188 5304 7228
rect 5905 7225 5917 7259
rect 5951 7256 5963 7259
rect 6914 7256 6920 7268
rect 5951 7228 6920 7256
rect 5951 7225 5963 7228
rect 5905 7219 5963 7225
rect 6914 7216 6920 7228
rect 6972 7216 6978 7268
rect 7368 7259 7426 7265
rect 7368 7225 7380 7259
rect 7414 7256 7426 7259
rect 8220 7256 8248 7352
rect 8570 7284 8576 7336
rect 8628 7324 8634 7336
rect 10229 7327 10287 7333
rect 10229 7324 10241 7327
rect 8628 7296 10241 7324
rect 8628 7284 8634 7296
rect 10229 7293 10241 7296
rect 10275 7293 10287 7327
rect 10229 7287 10287 7293
rect 11241 7327 11299 7333
rect 11241 7293 11253 7327
rect 11287 7324 11299 7327
rect 11532 7324 11560 7364
rect 11606 7352 11612 7364
rect 11664 7352 11670 7404
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7392 11943 7395
rect 12066 7392 12072 7404
rect 11931 7364 12072 7392
rect 11931 7361 11943 7364
rect 11885 7355 11943 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 12434 7392 12440 7404
rect 12395 7364 12440 7392
rect 12434 7352 12440 7364
rect 12492 7352 12498 7404
rect 13832 7392 13860 7423
rect 14090 7420 14096 7432
rect 14148 7420 14154 7472
rect 14366 7392 14372 7404
rect 13832 7364 14372 7392
rect 14366 7352 14372 7364
rect 14424 7352 14430 7404
rect 14476 7333 14504 7500
rect 15105 7497 15117 7531
rect 15151 7528 15163 7531
rect 16022 7528 16028 7540
rect 15151 7500 16028 7528
rect 15151 7497 15163 7500
rect 15105 7491 15163 7497
rect 16022 7488 16028 7500
rect 16080 7488 16086 7540
rect 16206 7488 16212 7540
rect 16264 7528 16270 7540
rect 16393 7531 16451 7537
rect 16393 7528 16405 7531
rect 16264 7500 16405 7528
rect 16264 7488 16270 7500
rect 16393 7497 16405 7500
rect 16439 7497 16451 7531
rect 16393 7491 16451 7497
rect 16850 7488 16856 7540
rect 16908 7528 16914 7540
rect 17589 7531 17647 7537
rect 16908 7500 17540 7528
rect 16908 7488 16914 7500
rect 14918 7420 14924 7472
rect 14976 7460 14982 7472
rect 17512 7460 17540 7500
rect 17589 7497 17601 7531
rect 17635 7528 17647 7531
rect 17770 7528 17776 7540
rect 17635 7500 17776 7528
rect 17635 7497 17647 7500
rect 17589 7491 17647 7497
rect 17770 7488 17776 7500
rect 17828 7488 17834 7540
rect 17862 7488 17868 7540
rect 17920 7528 17926 7540
rect 18049 7531 18107 7537
rect 18049 7528 18061 7531
rect 17920 7500 18061 7528
rect 17920 7488 17926 7500
rect 18049 7497 18061 7500
rect 18095 7497 18107 7531
rect 18049 7491 18107 7497
rect 18506 7488 18512 7540
rect 18564 7528 18570 7540
rect 20073 7531 20131 7537
rect 18564 7500 18644 7528
rect 18564 7488 18570 7500
rect 17954 7460 17960 7472
rect 14976 7432 16988 7460
rect 17512 7432 17960 7460
rect 14976 7420 14982 7432
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7392 14795 7395
rect 15194 7392 15200 7404
rect 14783 7364 15200 7392
rect 14783 7361 14795 7364
rect 14737 7355 14795 7361
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 15378 7352 15384 7404
rect 15436 7392 15442 7404
rect 16025 7395 16083 7401
rect 16025 7392 16037 7395
rect 15436 7364 16037 7392
rect 15436 7352 15442 7364
rect 16025 7361 16037 7364
rect 16071 7392 16083 7395
rect 16482 7392 16488 7404
rect 16071 7364 16488 7392
rect 16071 7361 16083 7364
rect 16025 7355 16083 7361
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 16850 7392 16856 7404
rect 16811 7364 16856 7392
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 16960 7401 16988 7432
rect 17954 7420 17960 7432
rect 18012 7420 18018 7472
rect 16945 7395 17003 7401
rect 16945 7361 16957 7395
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 17678 7352 17684 7404
rect 17736 7392 17742 7404
rect 18616 7401 18644 7500
rect 20073 7497 20085 7531
rect 20119 7528 20131 7531
rect 20162 7528 20168 7540
rect 20119 7500 20168 7528
rect 20119 7497 20131 7500
rect 20073 7491 20131 7497
rect 20162 7488 20168 7500
rect 20220 7488 20226 7540
rect 19061 7463 19119 7469
rect 19061 7429 19073 7463
rect 19107 7460 19119 7463
rect 20530 7460 20536 7472
rect 19107 7432 20536 7460
rect 19107 7429 19119 7432
rect 19061 7423 19119 7429
rect 20530 7420 20536 7432
rect 20588 7420 20594 7472
rect 18509 7395 18567 7401
rect 18509 7392 18521 7395
rect 17736 7364 18521 7392
rect 17736 7352 17742 7364
rect 18509 7361 18521 7364
rect 18555 7361 18567 7395
rect 18509 7355 18567 7361
rect 18601 7395 18659 7401
rect 18601 7361 18613 7395
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 18874 7352 18880 7404
rect 18932 7392 18938 7404
rect 19702 7392 19708 7404
rect 18932 7364 19472 7392
rect 19663 7364 19708 7392
rect 18932 7352 18938 7364
rect 14461 7327 14519 7333
rect 11287 7296 11560 7324
rect 11624 7296 14412 7324
rect 11287 7293 11299 7296
rect 11241 7287 11299 7293
rect 9030 7256 9036 7268
rect 7414 7228 8248 7256
rect 8772 7228 9036 7256
rect 7414 7225 7426 7228
rect 7368 7219 7426 7225
rect 5994 7188 6000 7200
rect 5276 7160 6000 7188
rect 5994 7148 6000 7160
rect 6052 7148 6058 7200
rect 6362 7148 6368 7200
rect 6420 7188 6426 7200
rect 8772 7188 8800 7228
rect 9030 7216 9036 7228
rect 9088 7216 9094 7268
rect 9309 7259 9367 7265
rect 9309 7225 9321 7259
rect 9355 7256 9367 7259
rect 9398 7256 9404 7268
rect 9355 7228 9404 7256
rect 9355 7225 9367 7228
rect 9309 7219 9367 7225
rect 9398 7216 9404 7228
rect 9456 7216 9462 7268
rect 9677 7259 9735 7265
rect 9677 7225 9689 7259
rect 9723 7225 9735 7259
rect 9677 7219 9735 7225
rect 6420 7160 8800 7188
rect 6420 7148 6426 7160
rect 8846 7148 8852 7200
rect 8904 7188 8910 7200
rect 9217 7191 9275 7197
rect 9217 7188 9229 7191
rect 8904 7160 9229 7188
rect 8904 7148 8910 7160
rect 9217 7157 9229 7160
rect 9263 7188 9275 7191
rect 9692 7188 9720 7219
rect 10502 7216 10508 7268
rect 10560 7256 10566 7268
rect 10560 7228 10999 7256
rect 10560 7216 10566 7228
rect 9263 7160 9720 7188
rect 9861 7191 9919 7197
rect 9263 7157 9275 7160
rect 9217 7151 9275 7157
rect 9861 7157 9873 7191
rect 9907 7188 9919 7191
rect 10410 7188 10416 7200
rect 9907 7160 10416 7188
rect 9907 7157 9919 7160
rect 9861 7151 9919 7157
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 10870 7188 10876 7200
rect 10831 7160 10876 7188
rect 10870 7148 10876 7160
rect 10928 7148 10934 7200
rect 10971 7188 10999 7228
rect 11054 7216 11060 7268
rect 11112 7256 11118 7268
rect 11333 7259 11391 7265
rect 11333 7256 11345 7259
rect 11112 7228 11345 7256
rect 11112 7216 11118 7228
rect 11333 7225 11345 7228
rect 11379 7225 11391 7259
rect 11333 7219 11391 7225
rect 11422 7216 11428 7268
rect 11480 7256 11486 7268
rect 11624 7256 11652 7296
rect 14384 7268 14412 7296
rect 14461 7293 14473 7327
rect 14507 7293 14519 7327
rect 14461 7287 14519 7293
rect 14642 7284 14648 7336
rect 14700 7324 14706 7336
rect 15289 7327 15347 7333
rect 15289 7324 15301 7327
rect 14700 7296 15301 7324
rect 14700 7284 14706 7296
rect 15289 7293 15301 7296
rect 15335 7293 15347 7327
rect 17405 7327 17463 7333
rect 15289 7287 15347 7293
rect 15396 7296 15976 7324
rect 11480 7228 11652 7256
rect 12704 7259 12762 7265
rect 11480 7216 11486 7228
rect 12704 7225 12716 7259
rect 12750 7256 12762 7259
rect 14182 7256 14188 7268
rect 12750 7228 14188 7256
rect 12750 7225 12762 7228
rect 12704 7219 12762 7225
rect 14182 7216 14188 7228
rect 14240 7216 14246 7268
rect 14366 7216 14372 7268
rect 14424 7216 14430 7268
rect 14550 7256 14556 7268
rect 14511 7228 14556 7256
rect 14550 7216 14556 7228
rect 14608 7216 14614 7268
rect 15102 7216 15108 7268
rect 15160 7256 15166 7268
rect 15396 7256 15424 7296
rect 15160 7228 15424 7256
rect 15160 7216 15166 7228
rect 15470 7216 15476 7268
rect 15528 7256 15534 7268
rect 15841 7259 15899 7265
rect 15841 7256 15853 7259
rect 15528 7228 15853 7256
rect 15528 7216 15534 7228
rect 15841 7225 15853 7228
rect 15887 7225 15899 7259
rect 15948 7256 15976 7296
rect 17405 7293 17417 7327
rect 17451 7324 17463 7327
rect 19334 7324 19340 7336
rect 17451 7296 19340 7324
rect 17451 7293 17463 7296
rect 17405 7287 17463 7293
rect 19334 7284 19340 7296
rect 19392 7284 19398 7336
rect 19444 7333 19472 7364
rect 19702 7352 19708 7364
rect 19760 7352 19766 7404
rect 20625 7395 20683 7401
rect 20625 7361 20637 7395
rect 20671 7361 20683 7395
rect 20625 7355 20683 7361
rect 19429 7327 19487 7333
rect 19429 7293 19441 7327
rect 19475 7293 19487 7327
rect 20640 7324 20668 7355
rect 19429 7287 19487 7293
rect 19628 7296 20668 7324
rect 18417 7259 18475 7265
rect 18417 7256 18429 7259
rect 15948 7228 18429 7256
rect 15841 7219 15899 7225
rect 18417 7225 18429 7228
rect 18463 7225 18475 7259
rect 19521 7259 19579 7265
rect 19521 7256 19533 7259
rect 18417 7219 18475 7225
rect 18524 7228 19533 7256
rect 11440 7188 11468 7216
rect 10971 7160 11468 7188
rect 12158 7148 12164 7200
rect 12216 7188 12222 7200
rect 15286 7188 15292 7200
rect 12216 7160 15292 7188
rect 12216 7148 12222 7160
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 15381 7191 15439 7197
rect 15381 7157 15393 7191
rect 15427 7188 15439 7191
rect 15654 7188 15660 7200
rect 15427 7160 15660 7188
rect 15427 7157 15439 7160
rect 15381 7151 15439 7157
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 15749 7191 15807 7197
rect 15749 7157 15761 7191
rect 15795 7188 15807 7191
rect 16206 7188 16212 7200
rect 15795 7160 16212 7188
rect 15795 7157 15807 7160
rect 15749 7151 15807 7157
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 16574 7148 16580 7200
rect 16632 7188 16638 7200
rect 16761 7191 16819 7197
rect 16761 7188 16773 7191
rect 16632 7160 16773 7188
rect 16632 7148 16638 7160
rect 16761 7157 16773 7160
rect 16807 7157 16819 7191
rect 16761 7151 16819 7157
rect 17218 7148 17224 7200
rect 17276 7188 17282 7200
rect 18524 7188 18552 7228
rect 19521 7225 19533 7228
rect 19567 7225 19579 7259
rect 19521 7219 19579 7225
rect 17276 7160 18552 7188
rect 17276 7148 17282 7160
rect 18690 7148 18696 7200
rect 18748 7188 18754 7200
rect 19628 7188 19656 7296
rect 20533 7259 20591 7265
rect 20533 7225 20545 7259
rect 20579 7256 20591 7259
rect 20622 7256 20628 7268
rect 20579 7228 20628 7256
rect 20579 7225 20591 7228
rect 20533 7219 20591 7225
rect 20622 7216 20628 7228
rect 20680 7216 20686 7268
rect 20438 7188 20444 7200
rect 18748 7160 19656 7188
rect 20399 7160 20444 7188
rect 18748 7148 18754 7160
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 1394 6944 1400 6996
rect 1452 6984 1458 6996
rect 2501 6987 2559 6993
rect 2501 6984 2513 6987
rect 1452 6956 2513 6984
rect 1452 6944 1458 6956
rect 2501 6953 2513 6956
rect 2547 6953 2559 6987
rect 2501 6947 2559 6953
rect 2593 6987 2651 6993
rect 2593 6953 2605 6987
rect 2639 6984 2651 6987
rect 4065 6987 4123 6993
rect 4065 6984 4077 6987
rect 2639 6956 4077 6984
rect 2639 6953 2651 6956
rect 2593 6947 2651 6953
rect 4065 6953 4077 6956
rect 4111 6953 4123 6987
rect 4065 6947 4123 6953
rect 5902 6944 5908 6996
rect 5960 6984 5966 6996
rect 6362 6984 6368 6996
rect 5960 6956 6368 6984
rect 5960 6944 5966 6956
rect 6362 6944 6368 6956
rect 6420 6944 6426 6996
rect 6454 6944 6460 6996
rect 6512 6984 6518 6996
rect 6641 6987 6699 6993
rect 6641 6984 6653 6987
rect 6512 6956 6653 6984
rect 6512 6944 6518 6956
rect 6641 6953 6653 6956
rect 6687 6953 6699 6987
rect 6641 6947 6699 6953
rect 7190 6944 7196 6996
rect 7248 6984 7254 6996
rect 7285 6987 7343 6993
rect 7285 6984 7297 6987
rect 7248 6956 7297 6984
rect 7248 6944 7254 6956
rect 7285 6953 7297 6956
rect 7331 6953 7343 6987
rect 7285 6947 7343 6953
rect 7374 6944 7380 6996
rect 7432 6984 7438 6996
rect 7561 6987 7619 6993
rect 7561 6984 7573 6987
rect 7432 6956 7573 6984
rect 7432 6944 7438 6956
rect 7561 6953 7573 6956
rect 7607 6953 7619 6987
rect 7561 6947 7619 6953
rect 7650 6944 7656 6996
rect 7708 6984 7714 6996
rect 7929 6987 7987 6993
rect 7929 6984 7941 6987
rect 7708 6956 7941 6984
rect 7708 6944 7714 6956
rect 7929 6953 7941 6956
rect 7975 6953 7987 6987
rect 8570 6984 8576 6996
rect 8531 6956 8576 6984
rect 7929 6947 7987 6953
rect 8570 6944 8576 6956
rect 8628 6944 8634 6996
rect 9030 6984 9036 6996
rect 8943 6956 9036 6984
rect 9030 6944 9036 6956
rect 9088 6984 9094 6996
rect 9582 6984 9588 6996
rect 9088 6956 9588 6984
rect 9088 6944 9094 6956
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 9769 6987 9827 6993
rect 9769 6953 9781 6987
rect 9815 6984 9827 6987
rect 10229 6987 10287 6993
rect 10229 6984 10241 6987
rect 9815 6956 10241 6984
rect 9815 6953 9827 6956
rect 9769 6947 9827 6953
rect 10229 6953 10241 6956
rect 10275 6953 10287 6987
rect 10229 6947 10287 6953
rect 10321 6987 10379 6993
rect 10321 6953 10333 6987
rect 10367 6984 10379 6987
rect 10870 6984 10876 6996
rect 10367 6956 10876 6984
rect 10367 6953 10379 6956
rect 10321 6947 10379 6953
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 11238 6984 11244 6996
rect 11151 6956 11244 6984
rect 11238 6944 11244 6956
rect 11296 6984 11302 6996
rect 11793 6987 11851 6993
rect 11296 6956 11744 6984
rect 11296 6944 11302 6956
rect 2958 6876 2964 6928
rect 3016 6916 3022 6928
rect 3602 6916 3608 6928
rect 3016 6888 3608 6916
rect 3016 6876 3022 6888
rect 3602 6876 3608 6888
rect 3660 6916 3666 6928
rect 4433 6919 4491 6925
rect 4433 6916 4445 6919
rect 3660 6888 4445 6916
rect 3660 6876 3666 6888
rect 4433 6885 4445 6888
rect 4479 6885 4491 6919
rect 4433 6879 4491 6885
rect 5445 6919 5503 6925
rect 5445 6885 5457 6919
rect 5491 6916 5503 6919
rect 6178 6916 6184 6928
rect 5491 6888 6184 6916
rect 5491 6885 5503 6888
rect 5445 6879 5503 6885
rect 6178 6876 6184 6888
rect 6236 6876 6242 6928
rect 6270 6876 6276 6928
rect 6328 6916 6334 6928
rect 6328 6888 7512 6916
rect 6328 6876 6334 6888
rect 1581 6851 1639 6857
rect 1581 6817 1593 6851
rect 1627 6848 1639 6851
rect 1762 6848 1768 6860
rect 1627 6820 1768 6848
rect 1627 6817 1639 6820
rect 1581 6811 1639 6817
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 3421 6851 3479 6857
rect 3421 6817 3433 6851
rect 3467 6848 3479 6851
rect 3694 6848 3700 6860
rect 3467 6820 3700 6848
rect 3467 6817 3479 6820
rect 3421 6811 3479 6817
rect 3694 6808 3700 6820
rect 3752 6808 3758 6860
rect 4525 6851 4583 6857
rect 4525 6817 4537 6851
rect 4571 6848 4583 6851
rect 5810 6848 5816 6860
rect 4571 6820 5816 6848
rect 4571 6817 4583 6820
rect 4525 6811 4583 6817
rect 5810 6808 5816 6820
rect 5868 6808 5874 6860
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 7484 6857 7512 6888
rect 7742 6876 7748 6928
rect 7800 6916 7806 6928
rect 8110 6916 8116 6928
rect 7800 6888 8116 6916
rect 7800 6876 7806 6888
rect 8110 6876 8116 6888
rect 8168 6876 8174 6928
rect 8662 6916 8668 6928
rect 8220 6888 8668 6916
rect 7469 6851 7527 6857
rect 6788 6820 6833 6848
rect 6788 6808 6794 6820
rect 7469 6817 7481 6851
rect 7515 6817 7527 6851
rect 7469 6811 7527 6817
rect 2682 6780 2688 6792
rect 2643 6752 2688 6780
rect 2682 6740 2688 6752
rect 2740 6740 2746 6792
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6780 3387 6783
rect 4246 6780 4252 6792
rect 3375 6752 4252 6780
rect 3375 6749 3387 6752
rect 3329 6743 3387 6749
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6780 4767 6783
rect 5074 6780 5080 6792
rect 4755 6752 5080 6780
rect 4755 6749 4767 6752
rect 4709 6743 4767 6749
rect 5074 6740 5080 6752
rect 5132 6740 5138 6792
rect 5534 6780 5540 6792
rect 5495 6752 5540 6780
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 5721 6783 5779 6789
rect 5721 6749 5733 6783
rect 5767 6780 5779 6783
rect 5902 6780 5908 6792
rect 5767 6752 5908 6780
rect 5767 6749 5779 6752
rect 5721 6743 5779 6749
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6780 6239 6783
rect 6748 6780 6776 6808
rect 6227 6752 6776 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 6822 6740 6828 6792
rect 6880 6780 6886 6792
rect 6880 6752 6925 6780
rect 6880 6740 6886 6752
rect 7558 6740 7564 6792
rect 7616 6780 7622 6792
rect 8018 6780 8024 6792
rect 7616 6752 8024 6780
rect 7616 6740 7622 6752
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 8220 6789 8248 6888
rect 8662 6876 8668 6888
rect 8720 6876 8726 6928
rect 8941 6919 8999 6925
rect 8941 6885 8953 6919
rect 8987 6916 8999 6919
rect 11514 6916 11520 6928
rect 8987 6888 11520 6916
rect 8987 6885 8999 6888
rect 8941 6879 8999 6885
rect 11514 6876 11520 6888
rect 11572 6876 11578 6928
rect 11716 6916 11744 6956
rect 11793 6953 11805 6987
rect 11839 6984 11851 6987
rect 11885 6987 11943 6993
rect 11885 6984 11897 6987
rect 11839 6956 11897 6984
rect 11839 6953 11851 6956
rect 11793 6947 11851 6953
rect 11885 6953 11897 6956
rect 11931 6953 11943 6987
rect 12158 6984 12164 6996
rect 11885 6947 11943 6953
rect 11992 6956 12164 6984
rect 11992 6916 12020 6956
rect 12158 6944 12164 6956
rect 12216 6944 12222 6996
rect 12345 6987 12403 6993
rect 12345 6953 12357 6987
rect 12391 6984 12403 6987
rect 12802 6984 12808 6996
rect 12391 6956 12808 6984
rect 12391 6953 12403 6956
rect 12345 6947 12403 6953
rect 12802 6944 12808 6956
rect 12860 6944 12866 6996
rect 13170 6944 13176 6996
rect 13228 6984 13234 6996
rect 15470 6984 15476 6996
rect 13228 6956 15476 6984
rect 13228 6944 13234 6956
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 15654 6984 15660 6996
rect 15615 6956 15660 6984
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 16850 6944 16856 6996
rect 16908 6984 16914 6996
rect 17034 6984 17040 6996
rect 16908 6956 17040 6984
rect 16908 6944 16914 6956
rect 17034 6944 17040 6956
rect 17092 6984 17098 6996
rect 17862 6984 17868 6996
rect 17092 6956 17724 6984
rect 17823 6956 17868 6984
rect 17092 6944 17098 6956
rect 11716 6888 12020 6916
rect 12066 6876 12072 6928
rect 12124 6916 12130 6928
rect 12253 6919 12311 6925
rect 12253 6916 12265 6919
rect 12124 6888 12265 6916
rect 12124 6876 12130 6888
rect 12253 6885 12265 6888
rect 12299 6885 12311 6919
rect 12894 6916 12900 6928
rect 12253 6879 12311 6885
rect 12452 6888 12900 6916
rect 9490 6848 9496 6860
rect 9232 6820 9496 6848
rect 9232 6789 9260 6820
rect 9490 6808 9496 6820
rect 9548 6848 9554 6860
rect 9548 6820 11560 6848
rect 9548 6808 9554 6820
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 9582 6740 9588 6792
rect 9640 6780 9646 6792
rect 9769 6783 9827 6789
rect 9769 6780 9781 6783
rect 9640 6752 9781 6780
rect 9640 6740 9646 6752
rect 9769 6749 9781 6752
rect 9815 6749 9827 6783
rect 10410 6780 10416 6792
rect 10371 6752 10416 6780
rect 9769 6743 9827 6749
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 11333 6783 11391 6789
rect 10520 6752 11192 6780
rect 1762 6712 1768 6724
rect 1723 6684 1768 6712
rect 1762 6672 1768 6684
rect 1820 6672 1826 6724
rect 10520 6712 10548 6752
rect 4163 6684 10548 6712
rect 10873 6715 10931 6721
rect 2133 6647 2191 6653
rect 2133 6613 2145 6647
rect 2179 6644 2191 6647
rect 3329 6647 3387 6653
rect 3329 6644 3341 6647
rect 2179 6616 3341 6644
rect 2179 6613 2191 6616
rect 2133 6607 2191 6613
rect 3329 6613 3341 6616
rect 3375 6613 3387 6647
rect 3602 6644 3608 6656
rect 3563 6616 3608 6644
rect 3329 6607 3387 6613
rect 3602 6604 3608 6616
rect 3660 6604 3666 6656
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 4163 6644 4191 6684
rect 10873 6681 10885 6715
rect 10919 6712 10931 6715
rect 11054 6712 11060 6724
rect 10919 6684 11060 6712
rect 10919 6681 10931 6684
rect 10873 6675 10931 6681
rect 11054 6672 11060 6684
rect 11112 6672 11118 6724
rect 11164 6712 11192 6752
rect 11333 6749 11345 6783
rect 11379 6780 11391 6783
rect 11422 6780 11428 6792
rect 11379 6752 11428 6780
rect 11379 6749 11391 6752
rect 11333 6743 11391 6749
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 11532 6789 11560 6820
rect 11606 6808 11612 6860
rect 11664 6848 11670 6860
rect 11793 6851 11851 6857
rect 11793 6848 11805 6851
rect 11664 6820 11805 6848
rect 11664 6808 11670 6820
rect 11793 6817 11805 6820
rect 11839 6817 11851 6851
rect 11793 6811 11851 6817
rect 11882 6808 11888 6860
rect 11940 6848 11946 6860
rect 12452 6848 12480 6888
rect 12894 6876 12900 6888
rect 12952 6876 12958 6928
rect 13078 6876 13084 6928
rect 13136 6916 13142 6928
rect 13265 6919 13323 6925
rect 13265 6916 13277 6919
rect 13136 6888 13277 6916
rect 13136 6876 13142 6888
rect 13265 6885 13277 6888
rect 13311 6916 13323 6919
rect 14182 6916 14188 6928
rect 13311 6888 14188 6916
rect 13311 6885 13323 6888
rect 13265 6879 13323 6885
rect 14182 6876 14188 6888
rect 14240 6876 14246 6928
rect 14366 6876 14372 6928
rect 14424 6916 14430 6928
rect 14553 6919 14611 6925
rect 14553 6916 14565 6919
rect 14424 6888 14565 6916
rect 14424 6876 14430 6888
rect 14553 6885 14565 6888
rect 14599 6916 14611 6919
rect 15102 6916 15108 6928
rect 14599 6888 15108 6916
rect 14599 6885 14611 6888
rect 14553 6879 14611 6885
rect 15102 6876 15108 6888
rect 15160 6876 15166 6928
rect 15746 6876 15752 6928
rect 15804 6916 15810 6928
rect 17218 6916 17224 6928
rect 15804 6888 16344 6916
rect 17179 6888 17224 6916
rect 15804 6876 15810 6888
rect 11940 6820 12480 6848
rect 11940 6808 11946 6820
rect 12526 6808 12532 6860
rect 12584 6848 12590 6860
rect 13906 6848 13912 6860
rect 12584 6820 13912 6848
rect 12584 6808 12590 6820
rect 13906 6808 13912 6820
rect 13964 6808 13970 6860
rect 16316 6857 16344 6888
rect 17218 6876 17224 6888
rect 17276 6876 17282 6928
rect 17696 6916 17724 6956
rect 17862 6944 17868 6956
rect 17920 6944 17926 6996
rect 18230 6984 18236 6996
rect 18191 6956 18236 6984
rect 18230 6944 18236 6956
rect 18288 6944 18294 6996
rect 18322 6944 18328 6996
rect 18380 6984 18386 6996
rect 18380 6956 18425 6984
rect 18380 6944 18386 6956
rect 18506 6944 18512 6996
rect 18564 6984 18570 6996
rect 18690 6984 18696 6996
rect 18564 6956 18696 6984
rect 18564 6944 18570 6956
rect 18690 6944 18696 6956
rect 18748 6944 18754 6996
rect 18782 6944 18788 6996
rect 18840 6984 18846 6996
rect 19334 6984 19340 6996
rect 18840 6956 19340 6984
rect 18840 6944 18846 6956
rect 19334 6944 19340 6956
rect 19392 6944 19398 6996
rect 19061 6919 19119 6925
rect 19061 6916 19073 6919
rect 17696 6888 19073 6916
rect 19061 6885 19073 6888
rect 19107 6885 19119 6919
rect 19518 6916 19524 6928
rect 19061 6879 19119 6885
rect 19159 6888 19524 6916
rect 14645 6851 14703 6857
rect 14645 6817 14657 6851
rect 14691 6848 14703 6851
rect 16301 6851 16359 6857
rect 14691 6820 16160 6848
rect 14691 6817 14703 6820
rect 14645 6811 14703 6817
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6780 11575 6783
rect 11974 6780 11980 6792
rect 11563 6752 11980 6780
rect 11563 6749 11575 6752
rect 11517 6743 11575 6749
rect 11974 6740 11980 6752
rect 12032 6780 12038 6792
rect 12437 6783 12495 6789
rect 12437 6780 12449 6783
rect 12032 6752 12449 6780
rect 12032 6740 12038 6752
rect 12437 6749 12449 6752
rect 12483 6749 12495 6783
rect 12437 6743 12495 6749
rect 13170 6740 13176 6792
rect 13228 6780 13234 6792
rect 13357 6783 13415 6789
rect 13357 6780 13369 6783
rect 13228 6752 13369 6780
rect 13228 6740 13234 6752
rect 13357 6749 13369 6752
rect 13403 6749 13415 6783
rect 13538 6780 13544 6792
rect 13499 6752 13544 6780
rect 13357 6743 13415 6749
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 14090 6780 14096 6792
rect 14003 6752 14096 6780
rect 14090 6740 14096 6752
rect 14148 6780 14154 6792
rect 14660 6780 14688 6811
rect 14148 6752 14688 6780
rect 14829 6783 14887 6789
rect 14148 6740 14154 6752
rect 14829 6749 14841 6783
rect 14875 6780 14887 6783
rect 15378 6780 15384 6792
rect 14875 6752 15384 6780
rect 14875 6749 14887 6752
rect 14829 6743 14887 6749
rect 15378 6740 15384 6752
rect 15436 6740 15442 6792
rect 15749 6783 15807 6789
rect 15749 6749 15761 6783
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 15933 6783 15991 6789
rect 15933 6749 15945 6783
rect 15979 6780 15991 6783
rect 16022 6780 16028 6792
rect 15979 6752 16028 6780
rect 15979 6749 15991 6752
rect 15933 6743 15991 6749
rect 14185 6715 14243 6721
rect 11164 6684 14136 6712
rect 4028 6616 4191 6644
rect 5077 6647 5135 6653
rect 4028 6604 4034 6616
rect 5077 6613 5089 6647
rect 5123 6644 5135 6647
rect 5994 6644 6000 6656
rect 5123 6616 6000 6644
rect 5123 6613 5135 6616
rect 5077 6607 5135 6613
rect 5994 6604 6000 6616
rect 6052 6604 6058 6656
rect 6270 6644 6276 6656
rect 6231 6616 6276 6644
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 8018 6604 8024 6656
rect 8076 6644 8082 6656
rect 9214 6644 9220 6656
rect 8076 6616 9220 6644
rect 8076 6604 8082 6616
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 9766 6644 9772 6656
rect 9364 6616 9772 6644
rect 9364 6604 9370 6616
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 9861 6647 9919 6653
rect 9861 6613 9873 6647
rect 9907 6644 9919 6647
rect 10686 6644 10692 6656
rect 9907 6616 10692 6644
rect 9907 6613 9919 6616
rect 9861 6607 9919 6613
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 12897 6647 12955 6653
rect 12897 6644 12909 6647
rect 11664 6616 12909 6644
rect 11664 6604 11670 6616
rect 12897 6613 12909 6616
rect 12943 6613 12955 6647
rect 12897 6607 12955 6613
rect 13354 6604 13360 6656
rect 13412 6644 13418 6656
rect 13538 6644 13544 6656
rect 13412 6616 13544 6644
rect 13412 6604 13418 6616
rect 13538 6604 13544 6616
rect 13596 6604 13602 6656
rect 14108 6644 14136 6684
rect 14185 6681 14197 6715
rect 14231 6712 14243 6715
rect 15764 6712 15792 6743
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 16132 6780 16160 6820
rect 16301 6817 16313 6851
rect 16347 6817 16359 6851
rect 17678 6848 17684 6860
rect 16301 6811 16359 6817
rect 16408 6820 17684 6848
rect 16408 6780 16436 6820
rect 17678 6808 17684 6820
rect 17736 6808 17742 6860
rect 19159 6848 19187 6888
rect 19518 6876 19524 6888
rect 19576 6876 19582 6928
rect 18432 6820 19187 6848
rect 16132 6752 16436 6780
rect 17313 6783 17371 6789
rect 17313 6749 17325 6783
rect 17359 6749 17371 6783
rect 17313 6743 17371 6749
rect 17497 6783 17555 6789
rect 17497 6749 17509 6783
rect 17543 6749 17555 6783
rect 17497 6743 17555 6749
rect 17328 6712 17356 6743
rect 14231 6684 15792 6712
rect 16316 6684 17356 6712
rect 17512 6712 17540 6743
rect 18322 6740 18328 6792
rect 18380 6780 18386 6792
rect 18432 6789 18460 6820
rect 19242 6808 19248 6860
rect 19300 6848 19306 6860
rect 19409 6851 19467 6857
rect 19409 6848 19421 6851
rect 19300 6820 19421 6848
rect 19300 6808 19306 6820
rect 19409 6817 19421 6820
rect 19455 6817 19467 6851
rect 19409 6811 19467 6817
rect 20901 6851 20959 6857
rect 20901 6817 20913 6851
rect 20947 6848 20959 6851
rect 21082 6848 21088 6860
rect 20947 6820 21088 6848
rect 20947 6817 20959 6820
rect 20901 6811 20959 6817
rect 21082 6808 21088 6820
rect 21140 6808 21146 6860
rect 18417 6783 18475 6789
rect 18417 6780 18429 6783
rect 18380 6752 18429 6780
rect 18380 6740 18386 6752
rect 18417 6749 18429 6752
rect 18463 6749 18475 6783
rect 18417 6743 18475 6749
rect 19061 6783 19119 6789
rect 19061 6749 19073 6783
rect 19107 6780 19119 6783
rect 19150 6780 19156 6792
rect 19107 6752 19156 6780
rect 19107 6749 19119 6752
rect 19061 6743 19119 6749
rect 19150 6740 19156 6752
rect 19208 6740 19214 6792
rect 17678 6712 17684 6724
rect 17512 6684 17684 6712
rect 14231 6681 14243 6684
rect 14185 6675 14243 6681
rect 15102 6644 15108 6656
rect 14108 6616 15108 6644
rect 15102 6604 15108 6616
rect 15160 6604 15166 6656
rect 15289 6647 15347 6653
rect 15289 6613 15301 6647
rect 15335 6644 15347 6647
rect 16316 6644 16344 6684
rect 17678 6672 17684 6684
rect 17736 6672 17742 6724
rect 15335 6616 16344 6644
rect 16485 6647 16543 6653
rect 15335 6613 15347 6616
rect 15289 6607 15347 6613
rect 16485 6613 16497 6647
rect 16531 6644 16543 6647
rect 16758 6644 16764 6656
rect 16531 6616 16764 6644
rect 16531 6613 16543 6616
rect 16485 6607 16543 6613
rect 16758 6604 16764 6616
rect 16816 6604 16822 6656
rect 16853 6647 16911 6653
rect 16853 6613 16865 6647
rect 16899 6644 16911 6647
rect 17402 6644 17408 6656
rect 16899 6616 17408 6644
rect 16899 6613 16911 6616
rect 16853 6607 16911 6613
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 17586 6604 17592 6656
rect 17644 6644 17650 6656
rect 20254 6644 20260 6656
rect 17644 6616 20260 6644
rect 17644 6604 17650 6616
rect 20254 6604 20260 6616
rect 20312 6644 20318 6656
rect 20533 6647 20591 6653
rect 20533 6644 20545 6647
rect 20312 6616 20545 6644
rect 20312 6604 20318 6616
rect 20533 6613 20545 6616
rect 20579 6613 20591 6647
rect 20533 6607 20591 6613
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 2130 6400 2136 6452
rect 2188 6440 2194 6452
rect 2869 6443 2927 6449
rect 2869 6440 2881 6443
rect 2188 6412 2881 6440
rect 2188 6400 2194 6412
rect 2869 6409 2881 6412
rect 2915 6409 2927 6443
rect 2869 6403 2927 6409
rect 4246 6400 4252 6452
rect 4304 6440 4310 6452
rect 13262 6440 13268 6452
rect 4304 6412 13268 6440
rect 4304 6400 4310 6412
rect 13262 6400 13268 6412
rect 13320 6400 13326 6452
rect 13354 6400 13360 6452
rect 13412 6440 13418 6452
rect 13998 6440 14004 6452
rect 13412 6412 13676 6440
rect 13959 6412 14004 6440
rect 13412 6400 13418 6412
rect 1762 6332 1768 6384
rect 1820 6372 1826 6384
rect 2314 6372 2320 6384
rect 1820 6344 2320 6372
rect 1820 6332 1826 6344
rect 2314 6332 2320 6344
rect 2372 6332 2378 6384
rect 3602 6332 3608 6384
rect 3660 6372 3666 6384
rect 4062 6372 4068 6384
rect 3660 6344 4068 6372
rect 3660 6332 3666 6344
rect 4062 6332 4068 6344
rect 4120 6332 4126 6384
rect 4985 6375 5043 6381
rect 4985 6341 4997 6375
rect 5031 6372 5043 6375
rect 5077 6375 5135 6381
rect 5077 6372 5089 6375
rect 5031 6344 5089 6372
rect 5031 6341 5043 6344
rect 4985 6335 5043 6341
rect 5077 6341 5089 6344
rect 5123 6341 5135 6375
rect 6270 6372 6276 6384
rect 5077 6335 5135 6341
rect 5552 6344 6276 6372
rect 2222 6264 2228 6316
rect 2280 6304 2286 6316
rect 2501 6307 2559 6313
rect 2501 6304 2513 6307
rect 2280 6276 2513 6304
rect 2280 6264 2286 6276
rect 2501 6273 2513 6276
rect 2547 6273 2559 6307
rect 3510 6304 3516 6316
rect 3471 6276 3516 6304
rect 2501 6267 2559 6273
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 3786 6264 3792 6316
rect 3844 6304 3850 6316
rect 4525 6307 4583 6313
rect 4525 6304 4537 6307
rect 3844 6276 4537 6304
rect 3844 6264 3850 6276
rect 4525 6273 4537 6276
rect 4571 6273 4583 6307
rect 4706 6304 4712 6316
rect 4667 6276 4712 6304
rect 4525 6267 4583 6273
rect 4706 6264 4712 6276
rect 4764 6264 4770 6316
rect 5552 6313 5580 6344
rect 6270 6332 6276 6344
rect 6328 6332 6334 6384
rect 6638 6372 6644 6384
rect 6380 6344 6644 6372
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 5718 6264 5724 6316
rect 5776 6304 5782 6316
rect 6380 6313 6408 6344
rect 6638 6332 6644 6344
rect 6696 6332 6702 6384
rect 7650 6372 7656 6384
rect 7611 6344 7656 6372
rect 7650 6332 7656 6344
rect 7708 6372 7714 6384
rect 8018 6372 8024 6384
rect 7708 6344 8024 6372
rect 7708 6332 7714 6344
rect 8018 6332 8024 6344
rect 8076 6332 8082 6384
rect 8110 6332 8116 6384
rect 8168 6372 8174 6384
rect 8168 6344 8248 6372
rect 8168 6332 8174 6344
rect 6365 6307 6423 6313
rect 5776 6276 5821 6304
rect 5776 6264 5782 6276
rect 6365 6273 6377 6307
rect 6411 6273 6423 6307
rect 6546 6304 6552 6316
rect 6507 6276 6552 6304
rect 6365 6267 6423 6273
rect 6546 6264 6552 6276
rect 6604 6304 6610 6316
rect 6822 6304 6828 6316
rect 6604 6276 6828 6304
rect 6604 6264 6610 6276
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 3973 6239 4031 6245
rect 3973 6205 3985 6239
rect 4019 6236 4031 6239
rect 4433 6239 4491 6245
rect 4433 6236 4445 6239
rect 4019 6208 4445 6236
rect 4019 6205 4031 6208
rect 3973 6199 4031 6205
rect 4433 6205 4445 6208
rect 4479 6236 4491 6239
rect 7926 6236 7932 6248
rect 4479 6208 7932 6236
rect 4479 6205 4491 6208
rect 4433 6199 4491 6205
rect 7926 6196 7932 6208
rect 7984 6196 7990 6248
rect 8220 6245 8248 6344
rect 9030 6332 9036 6384
rect 9088 6372 9094 6384
rect 9088 6344 9812 6372
rect 9088 6332 9094 6344
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 8404 6276 8493 6304
rect 8404 6248 8432 6276
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 9784 6313 9812 6344
rect 11054 6332 11060 6384
rect 11112 6372 11118 6384
rect 11882 6372 11888 6384
rect 11112 6344 11888 6372
rect 11112 6332 11118 6344
rect 11882 6332 11888 6344
rect 11940 6332 11946 6384
rect 9769 6307 9827 6313
rect 8628 6276 9720 6304
rect 8628 6264 8634 6276
rect 8205 6239 8263 6245
rect 8205 6205 8217 6239
rect 8251 6205 8263 6239
rect 8205 6199 8263 6205
rect 8386 6196 8392 6248
rect 8444 6196 8450 6248
rect 9214 6236 9220 6248
rect 9175 6208 9220 6236
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 9692 6236 9720 6276
rect 9769 6273 9781 6307
rect 9815 6273 9827 6307
rect 11974 6304 11980 6316
rect 9769 6267 9827 6273
rect 10796 6276 11980 6304
rect 10796 6236 10824 6276
rect 11974 6264 11980 6276
rect 12032 6264 12038 6316
rect 13648 6304 13676 6412
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 16945 6443 17003 6449
rect 16945 6409 16957 6443
rect 16991 6440 17003 6443
rect 17494 6440 17500 6452
rect 16991 6412 17500 6440
rect 16991 6409 17003 6412
rect 16945 6403 17003 6409
rect 17494 6400 17500 6412
rect 17552 6400 17558 6452
rect 19242 6400 19248 6452
rect 19300 6440 19306 6452
rect 20717 6443 20775 6449
rect 20717 6440 20729 6443
rect 19300 6412 20729 6440
rect 19300 6400 19306 6412
rect 20717 6409 20729 6412
rect 20763 6409 20775 6443
rect 20717 6403 20775 6409
rect 13906 6332 13912 6384
rect 13964 6372 13970 6384
rect 14366 6372 14372 6384
rect 13964 6344 14372 6372
rect 13964 6332 13970 6344
rect 14366 6332 14372 6344
rect 14424 6332 14430 6384
rect 16022 6332 16028 6384
rect 16080 6372 16086 6384
rect 16393 6375 16451 6381
rect 16393 6372 16405 6375
rect 16080 6344 16405 6372
rect 16080 6332 16086 6344
rect 16393 6341 16405 6344
rect 16439 6372 16451 6375
rect 16439 6344 18644 6372
rect 16439 6341 16451 6344
rect 16393 6335 16451 6341
rect 15013 6307 15071 6313
rect 15013 6304 15025 6307
rect 13648 6276 15025 6304
rect 15013 6273 15025 6276
rect 15059 6273 15071 6307
rect 17402 6304 17408 6316
rect 17363 6276 17408 6304
rect 15013 6267 15071 6273
rect 17402 6264 17408 6276
rect 17460 6264 17466 6316
rect 17497 6307 17555 6313
rect 17497 6273 17509 6307
rect 17543 6304 17555 6307
rect 17543 6276 17632 6304
rect 17543 6273 17555 6276
rect 17497 6267 17555 6273
rect 17604 6248 17632 6276
rect 17954 6264 17960 6316
rect 18012 6304 18018 6316
rect 18322 6304 18328 6316
rect 18012 6276 18328 6304
rect 18012 6264 18018 6276
rect 18322 6264 18328 6276
rect 18380 6304 18386 6316
rect 18616 6313 18644 6344
rect 18509 6307 18567 6313
rect 18509 6304 18521 6307
rect 18380 6276 18521 6304
rect 18380 6264 18386 6276
rect 18509 6273 18521 6276
rect 18555 6273 18567 6307
rect 18509 6267 18567 6273
rect 18601 6307 18659 6313
rect 18601 6273 18613 6307
rect 18647 6273 18659 6307
rect 18601 6267 18659 6273
rect 9692 6208 10824 6236
rect 11793 6239 11851 6245
rect 11793 6205 11805 6239
rect 11839 6236 11851 6239
rect 11839 6208 12480 6236
rect 11839 6205 11851 6208
rect 11793 6199 11851 6205
rect 3329 6171 3387 6177
rect 3329 6137 3341 6171
rect 3375 6168 3387 6171
rect 4985 6171 5043 6177
rect 4985 6168 4997 6171
rect 3375 6140 4997 6168
rect 3375 6137 3387 6140
rect 3329 6131 3387 6137
rect 4985 6137 4997 6140
rect 5031 6137 5043 6171
rect 4985 6131 5043 6137
rect 6086 6128 6092 6180
rect 6144 6168 6150 6180
rect 6144 6140 7972 6168
rect 6144 6128 6150 6140
rect 1946 6100 1952 6112
rect 1907 6072 1952 6100
rect 1946 6060 1952 6072
rect 2004 6060 2010 6112
rect 2314 6100 2320 6112
rect 2275 6072 2320 6100
rect 2314 6060 2320 6072
rect 2372 6060 2378 6112
rect 2406 6060 2412 6112
rect 2464 6100 2470 6112
rect 3234 6100 3240 6112
rect 2464 6072 2509 6100
rect 3195 6072 3240 6100
rect 2464 6060 2470 6072
rect 3234 6060 3240 6072
rect 3292 6060 3298 6112
rect 4062 6100 4068 6112
rect 4023 6072 4068 6100
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 5445 6103 5503 6109
rect 5445 6069 5457 6103
rect 5491 6100 5503 6103
rect 5905 6103 5963 6109
rect 5905 6100 5917 6103
rect 5491 6072 5917 6100
rect 5491 6069 5503 6072
rect 5445 6063 5503 6069
rect 5905 6069 5917 6072
rect 5951 6069 5963 6103
rect 5905 6063 5963 6069
rect 6273 6103 6331 6109
rect 6273 6069 6285 6103
rect 6319 6100 6331 6103
rect 6638 6100 6644 6112
rect 6319 6072 6644 6100
rect 6319 6069 6331 6072
rect 6273 6063 6331 6069
rect 6638 6060 6644 6072
rect 6696 6060 6702 6112
rect 6825 6103 6883 6109
rect 6825 6069 6837 6103
rect 6871 6100 6883 6103
rect 7374 6100 7380 6112
rect 6871 6072 7380 6100
rect 6871 6069 6883 6072
rect 6825 6063 6883 6069
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 7742 6060 7748 6112
rect 7800 6100 7806 6112
rect 7837 6103 7895 6109
rect 7837 6100 7849 6103
rect 7800 6072 7849 6100
rect 7800 6060 7806 6072
rect 7837 6069 7849 6072
rect 7883 6069 7895 6103
rect 7944 6100 7972 6140
rect 8018 6128 8024 6180
rect 8076 6168 8082 6180
rect 8297 6171 8355 6177
rect 8297 6168 8309 6171
rect 8076 6140 8309 6168
rect 8076 6128 8082 6140
rect 8297 6137 8309 6140
rect 8343 6168 8355 6171
rect 8570 6168 8576 6180
rect 8343 6140 8576 6168
rect 8343 6137 8355 6140
rect 8297 6131 8355 6137
rect 8570 6128 8576 6140
rect 8628 6128 8634 6180
rect 9490 6128 9496 6180
rect 9548 6168 9554 6180
rect 10014 6171 10072 6177
rect 10014 6168 10026 6171
rect 9548 6140 10026 6168
rect 9548 6128 9554 6140
rect 10014 6137 10026 6140
rect 10060 6137 10072 6171
rect 11882 6168 11888 6180
rect 10014 6131 10072 6137
rect 10980 6140 11888 6168
rect 9306 6100 9312 6112
rect 7944 6072 9312 6100
rect 7837 6063 7895 6069
rect 9306 6060 9312 6072
rect 9364 6060 9370 6112
rect 9401 6103 9459 6109
rect 9401 6069 9413 6103
rect 9447 6100 9459 6103
rect 10980 6100 11008 6140
rect 11882 6128 11888 6140
rect 11940 6128 11946 6180
rect 12452 6168 12480 6208
rect 12526 6196 12532 6248
rect 12584 6236 12590 6248
rect 12621 6239 12679 6245
rect 12621 6236 12633 6239
rect 12584 6208 12633 6236
rect 12584 6196 12590 6208
rect 12621 6205 12633 6208
rect 12667 6205 12679 6239
rect 12621 6199 12679 6205
rect 12888 6239 12946 6245
rect 12888 6205 12900 6239
rect 12934 6236 12946 6239
rect 13814 6236 13820 6248
rect 12934 6208 13820 6236
rect 12934 6205 12946 6208
rect 12888 6199 12946 6205
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 14458 6236 14464 6248
rect 14419 6208 14464 6236
rect 14458 6196 14464 6208
rect 14516 6196 14522 6248
rect 14568 6208 15516 6236
rect 12452 6140 12940 6168
rect 9447 6072 11008 6100
rect 9447 6069 9459 6072
rect 9401 6063 9459 6069
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 11149 6103 11207 6109
rect 11149 6100 11161 6103
rect 11112 6072 11161 6100
rect 11112 6060 11118 6072
rect 11149 6069 11161 6072
rect 11195 6069 11207 6103
rect 11149 6063 11207 6069
rect 11977 6103 12035 6109
rect 11977 6069 11989 6103
rect 12023 6100 12035 6103
rect 12802 6100 12808 6112
rect 12023 6072 12808 6100
rect 12023 6069 12035 6072
rect 11977 6063 12035 6069
rect 12802 6060 12808 6072
rect 12860 6060 12866 6112
rect 12912 6100 12940 6140
rect 12986 6128 12992 6180
rect 13044 6168 13050 6180
rect 14568 6168 14596 6208
rect 13044 6140 14596 6168
rect 15280 6171 15338 6177
rect 13044 6128 13050 6140
rect 15280 6137 15292 6171
rect 15326 6168 15338 6171
rect 15378 6168 15384 6180
rect 15326 6140 15384 6168
rect 15326 6137 15338 6140
rect 15280 6131 15338 6137
rect 15378 6128 15384 6140
rect 15436 6128 15442 6180
rect 15488 6168 15516 6208
rect 17586 6196 17592 6248
rect 17644 6196 17650 6248
rect 17696 6208 18543 6236
rect 17696 6168 17724 6208
rect 15488 6140 17724 6168
rect 17954 6128 17960 6180
rect 18012 6168 18018 6180
rect 18417 6171 18475 6177
rect 18417 6168 18429 6171
rect 18012 6140 18429 6168
rect 18012 6128 18018 6140
rect 18417 6137 18429 6140
rect 18463 6137 18475 6171
rect 18515 6168 18543 6208
rect 18874 6196 18880 6248
rect 18932 6236 18938 6248
rect 19150 6236 19156 6248
rect 18932 6208 19156 6236
rect 18932 6196 18938 6208
rect 19150 6196 19156 6208
rect 19208 6236 19214 6248
rect 19337 6239 19395 6245
rect 19337 6236 19349 6239
rect 19208 6208 19349 6236
rect 19208 6196 19214 6208
rect 19337 6205 19349 6208
rect 19383 6205 19395 6239
rect 20438 6236 20444 6248
rect 19337 6199 19395 6205
rect 19444 6208 20444 6236
rect 19444 6168 19472 6208
rect 20438 6196 20444 6208
rect 20496 6196 20502 6248
rect 18515 6140 19472 6168
rect 19604 6171 19662 6177
rect 18417 6131 18475 6137
rect 19604 6137 19616 6171
rect 19650 6168 19662 6171
rect 20254 6168 20260 6180
rect 19650 6140 20260 6168
rect 19650 6137 19662 6140
rect 19604 6131 19662 6137
rect 20254 6128 20260 6140
rect 20312 6128 20318 6180
rect 14090 6100 14096 6112
rect 12912 6072 14096 6100
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 14645 6103 14703 6109
rect 14645 6069 14657 6103
rect 14691 6100 14703 6103
rect 15194 6100 15200 6112
rect 14691 6072 15200 6100
rect 14691 6069 14703 6072
rect 14645 6063 14703 6069
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 17313 6103 17371 6109
rect 17313 6069 17325 6103
rect 17359 6100 17371 6103
rect 17770 6100 17776 6112
rect 17359 6072 17776 6100
rect 17359 6069 17371 6072
rect 17313 6063 17371 6069
rect 17770 6060 17776 6072
rect 17828 6060 17834 6112
rect 18046 6100 18052 6112
rect 18007 6072 18052 6100
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 18322 6060 18328 6112
rect 18380 6100 18386 6112
rect 20806 6100 20812 6112
rect 18380 6072 20812 6100
rect 18380 6060 18386 6072
rect 20806 6060 20812 6072
rect 20864 6060 20870 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 3694 5856 3700 5908
rect 3752 5896 3758 5908
rect 5721 5899 5779 5905
rect 3752 5868 5488 5896
rect 3752 5856 3758 5868
rect 1394 5788 1400 5840
rect 1452 5828 1458 5840
rect 1857 5831 1915 5837
rect 1857 5828 1869 5831
rect 1452 5800 1869 5828
rect 1452 5788 1458 5800
rect 1857 5797 1869 5800
rect 1903 5797 1915 5831
rect 4332 5831 4390 5837
rect 1857 5791 1915 5797
rect 2332 5800 4108 5828
rect 1581 5763 1639 5769
rect 1581 5729 1593 5763
rect 1627 5760 1639 5763
rect 1946 5760 1952 5772
rect 1627 5732 1952 5760
rect 1627 5729 1639 5732
rect 1581 5723 1639 5729
rect 1946 5720 1952 5732
rect 2004 5720 2010 5772
rect 1854 5652 1860 5704
rect 1912 5692 1918 5704
rect 2332 5701 2360 5800
rect 2584 5763 2642 5769
rect 2584 5729 2596 5763
rect 2630 5760 2642 5763
rect 3878 5760 3884 5772
rect 2630 5732 3884 5760
rect 2630 5729 2642 5732
rect 2584 5723 2642 5729
rect 3878 5720 3884 5732
rect 3936 5720 3942 5772
rect 4080 5769 4108 5800
rect 4332 5797 4344 5831
rect 4378 5828 4390 5831
rect 4706 5828 4712 5840
rect 4378 5800 4712 5828
rect 4378 5797 4390 5800
rect 4332 5791 4390 5797
rect 4706 5788 4712 5800
rect 4764 5788 4770 5840
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5760 4123 5763
rect 5460 5760 5488 5868
rect 5721 5865 5733 5899
rect 5767 5896 5779 5899
rect 6086 5896 6092 5908
rect 5767 5868 6092 5896
rect 5767 5865 5779 5868
rect 5721 5859 5779 5865
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 6178 5856 6184 5908
rect 6236 5896 6242 5908
rect 7193 5899 7251 5905
rect 7193 5896 7205 5899
rect 6236 5868 7205 5896
rect 6236 5856 6242 5868
rect 7193 5865 7205 5868
rect 7239 5865 7251 5899
rect 7193 5859 7251 5865
rect 7282 5856 7288 5908
rect 7340 5896 7346 5908
rect 7653 5899 7711 5905
rect 7653 5896 7665 5899
rect 7340 5868 7665 5896
rect 7340 5856 7346 5868
rect 7653 5865 7665 5868
rect 7699 5865 7711 5899
rect 7653 5859 7711 5865
rect 8205 5899 8263 5905
rect 8205 5865 8217 5899
rect 8251 5865 8263 5899
rect 8570 5896 8576 5908
rect 8531 5868 8576 5896
rect 8205 5859 8263 5865
rect 5534 5788 5540 5840
rect 5592 5828 5598 5840
rect 8220 5828 8248 5859
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 9306 5856 9312 5908
rect 9364 5896 9370 5908
rect 11793 5899 11851 5905
rect 9364 5868 11744 5896
rect 9364 5856 9370 5868
rect 9944 5831 10002 5837
rect 5592 5800 8248 5828
rect 8312 5800 9904 5828
rect 5592 5788 5598 5800
rect 6454 5760 6460 5772
rect 4111 5732 5396 5760
rect 5460 5732 6460 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 2317 5695 2375 5701
rect 2317 5692 2329 5695
rect 1912 5664 2329 5692
rect 1912 5652 1918 5664
rect 2317 5661 2329 5664
rect 2363 5661 2375 5695
rect 5368 5692 5396 5732
rect 6454 5720 6460 5732
rect 6512 5720 6518 5772
rect 6549 5763 6607 5769
rect 6549 5729 6561 5763
rect 6595 5729 6607 5763
rect 6549 5723 6607 5729
rect 6641 5763 6699 5769
rect 6641 5729 6653 5763
rect 6687 5760 6699 5763
rect 7282 5760 7288 5772
rect 6687 5732 7288 5760
rect 6687 5729 6699 5732
rect 6641 5723 6699 5729
rect 5718 5692 5724 5704
rect 5368 5664 5724 5692
rect 2317 5655 2375 5661
rect 5718 5652 5724 5664
rect 5776 5652 5782 5704
rect 5534 5584 5540 5636
rect 5592 5624 5598 5636
rect 6086 5624 6092 5636
rect 5592 5596 6092 5624
rect 5592 5584 5598 5596
rect 6086 5584 6092 5596
rect 6144 5584 6150 5636
rect 6564 5624 6592 5723
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 7374 5720 7380 5772
rect 7432 5760 7438 5772
rect 7561 5763 7619 5769
rect 7561 5760 7573 5763
rect 7432 5732 7573 5760
rect 7432 5720 7438 5732
rect 7561 5729 7573 5732
rect 7607 5729 7619 5763
rect 8312 5760 8340 5800
rect 7561 5723 7619 5729
rect 7760 5732 8340 5760
rect 8404 5732 8800 5760
rect 6730 5652 6736 5704
rect 6788 5692 6794 5704
rect 6788 5664 6833 5692
rect 6788 5652 6794 5664
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 7760 5692 7788 5732
rect 8404 5704 8432 5732
rect 7064 5664 7788 5692
rect 7837 5695 7895 5701
rect 7064 5652 7070 5664
rect 7837 5661 7849 5695
rect 7883 5692 7895 5695
rect 8386 5692 8392 5704
rect 7883 5664 8392 5692
rect 7883 5661 7895 5664
rect 7837 5655 7895 5661
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 8772 5701 8800 5732
rect 9030 5720 9036 5772
rect 9088 5760 9094 5772
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9088 5732 9689 5760
rect 9088 5720 9094 5732
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 9876 5760 9904 5800
rect 9944 5797 9956 5831
rect 9990 5828 10002 5831
rect 11054 5828 11060 5840
rect 9990 5800 11060 5828
rect 9990 5797 10002 5800
rect 9944 5791 10002 5797
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 11716 5837 11744 5868
rect 11793 5865 11805 5899
rect 11839 5896 11851 5899
rect 12342 5896 12348 5908
rect 11839 5868 12348 5896
rect 11839 5865 11851 5868
rect 11793 5859 11851 5865
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 12802 5856 12808 5908
rect 12860 5896 12866 5908
rect 12860 5868 14044 5896
rect 12860 5856 12866 5868
rect 11701 5831 11759 5837
rect 11701 5797 11713 5831
rect 11747 5828 11759 5831
rect 12986 5828 12992 5840
rect 11747 5800 12992 5828
rect 11747 5797 11759 5800
rect 11701 5791 11759 5797
rect 12986 5788 12992 5800
rect 13044 5788 13050 5840
rect 13354 5837 13360 5840
rect 13348 5791 13360 5837
rect 13412 5828 13418 5840
rect 14016 5828 14044 5868
rect 14090 5856 14096 5908
rect 14148 5896 14154 5908
rect 15010 5896 15016 5908
rect 14148 5868 15016 5896
rect 14148 5856 14154 5868
rect 15010 5856 15016 5868
rect 15068 5856 15074 5908
rect 15473 5899 15531 5905
rect 15473 5865 15485 5899
rect 15519 5865 15531 5899
rect 15473 5859 15531 5865
rect 15841 5899 15899 5905
rect 15841 5865 15853 5899
rect 15887 5896 15899 5899
rect 16114 5896 16120 5908
rect 15887 5868 16120 5896
rect 15887 5865 15899 5868
rect 15841 5859 15899 5865
rect 15488 5828 15516 5859
rect 16114 5856 16120 5868
rect 16172 5856 16178 5908
rect 17696 5868 17908 5896
rect 17696 5828 17724 5868
rect 13412 5800 13448 5828
rect 14016 5800 15424 5828
rect 15488 5800 17724 5828
rect 17880 5828 17908 5868
rect 18046 5856 18052 5908
rect 18104 5896 18110 5908
rect 18785 5899 18843 5905
rect 18785 5896 18797 5899
rect 18104 5868 18797 5896
rect 18104 5856 18110 5868
rect 18785 5865 18797 5868
rect 18831 5865 18843 5899
rect 19794 5896 19800 5908
rect 19755 5868 19800 5896
rect 18785 5859 18843 5865
rect 19794 5856 19800 5868
rect 19852 5896 19858 5908
rect 20622 5896 20628 5908
rect 19852 5868 20628 5896
rect 19852 5856 19858 5868
rect 20622 5856 20628 5868
rect 20680 5856 20686 5908
rect 18877 5831 18935 5837
rect 18877 5828 18889 5831
rect 17880 5800 18889 5828
rect 13354 5788 13360 5791
rect 13412 5788 13418 5800
rect 11606 5760 11612 5772
rect 9876 5732 11612 5760
rect 9677 5723 9735 5729
rect 11606 5720 11612 5732
rect 11664 5720 11670 5772
rect 12342 5720 12348 5772
rect 12400 5760 12406 5772
rect 12529 5763 12587 5769
rect 12529 5760 12541 5763
rect 12400 5732 12541 5760
rect 12400 5720 12406 5732
rect 12529 5729 12541 5732
rect 12575 5729 12587 5763
rect 12529 5723 12587 5729
rect 12618 5720 12624 5772
rect 12676 5760 12682 5772
rect 13081 5763 13139 5769
rect 13081 5760 13093 5763
rect 12676 5732 13093 5760
rect 12676 5720 12682 5732
rect 13081 5729 13093 5732
rect 13127 5760 13139 5763
rect 13170 5760 13176 5772
rect 13127 5732 13176 5760
rect 13127 5729 13139 5732
rect 13081 5723 13139 5729
rect 13170 5720 13176 5732
rect 13228 5720 13234 5772
rect 14182 5720 14188 5772
rect 14240 5760 14246 5772
rect 15102 5760 15108 5772
rect 14240 5732 15108 5760
rect 14240 5720 14246 5732
rect 15102 5720 15108 5732
rect 15160 5720 15166 5772
rect 15396 5760 15424 5800
rect 18877 5797 18889 5800
rect 18923 5797 18935 5831
rect 19886 5828 19892 5840
rect 19799 5800 19892 5828
rect 18877 5791 18935 5797
rect 19886 5788 19892 5800
rect 19944 5828 19950 5840
rect 21266 5828 21272 5840
rect 19944 5800 21272 5828
rect 19944 5788 19950 5800
rect 21266 5788 21272 5800
rect 21324 5788 21330 5840
rect 15746 5760 15752 5772
rect 15396 5732 15752 5760
rect 15746 5720 15752 5732
rect 15804 5720 15810 5772
rect 16761 5763 16819 5769
rect 16761 5729 16773 5763
rect 16807 5760 16819 5763
rect 16850 5760 16856 5772
rect 16807 5732 16856 5760
rect 16807 5729 16819 5732
rect 16761 5723 16819 5729
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 17034 5769 17040 5772
rect 17028 5760 17040 5769
rect 16995 5732 17040 5760
rect 17028 5723 17040 5732
rect 17034 5720 17040 5723
rect 17092 5720 17098 5772
rect 18322 5720 18328 5772
rect 18380 5760 18386 5772
rect 20438 5760 20444 5772
rect 18380 5732 20444 5760
rect 18380 5720 18386 5732
rect 20438 5720 20444 5732
rect 20496 5720 20502 5772
rect 8665 5695 8723 5701
rect 8665 5692 8677 5695
rect 8496 5664 8677 5692
rect 8110 5624 8116 5636
rect 6564 5596 8116 5624
rect 8110 5584 8116 5596
rect 8168 5584 8174 5636
rect 3510 5516 3516 5568
rect 3568 5556 3574 5568
rect 3697 5559 3755 5565
rect 3697 5556 3709 5559
rect 3568 5528 3709 5556
rect 3568 5516 3574 5528
rect 3697 5525 3709 5528
rect 3743 5525 3755 5559
rect 3697 5519 3755 5525
rect 3878 5516 3884 5568
rect 3936 5556 3942 5568
rect 5074 5556 5080 5568
rect 3936 5528 5080 5556
rect 3936 5516 3942 5528
rect 5074 5516 5080 5528
rect 5132 5556 5138 5568
rect 5445 5559 5503 5565
rect 5445 5556 5457 5559
rect 5132 5528 5457 5556
rect 5132 5516 5138 5528
rect 5445 5525 5457 5528
rect 5491 5525 5503 5559
rect 5445 5519 5503 5525
rect 6181 5559 6239 5565
rect 6181 5525 6193 5559
rect 6227 5556 6239 5559
rect 7006 5556 7012 5568
rect 6227 5528 7012 5556
rect 6227 5525 6239 5528
rect 6181 5519 6239 5525
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 7834 5516 7840 5568
rect 7892 5556 7898 5568
rect 8496 5556 8524 5664
rect 8665 5661 8677 5664
rect 8711 5661 8723 5695
rect 8665 5655 8723 5661
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5661 8815 5695
rect 8757 5655 8815 5661
rect 11977 5695 12035 5701
rect 11977 5661 11989 5695
rect 12023 5692 12035 5695
rect 12158 5692 12164 5704
rect 12023 5664 12164 5692
rect 12023 5661 12035 5664
rect 11977 5655 12035 5661
rect 12158 5652 12164 5664
rect 12216 5652 12222 5704
rect 14737 5695 14795 5701
rect 14737 5661 14749 5695
rect 14783 5661 14795 5695
rect 14737 5655 14795 5661
rect 10686 5584 10692 5636
rect 10744 5624 10750 5636
rect 12618 5624 12624 5636
rect 10744 5596 12624 5624
rect 10744 5584 10750 5596
rect 12618 5584 12624 5596
rect 12676 5584 12682 5636
rect 12713 5627 12771 5633
rect 12713 5593 12725 5627
rect 12759 5624 12771 5627
rect 13078 5624 13084 5636
rect 12759 5596 13084 5624
rect 12759 5593 12771 5596
rect 12713 5587 12771 5593
rect 13078 5584 13084 5596
rect 13136 5584 13142 5636
rect 14458 5624 14464 5636
rect 14419 5596 14464 5624
rect 14458 5584 14464 5596
rect 14516 5584 14522 5636
rect 14752 5624 14780 5655
rect 15194 5652 15200 5704
rect 15252 5692 15258 5704
rect 15933 5695 15991 5701
rect 15933 5692 15945 5695
rect 15252 5664 15945 5692
rect 15252 5652 15258 5664
rect 15933 5661 15945 5664
rect 15979 5661 15991 5695
rect 15933 5655 15991 5661
rect 16022 5652 16028 5704
rect 16080 5692 16086 5704
rect 16080 5664 16125 5692
rect 16080 5652 16086 5664
rect 18138 5652 18144 5704
rect 18196 5692 18202 5704
rect 18969 5695 19027 5701
rect 18969 5692 18981 5695
rect 18196 5664 18981 5692
rect 18196 5652 18202 5664
rect 18969 5661 18981 5664
rect 19015 5661 19027 5695
rect 18969 5655 19027 5661
rect 19518 5652 19524 5704
rect 19576 5692 19582 5704
rect 19981 5695 20039 5701
rect 19981 5692 19993 5695
rect 19576 5664 19993 5692
rect 19576 5652 19582 5664
rect 19981 5661 19993 5664
rect 20027 5661 20039 5695
rect 19981 5655 20039 5661
rect 16574 5624 16580 5636
rect 14752 5596 16580 5624
rect 16574 5584 16580 5596
rect 16632 5584 16638 5636
rect 17770 5584 17776 5636
rect 17828 5624 17834 5636
rect 18417 5627 18475 5633
rect 18417 5624 18429 5627
rect 17828 5596 18429 5624
rect 17828 5584 17834 5596
rect 18417 5593 18429 5596
rect 18463 5593 18475 5627
rect 18417 5587 18475 5593
rect 7892 5528 8524 5556
rect 7892 5516 7898 5528
rect 9582 5516 9588 5568
rect 9640 5556 9646 5568
rect 10410 5556 10416 5568
rect 9640 5528 10416 5556
rect 9640 5516 9646 5528
rect 10410 5516 10416 5528
rect 10468 5556 10474 5568
rect 11057 5559 11115 5565
rect 11057 5556 11069 5559
rect 10468 5528 11069 5556
rect 10468 5516 10474 5528
rect 11057 5525 11069 5528
rect 11103 5525 11115 5559
rect 11057 5519 11115 5525
rect 11146 5516 11152 5568
rect 11204 5556 11210 5568
rect 11333 5559 11391 5565
rect 11333 5556 11345 5559
rect 11204 5528 11345 5556
rect 11204 5516 11210 5528
rect 11333 5525 11345 5528
rect 11379 5525 11391 5559
rect 11333 5519 11391 5525
rect 12158 5516 12164 5568
rect 12216 5556 12222 5568
rect 12986 5556 12992 5568
rect 12216 5528 12992 5556
rect 12216 5516 12222 5528
rect 12986 5516 12992 5528
rect 13044 5516 13050 5568
rect 13722 5516 13728 5568
rect 13780 5556 13786 5568
rect 17494 5556 17500 5568
rect 13780 5528 17500 5556
rect 13780 5516 13786 5528
rect 17494 5516 17500 5528
rect 17552 5516 17558 5568
rect 17678 5516 17684 5568
rect 17736 5556 17742 5568
rect 18141 5559 18199 5565
rect 18141 5556 18153 5559
rect 17736 5528 18153 5556
rect 17736 5516 17742 5528
rect 18141 5525 18153 5528
rect 18187 5525 18199 5559
rect 18141 5519 18199 5525
rect 18690 5516 18696 5568
rect 18748 5556 18754 5568
rect 19429 5559 19487 5565
rect 19429 5556 19441 5559
rect 18748 5528 19441 5556
rect 18748 5516 18754 5528
rect 19429 5525 19441 5528
rect 19475 5525 19487 5559
rect 19429 5519 19487 5525
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 1578 5352 1584 5364
rect 1539 5324 1584 5352
rect 1578 5312 1584 5324
rect 1636 5312 1642 5364
rect 3234 5312 3240 5364
rect 3292 5352 3298 5364
rect 3605 5355 3663 5361
rect 3605 5352 3617 5355
rect 3292 5324 3617 5352
rect 3292 5312 3298 5324
rect 3605 5321 3617 5324
rect 3651 5321 3663 5355
rect 3605 5315 3663 5321
rect 4890 5312 4896 5364
rect 4948 5352 4954 5364
rect 5258 5352 5264 5364
rect 4948 5324 5264 5352
rect 4948 5312 4954 5324
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 5721 5355 5779 5361
rect 5721 5321 5733 5355
rect 5767 5352 5779 5355
rect 7190 5352 7196 5364
rect 5767 5324 7196 5352
rect 5767 5321 5779 5324
rect 5721 5315 5779 5321
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 8202 5352 8208 5364
rect 8163 5324 8208 5352
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 9030 5352 9036 5364
rect 8772 5324 9036 5352
rect 3326 5244 3332 5296
rect 3384 5284 3390 5296
rect 6270 5284 6276 5296
rect 3384 5256 6276 5284
rect 3384 5244 3390 5256
rect 6270 5244 6276 5256
rect 6328 5244 6334 5296
rect 1854 5176 1860 5228
rect 1912 5216 1918 5228
rect 1949 5219 2007 5225
rect 1949 5216 1961 5219
rect 1912 5188 1961 5216
rect 1912 5176 1918 5188
rect 1949 5185 1961 5188
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 3878 5176 3884 5228
rect 3936 5216 3942 5228
rect 4157 5219 4215 5225
rect 4157 5216 4169 5219
rect 3936 5188 4169 5216
rect 3936 5176 3942 5188
rect 4157 5185 4169 5188
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 4706 5176 4712 5228
rect 4764 5216 4770 5228
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 4764 5188 5181 5216
rect 4764 5176 4770 5188
rect 5169 5185 5181 5188
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 3694 5148 3700 5160
rect 1443 5120 3700 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 3973 5151 4031 5157
rect 3973 5117 3985 5151
rect 4019 5148 4031 5151
rect 4062 5148 4068 5160
rect 4019 5120 4068 5148
rect 4019 5117 4031 5120
rect 3973 5111 4031 5117
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 4246 5108 4252 5160
rect 4304 5148 4310 5160
rect 4985 5151 5043 5157
rect 4985 5148 4997 5151
rect 4304 5120 4997 5148
rect 4304 5108 4310 5120
rect 4985 5117 4997 5120
rect 5031 5148 5043 5151
rect 5074 5148 5080 5160
rect 5031 5120 5080 5148
rect 5031 5117 5043 5120
rect 4985 5111 5043 5117
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 6089 5151 6147 5157
rect 6089 5148 6101 5151
rect 6052 5120 6101 5148
rect 6052 5108 6058 5120
rect 6089 5117 6101 5120
rect 6135 5117 6147 5151
rect 6089 5111 6147 5117
rect 6178 5108 6184 5160
rect 6236 5148 6242 5160
rect 6236 5120 6281 5148
rect 6236 5108 6242 5120
rect 2222 5089 2228 5092
rect 2216 5080 2228 5089
rect 2183 5052 2228 5080
rect 2216 5043 2228 5052
rect 2222 5040 2228 5043
rect 2280 5040 2286 5092
rect 4338 5040 4344 5092
rect 4396 5080 4402 5092
rect 5534 5080 5540 5092
rect 4396 5052 5540 5080
rect 4396 5040 4402 5052
rect 5534 5040 5540 5052
rect 5592 5040 5598 5092
rect 6380 5080 6408 5179
rect 8110 5176 8116 5228
rect 8168 5216 8174 5228
rect 8662 5216 8668 5228
rect 8168 5188 8668 5216
rect 8168 5176 8174 5188
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 6822 5148 6828 5160
rect 6783 5120 6828 5148
rect 6822 5108 6828 5120
rect 6880 5148 6886 5160
rect 8772 5157 8800 5324
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 9122 5312 9128 5364
rect 9180 5352 9186 5364
rect 9180 5324 10640 5352
rect 9180 5312 9186 5324
rect 10612 5284 10640 5324
rect 10686 5312 10692 5364
rect 10744 5352 10750 5364
rect 10744 5324 12388 5352
rect 10744 5312 10750 5324
rect 12360 5284 12388 5324
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 14550 5352 14556 5364
rect 12492 5324 14556 5352
rect 12492 5312 12498 5324
rect 14550 5312 14556 5324
rect 14608 5312 14614 5364
rect 16850 5352 16856 5364
rect 15856 5324 16856 5352
rect 15657 5287 15715 5293
rect 15657 5284 15669 5287
rect 10612 5256 12296 5284
rect 12360 5256 15669 5284
rect 11609 5219 11667 5225
rect 11609 5185 11621 5219
rect 11655 5216 11667 5219
rect 12158 5216 12164 5228
rect 11655 5188 12164 5216
rect 11655 5185 11667 5188
rect 11609 5179 11667 5185
rect 12158 5176 12164 5188
rect 12216 5176 12222 5228
rect 12268 5216 12296 5256
rect 15657 5253 15669 5256
rect 15703 5253 15715 5287
rect 15657 5247 15715 5253
rect 12897 5219 12955 5225
rect 12897 5216 12909 5219
rect 12268 5188 12909 5216
rect 12897 5185 12909 5188
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 12986 5176 12992 5228
rect 13044 5216 13050 5228
rect 13081 5219 13139 5225
rect 13081 5216 13093 5219
rect 13044 5188 13093 5216
rect 13044 5176 13050 5188
rect 13081 5185 13093 5188
rect 13127 5216 13139 5219
rect 13354 5216 13360 5228
rect 13127 5188 13360 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 13354 5176 13360 5188
rect 13412 5216 13418 5228
rect 14369 5219 14427 5225
rect 14369 5216 14381 5219
rect 13412 5188 14381 5216
rect 13412 5176 13418 5188
rect 14369 5185 14381 5188
rect 14415 5216 14427 5219
rect 14550 5216 14556 5228
rect 14415 5188 14556 5216
rect 14415 5185 14427 5188
rect 14369 5179 14427 5185
rect 14550 5176 14556 5188
rect 14608 5176 14614 5228
rect 14642 5176 14648 5228
rect 14700 5216 14706 5228
rect 15289 5219 15347 5225
rect 15289 5216 15301 5219
rect 14700 5188 15301 5216
rect 14700 5176 14706 5188
rect 15289 5185 15301 5188
rect 15335 5185 15347 5219
rect 15289 5179 15347 5185
rect 15378 5176 15384 5228
rect 15436 5216 15442 5228
rect 15856 5225 15884 5324
rect 16850 5312 16856 5324
rect 16908 5312 16914 5364
rect 17034 5312 17040 5364
rect 17092 5352 17098 5364
rect 17221 5355 17279 5361
rect 17221 5352 17233 5355
rect 17092 5324 17233 5352
rect 17092 5312 17098 5324
rect 17221 5321 17233 5324
rect 17267 5321 17279 5355
rect 17221 5315 17279 5321
rect 17773 5355 17831 5361
rect 17773 5321 17785 5355
rect 17819 5352 17831 5355
rect 17954 5352 17960 5364
rect 17819 5324 17960 5352
rect 17819 5321 17831 5324
rect 17773 5315 17831 5321
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 19058 5312 19064 5364
rect 19116 5352 19122 5364
rect 20254 5352 20260 5364
rect 19116 5324 19932 5352
rect 20215 5324 20260 5352
rect 19116 5312 19122 5324
rect 15841 5219 15899 5225
rect 15436 5188 15481 5216
rect 15436 5176 15442 5188
rect 15841 5185 15853 5219
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 17497 5219 17555 5225
rect 17497 5185 17509 5219
rect 17543 5216 17555 5219
rect 17773 5219 17831 5225
rect 17773 5216 17785 5219
rect 17543 5188 17785 5216
rect 17543 5185 17555 5188
rect 17497 5179 17555 5185
rect 17773 5185 17785 5188
rect 17819 5185 17831 5219
rect 19904 5216 19932 5324
rect 20254 5312 20260 5324
rect 20312 5312 20318 5364
rect 20717 5219 20775 5225
rect 20717 5216 20729 5219
rect 17773 5179 17831 5185
rect 17880 5188 19012 5216
rect 19904 5188 20729 5216
rect 8757 5151 8815 5157
rect 8757 5148 8769 5151
rect 6880 5120 8769 5148
rect 6880 5108 6886 5120
rect 8757 5117 8769 5120
rect 8803 5117 8815 5151
rect 8757 5111 8815 5117
rect 9024 5151 9082 5157
rect 9024 5117 9036 5151
rect 9070 5148 9082 5151
rect 9582 5148 9588 5160
rect 9070 5120 9588 5148
rect 9070 5117 9082 5120
rect 9024 5111 9082 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 10134 5108 10140 5160
rect 10192 5148 10198 5160
rect 10413 5151 10471 5157
rect 10413 5148 10425 5151
rect 10192 5120 10425 5148
rect 10192 5108 10198 5120
rect 10413 5117 10425 5120
rect 10459 5117 10471 5151
rect 15197 5151 15255 5157
rect 15197 5148 15209 5151
rect 10413 5111 10471 5117
rect 11164 5120 15209 5148
rect 6730 5080 6736 5092
rect 6380 5052 6736 5080
rect 6730 5040 6736 5052
rect 6788 5080 6794 5092
rect 7098 5089 7104 5092
rect 7092 5080 7104 5089
rect 6788 5052 7104 5080
rect 6788 5040 6794 5052
rect 7092 5043 7104 5052
rect 7098 5040 7104 5043
rect 7156 5040 7162 5092
rect 7466 5040 7472 5092
rect 7524 5080 7530 5092
rect 8846 5080 8852 5092
rect 7524 5052 8852 5080
rect 7524 5040 7530 5052
rect 8846 5040 8852 5052
rect 8904 5040 8910 5092
rect 9398 5080 9404 5092
rect 8947 5052 9404 5080
rect 3329 5015 3387 5021
rect 3329 4981 3341 5015
rect 3375 5012 3387 5015
rect 3602 5012 3608 5024
rect 3375 4984 3608 5012
rect 3375 4981 3387 4984
rect 3329 4975 3387 4981
rect 3602 4972 3608 4984
rect 3660 4972 3666 5024
rect 4065 5015 4123 5021
rect 4065 4981 4077 5015
rect 4111 5012 4123 5015
rect 4617 5015 4675 5021
rect 4617 5012 4629 5015
rect 4111 4984 4629 5012
rect 4111 4981 4123 4984
rect 4065 4975 4123 4981
rect 4617 4981 4629 4984
rect 4663 4981 4675 5015
rect 4617 4975 4675 4981
rect 5077 5015 5135 5021
rect 5077 4981 5089 5015
rect 5123 5012 5135 5015
rect 8947 5012 8975 5052
rect 9398 5040 9404 5052
rect 9456 5080 9462 5092
rect 11164 5080 11192 5120
rect 15197 5117 15209 5120
rect 15243 5117 15255 5151
rect 17880 5148 17908 5188
rect 15197 5111 15255 5117
rect 15295 5120 17908 5148
rect 18049 5151 18107 5157
rect 9456 5052 11192 5080
rect 11333 5083 11391 5089
rect 9456 5040 9462 5052
rect 11333 5049 11345 5083
rect 11379 5080 11391 5083
rect 11606 5080 11612 5092
rect 11379 5052 11612 5080
rect 11379 5049 11391 5052
rect 11333 5043 11391 5049
rect 11606 5040 11612 5052
rect 11664 5080 11670 5092
rect 15295 5080 15323 5120
rect 18049 5117 18061 5151
rect 18095 5117 18107 5151
rect 18874 5148 18880 5160
rect 18835 5120 18880 5148
rect 18049 5111 18107 5117
rect 11664 5052 15323 5080
rect 15657 5083 15715 5089
rect 11664 5040 11670 5052
rect 15657 5049 15669 5083
rect 15703 5080 15715 5083
rect 15838 5080 15844 5092
rect 15703 5052 15844 5080
rect 15703 5049 15715 5052
rect 15657 5043 15715 5049
rect 15838 5040 15844 5052
rect 15896 5040 15902 5092
rect 16022 5040 16028 5092
rect 16080 5089 16086 5092
rect 16080 5083 16144 5089
rect 16080 5049 16098 5083
rect 16132 5049 16144 5083
rect 18064 5080 18092 5111
rect 18874 5108 18880 5120
rect 18932 5108 18938 5160
rect 18984 5148 19012 5188
rect 20717 5185 20729 5188
rect 20763 5185 20775 5219
rect 20717 5179 20775 5185
rect 20070 5148 20076 5160
rect 18984 5120 20076 5148
rect 20070 5108 20076 5120
rect 20128 5108 20134 5160
rect 20530 5148 20536 5160
rect 20491 5120 20536 5148
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 18782 5080 18788 5092
rect 18064 5052 18788 5080
rect 16080 5043 16144 5049
rect 16080 5040 16086 5043
rect 18782 5040 18788 5052
rect 18840 5040 18846 5092
rect 19144 5083 19202 5089
rect 19144 5049 19156 5083
rect 19190 5080 19202 5083
rect 19702 5080 19708 5092
rect 19190 5052 19708 5080
rect 19190 5049 19202 5052
rect 19144 5043 19202 5049
rect 19702 5040 19708 5052
rect 19760 5040 19766 5092
rect 5123 4984 8975 5012
rect 5123 4981 5135 4984
rect 5077 4975 5135 4981
rect 9030 4972 9036 5024
rect 9088 5012 9094 5024
rect 10042 5012 10048 5024
rect 9088 4984 10048 5012
rect 9088 4972 9094 4984
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 10137 5015 10195 5021
rect 10137 4981 10149 5015
rect 10183 5012 10195 5015
rect 10410 5012 10416 5024
rect 10183 4984 10416 5012
rect 10183 4981 10195 4984
rect 10137 4975 10195 4981
rect 10410 4972 10416 4984
rect 10468 4972 10474 5024
rect 10597 5015 10655 5021
rect 10597 4981 10609 5015
rect 10643 5012 10655 5015
rect 10778 5012 10784 5024
rect 10643 4984 10784 5012
rect 10643 4981 10655 4984
rect 10597 4975 10655 4981
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 10870 4972 10876 5024
rect 10928 5012 10934 5024
rect 10965 5015 11023 5021
rect 10965 5012 10977 5015
rect 10928 4984 10977 5012
rect 10928 4972 10934 4984
rect 10965 4981 10977 4984
rect 11011 4981 11023 5015
rect 11422 5012 11428 5024
rect 11383 4984 11428 5012
rect 10965 4975 11023 4981
rect 11422 4972 11428 4984
rect 11480 4972 11486 5024
rect 12434 5012 12440 5024
rect 12395 4984 12440 5012
rect 12434 4972 12440 4984
rect 12492 4972 12498 5024
rect 12805 5015 12863 5021
rect 12805 4981 12817 5015
rect 12851 5012 12863 5015
rect 13262 5012 13268 5024
rect 12851 4984 13268 5012
rect 12851 4981 12863 4984
rect 12805 4975 12863 4981
rect 13262 4972 13268 4984
rect 13320 4972 13326 5024
rect 13725 5015 13783 5021
rect 13725 4981 13737 5015
rect 13771 5012 13783 5015
rect 13906 5012 13912 5024
rect 13771 4984 13912 5012
rect 13771 4981 13783 4984
rect 13725 4975 13783 4981
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 14090 5012 14096 5024
rect 14051 4984 14096 5012
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 14829 5015 14887 5021
rect 14240 4984 14285 5012
rect 14240 4972 14246 4984
rect 14829 4981 14841 5015
rect 14875 5012 14887 5015
rect 15194 5012 15200 5024
rect 14875 4984 15200 5012
rect 14875 4981 14887 4984
rect 14829 4975 14887 4981
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 18233 5015 18291 5021
rect 18233 4981 18245 5015
rect 18279 5012 18291 5015
rect 18506 5012 18512 5024
rect 18279 4984 18512 5012
rect 18279 4981 18291 4984
rect 18233 4975 18291 4981
rect 18506 4972 18512 4984
rect 18564 4972 18570 5024
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 2222 4768 2228 4820
rect 2280 4808 2286 4820
rect 2869 4811 2927 4817
rect 2869 4808 2881 4811
rect 2280 4780 2881 4808
rect 2280 4768 2286 4780
rect 2869 4777 2881 4780
rect 2915 4777 2927 4811
rect 3326 4808 3332 4820
rect 3287 4780 3332 4808
rect 2869 4771 2927 4777
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 4982 4808 4988 4820
rect 3752 4780 4988 4808
rect 3752 4768 3758 4780
rect 4982 4768 4988 4780
rect 5040 4768 5046 4820
rect 5077 4811 5135 4817
rect 5077 4777 5089 4811
rect 5123 4808 5135 4811
rect 5166 4808 5172 4820
rect 5123 4780 5172 4808
rect 5123 4777 5135 4780
rect 5077 4771 5135 4777
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 7098 4808 7104 4820
rect 5552 4780 6408 4808
rect 7059 4780 7104 4808
rect 1854 4740 1860 4752
rect 1504 4712 1860 4740
rect 1504 4681 1532 4712
rect 1854 4700 1860 4712
rect 1912 4700 1918 4752
rect 2884 4712 4108 4740
rect 2884 4684 2912 4712
rect 1489 4675 1547 4681
rect 1489 4641 1501 4675
rect 1535 4641 1547 4675
rect 1489 4635 1547 4641
rect 1756 4675 1814 4681
rect 1756 4641 1768 4675
rect 1802 4672 1814 4675
rect 2222 4672 2228 4684
rect 1802 4644 2228 4672
rect 1802 4641 1814 4644
rect 1756 4635 1814 4641
rect 2222 4632 2228 4644
rect 2280 4632 2286 4684
rect 2866 4632 2872 4684
rect 2924 4632 2930 4684
rect 4080 4681 4108 4712
rect 3421 4675 3479 4681
rect 3421 4641 3433 4675
rect 3467 4672 3479 4675
rect 4065 4675 4123 4681
rect 3467 4644 4016 4672
rect 3467 4641 3479 4644
rect 3421 4635 3479 4641
rect 3602 4604 3608 4616
rect 3563 4576 3608 4604
rect 3602 4564 3608 4576
rect 3660 4564 3666 4616
rect 3988 4604 4016 4644
rect 4065 4641 4077 4675
rect 4111 4672 4123 4675
rect 4246 4672 4252 4684
rect 4111 4644 4252 4672
rect 4111 4641 4123 4644
rect 4065 4635 4123 4641
rect 4246 4632 4252 4644
rect 4304 4632 4310 4684
rect 4706 4632 4712 4684
rect 4764 4672 4770 4684
rect 4985 4675 5043 4681
rect 4985 4672 4997 4675
rect 4764 4644 4997 4672
rect 4764 4632 4770 4644
rect 4985 4641 4997 4644
rect 5031 4672 5043 4675
rect 5442 4672 5448 4684
rect 5031 4644 5448 4672
rect 5031 4641 5043 4644
rect 4985 4635 5043 4641
rect 5442 4632 5448 4644
rect 5500 4632 5506 4684
rect 3988 4576 5120 4604
rect 3142 4496 3148 4548
rect 3200 4536 3206 4548
rect 4617 4539 4675 4545
rect 4617 4536 4629 4539
rect 3200 4508 4629 4536
rect 3200 4496 3206 4508
rect 4617 4505 4629 4508
rect 4663 4505 4675 4539
rect 5092 4536 5120 4576
rect 5166 4564 5172 4616
rect 5224 4604 5230 4616
rect 5261 4607 5319 4613
rect 5261 4604 5273 4607
rect 5224 4576 5273 4604
rect 5224 4564 5230 4576
rect 5261 4573 5273 4576
rect 5307 4604 5319 4607
rect 5552 4604 5580 4780
rect 5902 4700 5908 4752
rect 5960 4749 5966 4752
rect 5960 4743 6024 4749
rect 5960 4709 5978 4743
rect 6012 4740 6024 4743
rect 6270 4740 6276 4752
rect 6012 4712 6276 4740
rect 6012 4709 6024 4712
rect 5960 4703 6024 4709
rect 5960 4700 5966 4703
rect 6270 4700 6276 4712
rect 6328 4700 6334 4752
rect 6380 4740 6408 4780
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 7374 4808 7380 4820
rect 7335 4780 7380 4808
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 7742 4808 7748 4820
rect 7703 4780 7748 4808
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 7837 4811 7895 4817
rect 7837 4777 7849 4811
rect 7883 4808 7895 4811
rect 8389 4811 8447 4817
rect 8389 4808 8401 4811
rect 7883 4780 8401 4808
rect 7883 4777 7895 4780
rect 7837 4771 7895 4777
rect 8389 4777 8401 4780
rect 8435 4777 8447 4811
rect 8389 4771 8447 4777
rect 8757 4811 8815 4817
rect 8757 4777 8769 4811
rect 8803 4808 8815 4811
rect 8846 4808 8852 4820
rect 8803 4780 8852 4808
rect 8803 4777 8815 4780
rect 8757 4771 8815 4777
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 10134 4808 10140 4820
rect 10095 4780 10140 4808
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 10505 4811 10563 4817
rect 10505 4777 10517 4811
rect 10551 4777 10563 4811
rect 10870 4808 10876 4820
rect 10831 4780 10876 4808
rect 10505 4771 10563 4777
rect 10410 4740 10416 4752
rect 6380 4712 10416 4740
rect 10410 4700 10416 4712
rect 10468 4700 10474 4752
rect 10520 4740 10548 4771
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 10965 4811 11023 4817
rect 10965 4777 10977 4811
rect 11011 4808 11023 4811
rect 11146 4808 11152 4820
rect 11011 4780 11152 4808
rect 11011 4777 11023 4780
rect 10965 4771 11023 4777
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 11422 4768 11428 4820
rect 11480 4808 11486 4820
rect 12066 4808 12072 4820
rect 11480 4780 12072 4808
rect 11480 4768 11486 4780
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 12989 4811 13047 4817
rect 12989 4808 13001 4811
rect 12492 4780 13001 4808
rect 12492 4768 12498 4780
rect 12989 4777 13001 4780
rect 13035 4777 13047 4811
rect 13906 4808 13912 4820
rect 13867 4780 13912 4808
rect 12989 4771 13047 4777
rect 13906 4768 13912 4780
rect 13964 4768 13970 4820
rect 14001 4811 14059 4817
rect 14001 4777 14013 4811
rect 14047 4808 14059 4811
rect 15194 4808 15200 4820
rect 14047 4780 15200 4808
rect 14047 4777 14059 4780
rect 14001 4771 14059 4777
rect 15194 4768 15200 4780
rect 15252 4768 15258 4820
rect 16022 4768 16028 4820
rect 16080 4808 16086 4820
rect 16080 4780 17172 4808
rect 16080 4768 16086 4780
rect 11885 4743 11943 4749
rect 11885 4740 11897 4743
rect 10520 4712 11897 4740
rect 11885 4709 11897 4712
rect 11931 4709 11943 4743
rect 11885 4703 11943 4709
rect 12897 4743 12955 4749
rect 12897 4709 12909 4743
rect 12943 4740 12955 4743
rect 13078 4740 13084 4752
rect 12943 4712 13084 4740
rect 12943 4709 12955 4712
rect 12897 4703 12955 4709
rect 13078 4700 13084 4712
rect 13136 4700 13142 4752
rect 13357 4743 13415 4749
rect 13357 4709 13369 4743
rect 13403 4740 13415 4743
rect 17144 4740 17172 4780
rect 17218 4768 17224 4820
rect 17276 4808 17282 4820
rect 17405 4811 17463 4817
rect 17405 4808 17417 4811
rect 17276 4780 17417 4808
rect 17276 4768 17282 4780
rect 17405 4777 17417 4780
rect 17451 4777 17463 4811
rect 17770 4808 17776 4820
rect 17731 4780 17776 4808
rect 17405 4771 17463 4777
rect 17770 4768 17776 4780
rect 17828 4768 17834 4820
rect 18233 4811 18291 4817
rect 18233 4777 18245 4811
rect 18279 4808 18291 4811
rect 20349 4811 20407 4817
rect 20349 4808 20361 4811
rect 18279 4780 20361 4808
rect 18279 4777 18291 4780
rect 18233 4771 18291 4777
rect 20349 4777 20361 4780
rect 20395 4777 20407 4811
rect 20349 4771 20407 4777
rect 17313 4743 17371 4749
rect 17313 4740 17325 4743
rect 13403 4712 16896 4740
rect 17144 4712 17325 4740
rect 13403 4709 13415 4712
rect 13357 4703 13415 4709
rect 5718 4672 5724 4684
rect 5679 4644 5724 4672
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 6288 4672 6316 4700
rect 8849 4675 8907 4681
rect 6288 4644 7972 4672
rect 7944 4613 7972 4644
rect 8849 4641 8861 4675
rect 8895 4672 8907 4675
rect 9674 4672 9680 4684
rect 8895 4644 9680 4672
rect 8895 4641 8907 4644
rect 8849 4635 8907 4641
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 9953 4675 10011 4681
rect 9953 4641 9965 4675
rect 9999 4672 10011 4675
rect 10870 4672 10876 4684
rect 9999 4644 10876 4672
rect 9999 4641 10011 4644
rect 9953 4635 10011 4641
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 11072 4644 13124 4672
rect 11072 4616 11100 4644
rect 5307 4576 5580 4604
rect 7929 4607 7987 4613
rect 5307 4573 5319 4576
rect 5261 4567 5319 4573
rect 7929 4573 7941 4607
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 8386 4564 8392 4616
rect 8444 4604 8450 4616
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 8444 4576 8953 4604
rect 8444 4564 8450 4576
rect 8941 4573 8953 4576
rect 8987 4573 8999 4607
rect 11054 4604 11060 4616
rect 11015 4576 11060 4604
rect 8941 4567 8999 4573
rect 11054 4564 11060 4576
rect 11112 4564 11118 4616
rect 11977 4607 12035 4613
rect 11977 4573 11989 4607
rect 12023 4573 12035 4607
rect 12158 4604 12164 4616
rect 12119 4576 12164 4604
rect 11977 4567 12035 4573
rect 5626 4536 5632 4548
rect 5092 4508 5632 4536
rect 4617 4499 4675 4505
rect 5626 4496 5632 4508
rect 5684 4496 5690 4548
rect 7650 4496 7656 4548
rect 7708 4536 7714 4548
rect 8294 4536 8300 4548
rect 7708 4508 8300 4536
rect 7708 4496 7714 4508
rect 8294 4496 8300 4508
rect 8352 4496 8358 4548
rect 8846 4496 8852 4548
rect 8904 4536 8910 4548
rect 11422 4536 11428 4548
rect 8904 4508 11428 4536
rect 8904 4496 8910 4508
rect 11422 4496 11428 4508
rect 11480 4496 11486 4548
rect 11992 4536 12020 4567
rect 12158 4564 12164 4576
rect 12216 4564 12222 4616
rect 13096 4613 13124 4644
rect 14274 4632 14280 4684
rect 14332 4672 14338 4684
rect 14645 4675 14703 4681
rect 14645 4672 14657 4675
rect 14332 4644 14657 4672
rect 14332 4632 14338 4644
rect 14645 4641 14657 4644
rect 14691 4641 14703 4675
rect 14645 4635 14703 4641
rect 14734 4632 14740 4684
rect 14792 4672 14798 4684
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 14792 4644 15669 4672
rect 14792 4632 14798 4644
rect 15657 4641 15669 4644
rect 15703 4641 15715 4675
rect 15657 4635 15715 4641
rect 16206 4632 16212 4684
rect 16264 4672 16270 4684
rect 16761 4675 16819 4681
rect 16761 4672 16773 4675
rect 16264 4644 16773 4672
rect 16264 4632 16270 4644
rect 16761 4641 16773 4644
rect 16807 4641 16819 4675
rect 16868 4672 16896 4712
rect 17313 4709 17325 4712
rect 17359 4709 17371 4743
rect 17313 4703 17371 4709
rect 17865 4743 17923 4749
rect 17865 4709 17877 4743
rect 17911 4740 17923 4743
rect 18690 4740 18696 4752
rect 17911 4712 18696 4740
rect 17911 4709 17923 4712
rect 17865 4703 17923 4709
rect 18690 4700 18696 4712
rect 18748 4700 18754 4752
rect 18417 4675 18475 4681
rect 18417 4672 18429 4675
rect 16868 4644 18429 4672
rect 16761 4635 16819 4641
rect 18417 4641 18429 4644
rect 18463 4641 18475 4675
rect 18782 4672 18788 4684
rect 18417 4635 18475 4641
rect 18515 4644 18788 4672
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4604 13139 4607
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 13127 4576 14105 4604
rect 13127 4573 13139 4576
rect 13081 4567 13139 4573
rect 14093 4573 14105 4576
rect 14139 4604 14151 4607
rect 14182 4604 14188 4616
rect 14139 4576 14188 4604
rect 14139 4573 14151 4576
rect 14093 4567 14151 4573
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14458 4564 14464 4616
rect 14516 4604 14522 4616
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 14516 4576 15761 4604
rect 14516 4564 14522 4576
rect 15749 4573 15761 4576
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 15933 4607 15991 4613
rect 15933 4573 15945 4607
rect 15979 4604 15991 4607
rect 16022 4604 16028 4616
rect 15979 4576 16028 4604
rect 15979 4573 15991 4576
rect 15933 4567 15991 4573
rect 16022 4564 16028 4576
rect 16080 4564 16086 4616
rect 16850 4604 16856 4616
rect 16811 4576 16856 4604
rect 16850 4564 16856 4576
rect 16908 4564 16914 4616
rect 17034 4604 17040 4616
rect 16995 4576 17040 4604
rect 17034 4564 17040 4576
rect 17092 4564 17098 4616
rect 17313 4607 17371 4613
rect 17313 4573 17325 4607
rect 17359 4604 17371 4607
rect 17957 4607 18015 4613
rect 17957 4604 17969 4607
rect 17359 4576 17969 4604
rect 17359 4573 17371 4576
rect 17313 4567 17371 4573
rect 17957 4573 17969 4576
rect 18003 4573 18015 4607
rect 18515 4604 18543 4644
rect 18782 4632 18788 4644
rect 18840 4632 18846 4684
rect 19518 4672 19524 4684
rect 19479 4644 19524 4672
rect 19518 4632 19524 4644
rect 19576 4632 19582 4684
rect 19794 4632 19800 4684
rect 19852 4672 19858 4684
rect 20165 4675 20223 4681
rect 20165 4672 20177 4675
rect 19852 4644 20177 4672
rect 19852 4632 19858 4644
rect 20165 4641 20177 4644
rect 20211 4641 20223 4675
rect 20165 4635 20223 4641
rect 17957 4567 18015 4573
rect 18340 4576 18543 4604
rect 18693 4607 18751 4613
rect 13541 4539 13599 4545
rect 13541 4536 13553 4539
rect 11992 4508 13553 4536
rect 13541 4505 13553 4508
rect 13587 4505 13599 4539
rect 13541 4499 13599 4505
rect 15289 4539 15347 4545
rect 15289 4505 15301 4539
rect 15335 4536 15347 4539
rect 18340 4536 18368 4576
rect 18693 4573 18705 4607
rect 18739 4573 18751 4607
rect 19610 4604 19616 4616
rect 19571 4576 19616 4604
rect 18693 4567 18751 4573
rect 15335 4508 18368 4536
rect 18708 4536 18736 4567
rect 19610 4564 19616 4576
rect 19668 4564 19674 4616
rect 19702 4564 19708 4616
rect 19760 4604 19766 4616
rect 19760 4576 19805 4604
rect 19760 4564 19766 4576
rect 19886 4564 19892 4616
rect 19944 4604 19950 4616
rect 20901 4607 20959 4613
rect 20901 4604 20913 4607
rect 19944 4576 20913 4604
rect 19944 4564 19950 4576
rect 20901 4573 20913 4576
rect 20947 4573 20959 4607
rect 20901 4567 20959 4573
rect 20162 4536 20168 4548
rect 18708 4508 20168 4536
rect 15335 4505 15347 4508
rect 15289 4499 15347 4505
rect 20162 4496 20168 4508
rect 20220 4496 20226 4548
rect 2961 4471 3019 4477
rect 2961 4437 2973 4471
rect 3007 4468 3019 4471
rect 3970 4468 3976 4480
rect 3007 4440 3976 4468
rect 3007 4437 3019 4440
rect 2961 4431 3019 4437
rect 3970 4428 3976 4440
rect 4028 4428 4034 4480
rect 4249 4471 4307 4477
rect 4249 4437 4261 4471
rect 4295 4468 4307 4471
rect 10962 4468 10968 4480
rect 4295 4440 10968 4468
rect 4295 4437 4307 4440
rect 4249 4431 4307 4437
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 11517 4471 11575 4477
rect 11517 4437 11529 4471
rect 11563 4468 11575 4471
rect 11698 4468 11704 4480
rect 11563 4440 11704 4468
rect 11563 4437 11575 4440
rect 11517 4431 11575 4437
rect 11698 4428 11704 4440
rect 11756 4428 11762 4480
rect 12529 4471 12587 4477
rect 12529 4437 12541 4471
rect 12575 4468 12587 4471
rect 12894 4468 12900 4480
rect 12575 4440 12900 4468
rect 12575 4437 12587 4440
rect 12529 4431 12587 4437
rect 12894 4428 12900 4440
rect 12952 4428 12958 4480
rect 13078 4428 13084 4480
rect 13136 4468 13142 4480
rect 13357 4471 13415 4477
rect 13357 4468 13369 4471
rect 13136 4440 13369 4468
rect 13136 4428 13142 4440
rect 13357 4437 13369 4440
rect 13403 4437 13415 4471
rect 14826 4468 14832 4480
rect 14787 4440 14832 4468
rect 13357 4431 13415 4437
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 15102 4428 15108 4480
rect 15160 4468 15166 4480
rect 15654 4468 15660 4480
rect 15160 4440 15660 4468
rect 15160 4428 15166 4440
rect 15654 4428 15660 4440
rect 15712 4428 15718 4480
rect 16393 4471 16451 4477
rect 16393 4437 16405 4471
rect 16439 4468 16451 4471
rect 17310 4468 17316 4480
rect 16439 4440 17316 4468
rect 16439 4437 16451 4440
rect 16393 4431 16451 4437
rect 17310 4428 17316 4440
rect 17368 4428 17374 4480
rect 17402 4428 17408 4480
rect 17460 4468 17466 4480
rect 18233 4471 18291 4477
rect 18233 4468 18245 4471
rect 17460 4440 18245 4468
rect 17460 4428 17466 4440
rect 18233 4437 18245 4440
rect 18279 4437 18291 4471
rect 18233 4431 18291 4437
rect 19153 4471 19211 4477
rect 19153 4437 19165 4471
rect 19199 4468 19211 4471
rect 20070 4468 20076 4480
rect 19199 4440 20076 4468
rect 19199 4437 19211 4440
rect 19153 4431 19211 4437
rect 20070 4428 20076 4440
rect 20128 4428 20134 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 3602 4224 3608 4276
rect 3660 4264 3666 4276
rect 13722 4264 13728 4276
rect 3660 4236 13728 4264
rect 3660 4224 3666 4236
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 14645 4267 14703 4273
rect 14645 4233 14657 4267
rect 14691 4264 14703 4267
rect 14737 4267 14795 4273
rect 14737 4264 14749 4267
rect 14691 4236 14749 4264
rect 14691 4233 14703 4236
rect 14645 4227 14703 4233
rect 14737 4233 14749 4236
rect 14783 4233 14795 4267
rect 14737 4227 14795 4233
rect 14826 4224 14832 4276
rect 14884 4264 14890 4276
rect 17770 4264 17776 4276
rect 14884 4236 17776 4264
rect 14884 4224 14890 4236
rect 17770 4224 17776 4236
rect 17828 4224 17834 4276
rect 19705 4267 19763 4273
rect 17880 4236 19104 4264
rect 4709 4199 4767 4205
rect 4709 4165 4721 4199
rect 4755 4196 4767 4199
rect 5994 4196 6000 4208
rect 4755 4168 6000 4196
rect 4755 4165 4767 4168
rect 4709 4159 4767 4165
rect 5994 4156 6000 4168
rect 6052 4156 6058 4208
rect 6362 4156 6368 4208
rect 6420 4196 6426 4208
rect 6730 4196 6736 4208
rect 6420 4168 6736 4196
rect 6420 4156 6426 4168
rect 6730 4156 6736 4168
rect 6788 4156 6794 4208
rect 6825 4199 6883 4205
rect 6825 4165 6837 4199
rect 6871 4165 6883 4199
rect 8202 4196 8208 4208
rect 6825 4159 6883 4165
rect 7484 4168 8208 4196
rect 2222 4128 2228 4140
rect 2183 4100 2228 4128
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 3142 4128 3148 4140
rect 3103 4100 3148 4128
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 3326 4128 3332 4140
rect 3287 4100 3332 4128
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 5166 4128 5172 4140
rect 4295 4100 5172 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 5166 4088 5172 4100
rect 5224 4128 5230 4140
rect 5629 4131 5687 4137
rect 5629 4128 5641 4131
rect 5224 4100 5641 4128
rect 5224 4088 5230 4100
rect 5629 4097 5641 4100
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4060 2191 4063
rect 4338 4060 4344 4072
rect 2179 4032 4344 4060
rect 2179 4029 2191 4032
rect 2133 4023 2191 4029
rect 4338 4020 4344 4032
rect 4396 4020 4402 4072
rect 4525 4063 4583 4069
rect 4525 4029 4537 4063
rect 4571 4060 4583 4063
rect 5718 4060 5724 4072
rect 4571 4032 5724 4060
rect 4571 4029 4583 4032
rect 4525 4023 4583 4029
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 6181 4063 6239 4069
rect 6181 4029 6193 4063
rect 6227 4060 6239 4063
rect 6546 4060 6552 4072
rect 6227 4032 6552 4060
rect 6227 4029 6239 4032
rect 6181 4023 6239 4029
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 2041 3995 2099 4001
rect 2041 3961 2053 3995
rect 2087 3992 2099 3995
rect 3053 3995 3111 4001
rect 2087 3964 2728 3992
rect 2087 3961 2099 3964
rect 2041 3955 2099 3961
rect 1673 3927 1731 3933
rect 1673 3893 1685 3927
rect 1719 3924 1731 3927
rect 2406 3924 2412 3936
rect 1719 3896 2412 3924
rect 1719 3893 1731 3896
rect 1673 3887 1731 3893
rect 2406 3884 2412 3896
rect 2464 3884 2470 3936
rect 2700 3933 2728 3964
rect 3053 3961 3065 3995
rect 3099 3992 3111 3995
rect 4890 3992 4896 4004
rect 3099 3964 4896 3992
rect 3099 3961 3111 3964
rect 3053 3955 3111 3961
rect 4890 3952 4896 3964
rect 4948 3952 4954 4004
rect 5258 3952 5264 4004
rect 5316 3992 5322 4004
rect 5353 3995 5411 4001
rect 5353 3992 5365 3995
rect 5316 3964 5365 3992
rect 5316 3952 5322 3964
rect 5353 3961 5365 3964
rect 5399 3961 5411 3995
rect 5353 3955 5411 3961
rect 5445 3995 5503 4001
rect 5445 3961 5457 3995
rect 5491 3992 5503 3995
rect 5994 3992 6000 4004
rect 5491 3964 6000 3992
rect 5491 3961 5503 3964
rect 5445 3955 5503 3961
rect 5994 3952 6000 3964
rect 6052 3952 6058 4004
rect 6840 3992 6868 4159
rect 7006 4088 7012 4140
rect 7064 4128 7070 4140
rect 7484 4137 7512 4168
rect 8202 4156 8208 4168
rect 8260 4156 8266 4208
rect 8294 4156 8300 4208
rect 8352 4196 8358 4208
rect 8352 4168 8397 4196
rect 8352 4156 8358 4168
rect 9858 4156 9864 4208
rect 9916 4196 9922 4208
rect 10318 4196 10324 4208
rect 9916 4168 10324 4196
rect 9916 4156 9922 4168
rect 10318 4156 10324 4168
rect 10376 4156 10382 4208
rect 10520 4168 11836 4196
rect 7285 4131 7343 4137
rect 7285 4128 7297 4131
rect 7064 4100 7297 4128
rect 7064 4088 7070 4100
rect 7285 4097 7297 4100
rect 7331 4097 7343 4131
rect 7285 4091 7343 4097
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 7190 4060 7196 4072
rect 7151 4032 7196 4060
rect 7190 4020 7196 4032
rect 7248 4020 7254 4072
rect 7558 4020 7564 4072
rect 7616 4060 7622 4072
rect 8113 4063 8171 4069
rect 8113 4060 8125 4063
rect 7616 4032 8125 4060
rect 7616 4020 7622 4032
rect 8113 4029 8125 4032
rect 8159 4029 8171 4063
rect 8113 4023 8171 4029
rect 8202 4020 8208 4072
rect 8260 4060 8266 4072
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 8260 4032 8677 4060
rect 8260 4020 8266 4032
rect 8665 4029 8677 4032
rect 8711 4029 8723 4063
rect 10321 4063 10379 4069
rect 10321 4060 10333 4063
rect 8665 4023 8723 4029
rect 8763 4032 10333 4060
rect 8763 3992 8791 4032
rect 10321 4029 10333 4032
rect 10367 4029 10379 4063
rect 10321 4023 10379 4029
rect 6840 3964 8791 3992
rect 8932 3995 8990 4001
rect 8932 3961 8944 3995
rect 8978 3992 8990 3995
rect 10520 3992 10548 4168
rect 11698 4128 11704 4140
rect 11659 4100 11704 4128
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 11808 4137 11836 4168
rect 11882 4156 11888 4208
rect 11940 4196 11946 4208
rect 12437 4199 12495 4205
rect 11940 4168 12296 4196
rect 11940 4156 11946 4168
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4128 11851 4131
rect 12066 4128 12072 4140
rect 11839 4100 12072 4128
rect 11839 4097 11851 4100
rect 11793 4091 11851 4097
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12268 4128 12296 4168
rect 12437 4165 12449 4199
rect 12483 4196 12495 4199
rect 13078 4196 13084 4208
rect 12483 4168 13084 4196
rect 12483 4165 12495 4168
rect 12437 4159 12495 4165
rect 13078 4156 13084 4168
rect 13136 4156 13142 4208
rect 14182 4156 14188 4208
rect 14240 4196 14246 4208
rect 14461 4199 14519 4205
rect 14461 4196 14473 4199
rect 14240 4168 14473 4196
rect 14240 4156 14246 4168
rect 14461 4165 14473 4168
rect 14507 4165 14519 4199
rect 14461 4159 14519 4165
rect 14550 4156 14556 4208
rect 14608 4196 14614 4208
rect 14608 4168 15332 4196
rect 14608 4156 14614 4168
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12268 4100 13001 4128
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 14645 4131 14703 4137
rect 14645 4097 14657 4131
rect 14691 4128 14703 4131
rect 15194 4128 15200 4140
rect 14691 4100 15200 4128
rect 14691 4097 14703 4100
rect 14645 4091 14703 4097
rect 15194 4088 15200 4100
rect 15252 4088 15258 4140
rect 15304 4137 15332 4168
rect 17678 4156 17684 4208
rect 17736 4196 17742 4208
rect 17880 4196 17908 4236
rect 17736 4168 17908 4196
rect 17736 4156 17742 4168
rect 15289 4131 15347 4137
rect 15289 4097 15301 4131
rect 15335 4097 15347 4131
rect 15289 4091 15347 4097
rect 15672 4100 15884 4128
rect 10686 4020 10692 4072
rect 10744 4060 10750 4072
rect 11882 4060 11888 4072
rect 10744 4032 11888 4060
rect 10744 4020 10750 4032
rect 11882 4020 11888 4032
rect 11940 4020 11946 4072
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 12529 4063 12587 4069
rect 12529 4029 12541 4063
rect 12575 4060 12587 4063
rect 12802 4060 12808 4072
rect 12575 4032 12808 4060
rect 12575 4029 12587 4032
rect 12529 4023 12587 4029
rect 8978 3964 10548 3992
rect 8978 3961 8990 3964
rect 8932 3955 8990 3961
rect 10594 3952 10600 4004
rect 10652 3992 10658 4004
rect 12452 3992 12480 4023
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4060 13139 4063
rect 13170 4060 13176 4072
rect 13127 4032 13176 4060
rect 13127 4029 13139 4032
rect 13081 4023 13139 4029
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 15672 4060 15700 4100
rect 13280 4032 15700 4060
rect 15749 4063 15807 4069
rect 10652 3964 10697 3992
rect 10796 3964 12480 3992
rect 10652 3952 10658 3964
rect 2685 3927 2743 3933
rect 2685 3893 2697 3927
rect 2731 3893 2743 3927
rect 3694 3924 3700 3936
rect 3655 3896 3700 3924
rect 2685 3887 2743 3893
rect 3694 3884 3700 3896
rect 3752 3884 3758 3936
rect 3878 3884 3884 3936
rect 3936 3924 3942 3936
rect 4065 3927 4123 3933
rect 4065 3924 4077 3927
rect 3936 3896 4077 3924
rect 3936 3884 3942 3896
rect 4065 3893 4077 3896
rect 4111 3893 4123 3927
rect 4065 3887 4123 3893
rect 4154 3884 4160 3936
rect 4212 3924 4218 3936
rect 4798 3924 4804 3936
rect 4212 3896 4804 3924
rect 4212 3884 4218 3896
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 4982 3924 4988 3936
rect 4943 3896 4988 3924
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 6365 3927 6423 3933
rect 6365 3893 6377 3927
rect 6411 3924 6423 3927
rect 9858 3924 9864 3936
rect 6411 3896 9864 3924
rect 6411 3893 6423 3896
rect 6365 3887 6423 3893
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 10045 3927 10103 3933
rect 10045 3893 10057 3927
rect 10091 3924 10103 3927
rect 10226 3924 10232 3936
rect 10091 3896 10232 3924
rect 10091 3893 10103 3896
rect 10045 3887 10103 3893
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10318 3884 10324 3936
rect 10376 3924 10382 3936
rect 10796 3924 10824 3964
rect 12618 3952 12624 4004
rect 12676 3992 12682 4004
rect 13280 3992 13308 4032
rect 15749 4029 15761 4063
rect 15795 4029 15807 4063
rect 15856 4060 15884 4100
rect 16022 4088 16028 4140
rect 16080 4128 16086 4140
rect 16945 4131 17003 4137
rect 16945 4128 16957 4131
rect 16080 4100 16957 4128
rect 16080 4088 16086 4100
rect 16945 4097 16957 4100
rect 16991 4128 17003 4131
rect 17954 4128 17960 4140
rect 16991 4100 17960 4128
rect 16991 4097 17003 4100
rect 16945 4091 17003 4097
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 18046 4088 18052 4140
rect 18104 4128 18110 4140
rect 19076 4128 19104 4236
rect 19705 4233 19717 4267
rect 19751 4264 19763 4267
rect 20530 4264 20536 4276
rect 19751 4236 20536 4264
rect 19751 4233 19763 4236
rect 19705 4227 19763 4233
rect 20530 4224 20536 4236
rect 20588 4224 20594 4276
rect 20254 4156 20260 4208
rect 20312 4196 20318 4208
rect 20898 4196 20904 4208
rect 20312 4168 20392 4196
rect 20859 4168 20904 4196
rect 20312 4156 20318 4168
rect 19978 4128 19984 4140
rect 18104 4100 18149 4128
rect 19076 4100 19984 4128
rect 18104 4088 18110 4100
rect 19978 4088 19984 4100
rect 20036 4088 20042 4140
rect 20364 4137 20392 4168
rect 20898 4156 20904 4168
rect 20956 4156 20962 4208
rect 20349 4131 20407 4137
rect 20349 4097 20361 4131
rect 20395 4097 20407 4131
rect 20349 4091 20407 4097
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 15856 4032 17325 4060
rect 15749 4023 15807 4029
rect 17313 4029 17325 4032
rect 17359 4060 17371 4063
rect 17497 4063 17555 4069
rect 17497 4060 17509 4063
rect 17359 4032 17509 4060
rect 17359 4029 17371 4032
rect 17313 4023 17371 4029
rect 17497 4029 17509 4032
rect 17543 4029 17555 4063
rect 19794 4060 19800 4072
rect 17497 4023 17555 4029
rect 18156 4032 19800 4060
rect 13354 4001 13360 4004
rect 12676 3964 13308 3992
rect 12676 3952 12682 3964
rect 13348 3955 13360 4001
rect 13412 3992 13418 4004
rect 13412 3964 13448 3992
rect 13354 3952 13360 3955
rect 13412 3952 13418 3964
rect 14090 3952 14096 4004
rect 14148 3992 14154 4004
rect 15764 3992 15792 4023
rect 14148 3964 15792 3992
rect 16025 3995 16083 4001
rect 14148 3952 14154 3964
rect 16025 3961 16037 3995
rect 16071 3992 16083 3995
rect 18156 3992 18184 4032
rect 19794 4020 19800 4032
rect 19852 4020 19858 4072
rect 20165 4063 20223 4069
rect 20165 4029 20177 4063
rect 20211 4060 20223 4063
rect 20530 4060 20536 4072
rect 20211 4032 20536 4060
rect 20211 4029 20223 4032
rect 20165 4023 20223 4029
rect 20530 4020 20536 4032
rect 20588 4020 20594 4072
rect 20717 4063 20775 4069
rect 20717 4029 20729 4063
rect 20763 4029 20775 4063
rect 20717 4023 20775 4029
rect 16071 3964 18184 3992
rect 18294 3995 18352 4001
rect 16071 3961 16083 3964
rect 16025 3955 16083 3961
rect 18294 3961 18306 3995
rect 18340 3961 18352 3995
rect 18294 3955 18352 3961
rect 10376 3896 10824 3924
rect 11241 3927 11299 3933
rect 10376 3884 10382 3896
rect 11241 3893 11253 3927
rect 11287 3924 11299 3927
rect 11514 3924 11520 3936
rect 11287 3896 11520 3924
rect 11287 3893 11299 3896
rect 11241 3887 11299 3893
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 11609 3927 11667 3933
rect 11609 3893 11621 3927
rect 11655 3924 11667 3927
rect 12434 3924 12440 3936
rect 11655 3896 12440 3924
rect 11655 3893 11667 3896
rect 11609 3887 11667 3893
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 12713 3927 12771 3933
rect 12713 3893 12725 3927
rect 12759 3924 12771 3927
rect 12802 3924 12808 3936
rect 12759 3896 12808 3924
rect 12759 3893 12771 3896
rect 12713 3887 12771 3893
rect 12802 3884 12808 3896
rect 12860 3884 12866 3936
rect 12989 3927 13047 3933
rect 12989 3893 13001 3927
rect 13035 3924 13047 3927
rect 13998 3924 14004 3936
rect 13035 3896 14004 3924
rect 13035 3893 13047 3896
rect 12989 3887 13047 3893
rect 13998 3884 14004 3896
rect 14056 3884 14062 3936
rect 15102 3924 15108 3936
rect 15063 3896 15108 3924
rect 15102 3884 15108 3896
rect 15160 3884 15166 3936
rect 15194 3884 15200 3936
rect 15252 3924 15258 3936
rect 15252 3896 15297 3924
rect 15252 3884 15258 3896
rect 16298 3884 16304 3936
rect 16356 3924 16362 3936
rect 16666 3924 16672 3936
rect 16356 3896 16401 3924
rect 16627 3896 16672 3924
rect 16356 3884 16362 3896
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 16761 3927 16819 3933
rect 16761 3893 16773 3927
rect 16807 3924 16819 3927
rect 16942 3924 16948 3936
rect 16807 3896 16948 3924
rect 16807 3893 16819 3896
rect 16761 3887 16819 3893
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 17034 3884 17040 3936
rect 17092 3924 17098 3936
rect 18309 3924 18337 3955
rect 20346 3952 20352 4004
rect 20404 3992 20410 4004
rect 20732 3992 20760 4023
rect 20404 3964 20760 3992
rect 20404 3952 20410 3964
rect 19334 3924 19340 3936
rect 17092 3896 19340 3924
rect 17092 3884 17098 3896
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 19429 3927 19487 3933
rect 19429 3893 19441 3927
rect 19475 3924 19487 3927
rect 19702 3924 19708 3936
rect 19475 3896 19708 3924
rect 19475 3893 19487 3896
rect 19429 3887 19487 3893
rect 19702 3884 19708 3896
rect 19760 3924 19766 3936
rect 19978 3924 19984 3936
rect 19760 3896 19984 3924
rect 19760 3884 19766 3896
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 20070 3884 20076 3936
rect 20128 3924 20134 3936
rect 20128 3896 20173 3924
rect 20128 3884 20134 3896
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 2038 3720 2044 3732
rect 1412 3692 2044 3720
rect 1412 3593 1440 3692
rect 2038 3680 2044 3692
rect 2096 3680 2102 3732
rect 2222 3680 2228 3732
rect 2280 3720 2286 3732
rect 3513 3723 3571 3729
rect 3513 3720 3525 3723
rect 2280 3692 3525 3720
rect 2280 3680 2286 3692
rect 3513 3689 3525 3692
rect 3559 3689 3571 3723
rect 3513 3683 3571 3689
rect 3602 3680 3608 3732
rect 3660 3720 3666 3732
rect 3878 3720 3884 3732
rect 3660 3692 3884 3720
rect 3660 3680 3666 3692
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 4801 3723 4859 3729
rect 4801 3720 4813 3723
rect 4304 3692 4813 3720
rect 4304 3680 4310 3692
rect 4801 3689 4813 3692
rect 4847 3689 4859 3723
rect 4801 3683 4859 3689
rect 4982 3680 4988 3732
rect 5040 3720 5046 3732
rect 5813 3723 5871 3729
rect 5813 3720 5825 3723
rect 5040 3692 5825 3720
rect 5040 3680 5046 3692
rect 5813 3689 5825 3692
rect 5859 3689 5871 3723
rect 7006 3720 7012 3732
rect 6967 3692 7012 3720
rect 5813 3683 5871 3689
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 7653 3723 7711 3729
rect 7653 3689 7665 3723
rect 7699 3720 7711 3723
rect 9674 3720 9680 3732
rect 7699 3692 9076 3720
rect 9635 3692 9680 3720
rect 7699 3689 7711 3692
rect 7653 3683 7711 3689
rect 1670 3652 1676 3664
rect 1631 3624 1676 3652
rect 1670 3612 1676 3624
rect 1728 3612 1734 3664
rect 7098 3652 7104 3664
rect 3620 3624 6684 3652
rect 7011 3624 7104 3652
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 1854 3544 1860 3596
rect 1912 3584 1918 3596
rect 2133 3587 2191 3593
rect 2133 3584 2145 3587
rect 1912 3556 2145 3584
rect 1912 3544 1918 3556
rect 2133 3553 2145 3556
rect 2179 3553 2191 3587
rect 2133 3547 2191 3553
rect 2400 3587 2458 3593
rect 2400 3553 2412 3587
rect 2446 3584 2458 3587
rect 3326 3584 3332 3596
rect 2446 3556 3332 3584
rect 2446 3553 2458 3556
rect 2400 3547 2458 3553
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 3620 3593 3648 3624
rect 3605 3587 3663 3593
rect 3605 3553 3617 3587
rect 3651 3553 3663 3587
rect 3605 3547 3663 3553
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 4893 3587 4951 3593
rect 4893 3584 4905 3587
rect 4212 3556 4905 3584
rect 4212 3544 4218 3556
rect 4893 3553 4905 3556
rect 4939 3553 4951 3587
rect 6362 3584 6368 3596
rect 4893 3547 4951 3553
rect 5000 3556 6368 3584
rect 5000 3516 5028 3556
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 3804 3488 5028 3516
rect 5077 3519 5135 3525
rect 3804 3457 3832 3488
rect 5077 3485 5089 3519
rect 5123 3516 5135 3519
rect 5166 3516 5172 3528
rect 5123 3488 5172 3516
rect 5123 3485 5135 3488
rect 5077 3479 5135 3485
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 3789 3451 3847 3457
rect 3789 3417 3801 3451
rect 3835 3417 3847 3451
rect 3789 3411 3847 3417
rect 4154 3408 4160 3460
rect 4212 3448 4218 3460
rect 4249 3451 4307 3457
rect 4249 3448 4261 3451
rect 4212 3420 4261 3448
rect 4212 3408 4218 3420
rect 4249 3417 4261 3420
rect 4295 3417 4307 3451
rect 4249 3411 4307 3417
rect 4433 3451 4491 3457
rect 4433 3417 4445 3451
rect 4479 3448 4491 3451
rect 5920 3448 5948 3479
rect 5994 3476 6000 3528
rect 6052 3516 6058 3528
rect 6052 3488 6097 3516
rect 6052 3476 6058 3488
rect 4479 3420 5948 3448
rect 6656 3448 6684 3624
rect 7098 3612 7104 3624
rect 7156 3652 7162 3664
rect 7282 3652 7288 3664
rect 7156 3624 7288 3652
rect 7156 3612 7162 3624
rect 7282 3612 7288 3624
rect 7340 3612 7346 3664
rect 7374 3612 7380 3664
rect 7432 3652 7438 3664
rect 7432 3624 7972 3652
rect 7432 3612 7438 3624
rect 7944 3584 7972 3624
rect 8018 3612 8024 3664
rect 8076 3652 8082 3664
rect 8938 3652 8944 3664
rect 8076 3624 8944 3652
rect 8076 3612 8082 3624
rect 8938 3612 8944 3624
rect 8996 3612 9002 3664
rect 8113 3587 8171 3593
rect 8113 3584 8125 3587
rect 7944 3556 8125 3584
rect 8113 3553 8125 3556
rect 8159 3553 8171 3587
rect 8113 3547 8171 3553
rect 8478 3544 8484 3596
rect 8536 3584 8542 3596
rect 8849 3587 8907 3593
rect 8849 3584 8861 3587
rect 8536 3556 8861 3584
rect 8536 3544 8542 3556
rect 8849 3553 8861 3556
rect 8895 3553 8907 3587
rect 9048 3584 9076 3692
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 9766 3680 9772 3732
rect 9824 3720 9830 3732
rect 10137 3723 10195 3729
rect 9824 3692 10088 3720
rect 9824 3680 9830 3692
rect 9125 3655 9183 3661
rect 9125 3621 9137 3655
rect 9171 3652 9183 3655
rect 9950 3652 9956 3664
rect 9171 3624 9956 3652
rect 9171 3621 9183 3624
rect 9125 3615 9183 3621
rect 9950 3612 9956 3624
rect 10008 3612 10014 3664
rect 10060 3661 10088 3692
rect 10137 3689 10149 3723
rect 10183 3720 10195 3723
rect 10686 3720 10692 3732
rect 10183 3692 10692 3720
rect 10183 3689 10195 3692
rect 10137 3683 10195 3689
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 12434 3720 12440 3732
rect 12395 3692 12440 3720
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 12805 3723 12863 3729
rect 12805 3689 12817 3723
rect 12851 3720 12863 3723
rect 13449 3723 13507 3729
rect 13449 3720 13461 3723
rect 12851 3692 13461 3720
rect 12851 3689 12863 3692
rect 12805 3683 12863 3689
rect 13449 3689 13461 3692
rect 13495 3689 13507 3723
rect 13449 3683 13507 3689
rect 15289 3723 15347 3729
rect 15289 3689 15301 3723
rect 15335 3689 15347 3723
rect 15289 3683 15347 3689
rect 17037 3723 17095 3729
rect 17037 3689 17049 3723
rect 17083 3720 17095 3723
rect 18046 3720 18052 3732
rect 17083 3692 18052 3720
rect 17083 3689 17095 3692
rect 17037 3683 17095 3689
rect 11054 3661 11060 3664
rect 10045 3655 10103 3661
rect 10045 3621 10057 3655
rect 10091 3652 10103 3655
rect 10091 3624 10824 3652
rect 10091 3621 10103 3624
rect 10045 3615 10103 3621
rect 10796 3584 10824 3624
rect 11048 3615 11060 3661
rect 11112 3652 11118 3664
rect 11112 3624 11148 3652
rect 11054 3612 11060 3615
rect 11112 3612 11118 3624
rect 11238 3612 11244 3664
rect 11296 3652 11302 3664
rect 11296 3624 12848 3652
rect 11296 3612 11302 3624
rect 12820 3584 12848 3624
rect 12894 3612 12900 3664
rect 12952 3652 12958 3664
rect 15102 3652 15108 3664
rect 12952 3624 12997 3652
rect 13280 3624 15108 3652
rect 12952 3612 12958 3624
rect 13170 3584 13176 3596
rect 9048 3556 9996 3584
rect 10796 3556 12747 3584
rect 12820 3556 13176 3584
rect 8849 3547 8907 3553
rect 9968 3528 9996 3556
rect 7285 3519 7343 3525
rect 7285 3485 7297 3519
rect 7331 3516 7343 3519
rect 8297 3519 8355 3525
rect 8297 3516 8309 3519
rect 7331 3488 8309 3516
rect 7331 3485 7343 3488
rect 7285 3479 7343 3485
rect 8297 3485 8309 3488
rect 8343 3516 8355 3519
rect 8386 3516 8392 3528
rect 8343 3488 8392 3516
rect 8343 3485 8355 3488
rect 8297 3479 8355 3485
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 8570 3476 8576 3528
rect 8628 3516 8634 3528
rect 9766 3516 9772 3528
rect 8628 3488 9772 3516
rect 8628 3476 8634 3488
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 9950 3476 9956 3528
rect 10008 3476 10014 3528
rect 10226 3516 10232 3528
rect 10187 3488 10232 3516
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10686 3476 10692 3528
rect 10744 3516 10750 3528
rect 10781 3519 10839 3525
rect 10781 3516 10793 3519
rect 10744 3488 10793 3516
rect 10744 3476 10750 3488
rect 10781 3485 10793 3488
rect 10827 3485 10839 3519
rect 10781 3479 10839 3485
rect 10594 3448 10600 3460
rect 6656 3420 10600 3448
rect 4479 3417 4491 3420
rect 4433 3411 4491 3417
rect 4264 3380 4292 3411
rect 10594 3408 10600 3420
rect 10652 3408 10658 3460
rect 12719 3448 12747 3556
rect 13170 3544 13176 3556
rect 13228 3544 13234 3596
rect 12802 3476 12808 3528
rect 12860 3516 12866 3528
rect 12989 3519 13047 3525
rect 12989 3516 13001 3519
rect 12860 3488 13001 3516
rect 12860 3476 12866 3488
rect 12989 3485 13001 3488
rect 13035 3485 13047 3519
rect 12989 3479 13047 3485
rect 13280 3448 13308 3624
rect 15102 3612 15108 3624
rect 15160 3612 15166 3664
rect 15304 3652 15332 3683
rect 18046 3680 18052 3692
rect 18104 3680 18110 3732
rect 18509 3723 18567 3729
rect 18509 3689 18521 3723
rect 18555 3689 18567 3723
rect 18509 3683 18567 3689
rect 16850 3652 16856 3664
rect 15304 3624 16856 3652
rect 16850 3612 16856 3624
rect 16908 3612 16914 3664
rect 17396 3655 17454 3661
rect 17396 3621 17408 3655
rect 17442 3652 17454 3655
rect 17586 3652 17592 3664
rect 17442 3624 17592 3652
rect 17442 3621 17454 3624
rect 17396 3615 17454 3621
rect 17586 3612 17592 3624
rect 17644 3612 17650 3664
rect 17954 3612 17960 3664
rect 18012 3652 18018 3664
rect 18524 3652 18552 3683
rect 18690 3652 18696 3664
rect 18012 3624 18696 3652
rect 18012 3612 18018 3624
rect 18690 3612 18696 3624
rect 18748 3612 18754 3664
rect 19242 3612 19248 3664
rect 19300 3612 19306 3664
rect 20257 3655 20315 3661
rect 20257 3621 20269 3655
rect 20303 3652 20315 3655
rect 20346 3652 20352 3664
rect 20303 3624 20352 3652
rect 20303 3621 20315 3624
rect 20257 3615 20315 3621
rect 20346 3612 20352 3624
rect 20404 3612 20410 3664
rect 13817 3587 13875 3593
rect 13817 3553 13829 3587
rect 13863 3584 13875 3587
rect 14090 3584 14096 3596
rect 13863 3556 14096 3584
rect 13863 3553 13875 3556
rect 13817 3547 13875 3553
rect 14090 3544 14096 3556
rect 14148 3544 14154 3596
rect 14826 3584 14832 3596
rect 14787 3556 14832 3584
rect 14826 3544 14832 3556
rect 14884 3544 14890 3596
rect 15286 3544 15292 3596
rect 15344 3584 15350 3596
rect 15657 3587 15715 3593
rect 15657 3584 15669 3587
rect 15344 3556 15669 3584
rect 15344 3544 15350 3556
rect 15657 3553 15669 3556
rect 15703 3553 15715 3587
rect 15657 3547 15715 3553
rect 16393 3587 16451 3593
rect 16393 3553 16405 3587
rect 16439 3584 16451 3587
rect 16574 3584 16580 3596
rect 16439 3556 16580 3584
rect 16439 3553 16451 3556
rect 16393 3547 16451 3553
rect 16574 3544 16580 3556
rect 16632 3544 16638 3596
rect 16669 3587 16727 3593
rect 16669 3553 16681 3587
rect 16715 3584 16727 3587
rect 16715 3556 18184 3584
rect 16715 3553 16727 3556
rect 16669 3547 16727 3553
rect 13906 3516 13912 3528
rect 13819 3488 13912 3516
rect 13906 3476 13912 3488
rect 13964 3476 13970 3528
rect 14001 3519 14059 3525
rect 14001 3485 14013 3519
rect 14047 3516 14059 3519
rect 14182 3516 14188 3528
rect 14047 3488 14188 3516
rect 14047 3485 14059 3488
rect 14001 3479 14059 3485
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 14844 3516 14872 3544
rect 15749 3519 15807 3525
rect 15749 3516 15761 3519
rect 14844 3488 15761 3516
rect 15749 3485 15761 3488
rect 15795 3485 15807 3519
rect 15749 3479 15807 3485
rect 15933 3519 15991 3525
rect 15933 3485 15945 3519
rect 15979 3516 15991 3519
rect 16022 3516 16028 3528
rect 15979 3488 16028 3516
rect 15979 3485 15991 3488
rect 15933 3479 15991 3485
rect 11716 3420 12664 3448
rect 12719 3420 13308 3448
rect 13924 3448 13952 3476
rect 15764 3448 15792 3479
rect 16022 3476 16028 3488
rect 16080 3476 16086 3528
rect 16482 3476 16488 3528
rect 16540 3516 16546 3528
rect 17037 3519 17095 3525
rect 17037 3516 17049 3519
rect 16540 3488 17049 3516
rect 16540 3476 16546 3488
rect 17037 3485 17049 3488
rect 17083 3516 17095 3519
rect 17129 3519 17187 3525
rect 17129 3516 17141 3519
rect 17083 3488 17141 3516
rect 17083 3485 17095 3488
rect 17037 3479 17095 3485
rect 17129 3485 17141 3488
rect 17175 3485 17187 3519
rect 18156 3516 18184 3556
rect 18230 3544 18236 3596
rect 18288 3584 18294 3596
rect 18966 3584 18972 3596
rect 18288 3556 18972 3584
rect 18288 3544 18294 3556
rect 18966 3544 18972 3556
rect 19024 3544 19030 3596
rect 19153 3587 19211 3593
rect 19153 3584 19165 3587
rect 19076 3556 19165 3584
rect 18782 3516 18788 3528
rect 18156 3488 18788 3516
rect 17129 3479 17187 3485
rect 18782 3476 18788 3488
rect 18840 3476 18846 3528
rect 18874 3476 18880 3528
rect 18932 3516 18938 3528
rect 19076 3516 19104 3556
rect 19153 3553 19165 3556
rect 19199 3553 19211 3587
rect 19260 3584 19288 3612
rect 20165 3587 20223 3593
rect 20165 3584 20177 3587
rect 19260 3556 20177 3584
rect 19153 3547 19211 3553
rect 20165 3553 20177 3556
rect 20211 3553 20223 3587
rect 20165 3547 20223 3553
rect 19242 3516 19248 3528
rect 18932 3488 19104 3516
rect 19203 3488 19248 3516
rect 18932 3476 18938 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 20070 3516 20076 3528
rect 19392 3488 20076 3516
rect 19392 3476 19398 3488
rect 20070 3476 20076 3488
rect 20128 3516 20134 3528
rect 20349 3519 20407 3525
rect 20349 3516 20361 3519
rect 20128 3488 20361 3516
rect 20128 3476 20134 3488
rect 20349 3485 20361 3488
rect 20395 3485 20407 3519
rect 20349 3479 20407 3485
rect 16117 3451 16175 3457
rect 16117 3448 16129 3451
rect 13924 3420 14688 3448
rect 15764 3420 16129 3448
rect 5258 3380 5264 3392
rect 4264 3352 5264 3380
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 5442 3380 5448 3392
rect 5403 3352 5448 3380
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 6086 3340 6092 3392
rect 6144 3380 6150 3392
rect 6641 3383 6699 3389
rect 6641 3380 6653 3383
rect 6144 3352 6653 3380
rect 6144 3340 6150 3352
rect 6641 3349 6653 3352
rect 6687 3349 6699 3383
rect 6641 3343 6699 3349
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 7650 3380 7656 3392
rect 6972 3352 7656 3380
rect 6972 3340 6978 3352
rect 7650 3340 7656 3352
rect 7708 3340 7714 3392
rect 8294 3340 8300 3392
rect 8352 3380 8358 3392
rect 11716 3380 11744 3420
rect 12158 3380 12164 3392
rect 8352 3352 11744 3380
rect 12119 3352 12164 3380
rect 8352 3340 8358 3352
rect 12158 3340 12164 3352
rect 12216 3340 12222 3392
rect 12636 3380 12664 3420
rect 14550 3380 14556 3392
rect 12636 3352 14556 3380
rect 14550 3340 14556 3352
rect 14608 3340 14614 3392
rect 14660 3380 14688 3420
rect 16117 3417 16129 3420
rect 16163 3417 16175 3451
rect 16117 3411 16175 3417
rect 19610 3408 19616 3460
rect 19668 3448 19674 3460
rect 19797 3451 19855 3457
rect 19797 3448 19809 3451
rect 19668 3420 19809 3448
rect 19668 3408 19674 3420
rect 19797 3417 19809 3420
rect 19843 3417 19855 3451
rect 19797 3411 19855 3417
rect 17862 3380 17868 3392
rect 14660 3352 17868 3380
rect 17862 3340 17868 3352
rect 17920 3340 17926 3392
rect 18785 3383 18843 3389
rect 18785 3349 18797 3383
rect 18831 3380 18843 3383
rect 19702 3380 19708 3392
rect 18831 3352 19708 3380
rect 18831 3349 18843 3352
rect 18785 3343 18843 3349
rect 19702 3340 19708 3352
rect 19760 3340 19766 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 1854 3136 1860 3188
rect 1912 3176 1918 3188
rect 5721 3179 5779 3185
rect 1912 3148 3832 3176
rect 1912 3136 1918 3148
rect 1673 3111 1731 3117
rect 1673 3077 1685 3111
rect 1719 3108 1731 3111
rect 2314 3108 2320 3120
rect 1719 3080 2320 3108
rect 1719 3077 1731 3080
rect 1673 3071 1731 3077
rect 2314 3068 2320 3080
rect 2372 3068 2378 3120
rect 3694 3108 3700 3120
rect 3160 3080 3700 3108
rect 2222 3040 2228 3052
rect 2183 3012 2228 3040
rect 2222 3000 2228 3012
rect 2280 3000 2286 3052
rect 3160 3049 3188 3080
rect 3694 3068 3700 3080
rect 3752 3068 3758 3120
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3009 3203 3043
rect 3326 3040 3332 3052
rect 3287 3012 3332 3040
rect 3145 3003 3203 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 3804 3040 3832 3148
rect 5721 3145 5733 3179
rect 5767 3176 5779 3179
rect 6178 3176 6184 3188
rect 5767 3148 6184 3176
rect 5767 3145 5779 3148
rect 5721 3139 5779 3145
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 6270 3136 6276 3188
rect 6328 3176 6334 3188
rect 8202 3176 8208 3188
rect 6328 3148 8208 3176
rect 6328 3136 6334 3148
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 8846 3136 8852 3188
rect 8904 3176 8910 3188
rect 14001 3179 14059 3185
rect 8904 3148 13676 3176
rect 8904 3136 8910 3148
rect 5258 3108 5264 3120
rect 5171 3080 5264 3108
rect 5258 3068 5264 3080
rect 5316 3108 5322 3120
rect 5994 3108 6000 3120
rect 5316 3080 6000 3108
rect 5316 3068 5322 3080
rect 5994 3068 6000 3080
rect 6052 3068 6058 3120
rect 9950 3068 9956 3120
rect 10008 3108 10014 3120
rect 10502 3108 10508 3120
rect 10008 3080 10508 3108
rect 10008 3068 10014 3080
rect 10502 3068 10508 3080
rect 10560 3068 10566 3120
rect 12066 3108 12072 3120
rect 12027 3080 12072 3108
rect 12066 3068 12072 3080
rect 12124 3068 12130 3120
rect 12434 3108 12440 3120
rect 12395 3080 12440 3108
rect 12434 3068 12440 3080
rect 12492 3068 12498 3120
rect 3881 3043 3939 3049
rect 3881 3040 3893 3043
rect 3804 3012 3893 3040
rect 3881 3009 3893 3012
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2972 3571 2975
rect 3786 2972 3792 2984
rect 3559 2944 3792 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 3786 2932 3792 2944
rect 3844 2932 3850 2984
rect 3896 2972 3924 3003
rect 6270 3000 6276 3052
rect 6328 3040 6334 3052
rect 6328 3012 6373 3040
rect 6328 3000 6334 3012
rect 7834 3000 7840 3052
rect 7892 3040 7898 3052
rect 8110 3040 8116 3052
rect 7892 3012 8116 3040
rect 7892 3000 7898 3012
rect 8110 3000 8116 3012
rect 8168 3040 8174 3052
rect 8481 3043 8539 3049
rect 8481 3040 8493 3043
rect 8168 3012 8493 3040
rect 8168 3000 8174 3012
rect 8481 3009 8493 3012
rect 8527 3009 8539 3043
rect 10226 3040 10232 3052
rect 8481 3003 8539 3009
rect 10060 3012 10232 3040
rect 4430 2972 4436 2984
rect 3896 2944 4436 2972
rect 4430 2932 4436 2944
rect 4488 2932 4494 2984
rect 5350 2972 5356 2984
rect 5311 2944 5356 2972
rect 5350 2932 5356 2944
rect 5408 2932 5414 2984
rect 6086 2972 6092 2984
rect 6047 2944 6092 2972
rect 6086 2932 6092 2944
rect 6144 2932 6150 2984
rect 6822 2972 6828 2984
rect 6783 2944 6828 2972
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 8748 2975 8806 2981
rect 7024 2944 8432 2972
rect 4148 2907 4206 2913
rect 4148 2873 4160 2907
rect 4194 2904 4206 2907
rect 5166 2904 5172 2916
rect 4194 2876 5172 2904
rect 4194 2873 4206 2876
rect 4148 2867 4206 2873
rect 5166 2864 5172 2876
rect 5224 2864 5230 2916
rect 7024 2904 7052 2944
rect 5552 2876 7052 2904
rect 7092 2907 7150 2913
rect 2038 2836 2044 2848
rect 1999 2808 2044 2836
rect 2038 2796 2044 2808
rect 2096 2796 2102 2848
rect 2133 2839 2191 2845
rect 2133 2805 2145 2839
rect 2179 2836 2191 2839
rect 2685 2839 2743 2845
rect 2685 2836 2697 2839
rect 2179 2808 2697 2836
rect 2179 2805 2191 2808
rect 2133 2799 2191 2805
rect 2685 2805 2697 2808
rect 2731 2805 2743 2839
rect 3050 2836 3056 2848
rect 3011 2808 3056 2836
rect 2685 2799 2743 2805
rect 3050 2796 3056 2808
rect 3108 2796 3114 2848
rect 3694 2836 3700 2848
rect 3655 2808 3700 2836
rect 3694 2796 3700 2808
rect 3752 2796 3758 2848
rect 5552 2845 5580 2876
rect 7092 2873 7104 2907
rect 7138 2904 7150 2907
rect 8404 2904 8432 2944
rect 8748 2941 8760 2975
rect 8794 2972 8806 2975
rect 10060 2972 10088 3012
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 10686 3040 10692 3052
rect 10647 3012 10692 3040
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 12897 3043 12955 3049
rect 12897 3040 12909 3043
rect 11848 3012 12909 3040
rect 11848 3000 11854 3012
rect 12897 3009 12909 3012
rect 12943 3009 12955 3043
rect 13078 3040 13084 3052
rect 13039 3012 13084 3040
rect 12897 3003 12955 3009
rect 13078 3000 13084 3012
rect 13136 3000 13142 3052
rect 13648 3049 13676 3148
rect 14001 3145 14013 3179
rect 14047 3176 14059 3179
rect 14047 3148 16896 3176
rect 14047 3145 14059 3148
rect 14001 3139 14059 3145
rect 14274 3068 14280 3120
rect 14332 3108 14338 3120
rect 14332 3080 15240 3108
rect 14332 3068 14338 3080
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3009 13691 3043
rect 14090 3040 14096 3052
rect 14051 3012 14096 3040
rect 13633 3003 13691 3009
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 14918 3040 14924 3052
rect 14879 3012 14924 3040
rect 14918 3000 14924 3012
rect 14976 3000 14982 3052
rect 8794 2944 10088 2972
rect 10137 2975 10195 2981
rect 8794 2941 8806 2944
rect 8748 2935 8806 2941
rect 10137 2941 10149 2975
rect 10183 2972 10195 2975
rect 10318 2972 10324 2984
rect 10183 2944 10324 2972
rect 10183 2941 10195 2944
rect 10137 2935 10195 2941
rect 10318 2932 10324 2944
rect 10376 2932 10382 2984
rect 10956 2975 11014 2981
rect 10956 2941 10968 2975
rect 11002 2972 11014 2975
rect 12158 2972 12164 2984
rect 11002 2944 12164 2972
rect 11002 2941 11014 2944
rect 10956 2935 11014 2941
rect 12158 2932 12164 2944
rect 12216 2972 12222 2984
rect 12710 2972 12716 2984
rect 12216 2944 12716 2972
rect 12216 2932 12222 2944
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 12802 2932 12808 2984
rect 12860 2972 12866 2984
rect 13446 2972 13452 2984
rect 12860 2944 12905 2972
rect 13407 2944 13452 2972
rect 12860 2932 12866 2944
rect 13446 2932 13452 2944
rect 13504 2932 13510 2984
rect 15212 2981 15240 3080
rect 16868 3040 16896 3148
rect 17034 3136 17040 3188
rect 17092 3176 17098 3188
rect 17221 3179 17279 3185
rect 17221 3176 17233 3179
rect 17092 3148 17233 3176
rect 17092 3136 17098 3148
rect 17221 3145 17233 3148
rect 17267 3145 17279 3179
rect 17221 3139 17279 3145
rect 18141 3179 18199 3185
rect 18141 3145 18153 3179
rect 18187 3176 18199 3179
rect 18233 3179 18291 3185
rect 18233 3176 18245 3179
rect 18187 3148 18245 3176
rect 18187 3145 18199 3148
rect 18141 3139 18199 3145
rect 18233 3145 18245 3148
rect 18279 3145 18291 3179
rect 19518 3176 19524 3188
rect 18233 3139 18291 3145
rect 18616 3148 18920 3176
rect 19479 3148 19524 3176
rect 16942 3068 16948 3120
rect 17000 3108 17006 3120
rect 17678 3108 17684 3120
rect 17000 3080 17684 3108
rect 17000 3068 17006 3080
rect 17678 3068 17684 3080
rect 17736 3068 17742 3120
rect 17862 3068 17868 3120
rect 17920 3108 17926 3120
rect 18616 3108 18644 3148
rect 17920 3080 18644 3108
rect 18892 3108 18920 3148
rect 19518 3136 19524 3148
rect 19576 3136 19582 3188
rect 18892 3080 20024 3108
rect 17920 3068 17926 3080
rect 17218 3040 17224 3052
rect 16868 3012 17224 3040
rect 17218 3000 17224 3012
rect 17276 3000 17282 3052
rect 18141 3043 18199 3049
rect 18141 3009 18153 3043
rect 18187 3040 18199 3043
rect 18187 3012 18644 3040
rect 18187 3009 18199 3012
rect 18141 3003 18199 3009
rect 15197 2975 15255 2981
rect 15197 2941 15209 2975
rect 15243 2941 15255 2975
rect 15197 2935 15255 2941
rect 15841 2975 15899 2981
rect 15841 2941 15853 2975
rect 15887 2972 15899 2975
rect 16482 2972 16488 2984
rect 15887 2944 16488 2972
rect 15887 2941 15899 2944
rect 15841 2935 15899 2941
rect 16482 2932 16488 2944
rect 16540 2932 16546 2984
rect 18616 2972 18644 3012
rect 18690 3000 18696 3052
rect 18748 3040 18754 3052
rect 18785 3043 18843 3049
rect 18785 3040 18797 3043
rect 18748 3012 18797 3040
rect 18748 3000 18754 3012
rect 18785 3009 18797 3012
rect 18831 3009 18843 3043
rect 19242 3040 19248 3052
rect 18785 3003 18843 3009
rect 18892 3012 19248 3040
rect 18892 2972 18920 3012
rect 19242 3000 19248 3012
rect 19300 3000 19306 3052
rect 19996 3049 20024 3080
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3009 20039 3043
rect 19981 3003 20039 3009
rect 20070 3000 20076 3052
rect 20128 3040 20134 3052
rect 20128 3012 20173 3040
rect 20128 3000 20134 3012
rect 19886 2972 19892 2984
rect 18616 2944 18920 2972
rect 19847 2944 19892 2972
rect 19886 2932 19892 2944
rect 19944 2932 19950 2984
rect 20533 2975 20591 2981
rect 20533 2941 20545 2975
rect 20579 2941 20591 2975
rect 20533 2935 20591 2941
rect 11146 2904 11152 2916
rect 7138 2876 8239 2904
rect 8404 2876 11152 2904
rect 7138 2873 7150 2876
rect 7092 2867 7150 2873
rect 5537 2839 5595 2845
rect 5537 2805 5549 2839
rect 5583 2805 5595 2839
rect 5537 2799 5595 2805
rect 6178 2796 6184 2848
rect 6236 2836 6242 2848
rect 6236 2808 6281 2836
rect 6236 2796 6242 2808
rect 6822 2796 6828 2848
rect 6880 2836 6886 2848
rect 7742 2836 7748 2848
rect 6880 2808 7748 2836
rect 6880 2796 6886 2808
rect 7742 2796 7748 2808
rect 7800 2796 7806 2848
rect 8211 2836 8239 2876
rect 11146 2864 11152 2876
rect 11204 2864 11210 2916
rect 14001 2907 14059 2913
rect 14001 2904 14013 2907
rect 11808 2876 14013 2904
rect 8386 2836 8392 2848
rect 8211 2808 8392 2836
rect 8386 2796 8392 2808
rect 8444 2836 8450 2848
rect 8570 2836 8576 2848
rect 8444 2808 8576 2836
rect 8444 2796 8450 2808
rect 8570 2796 8576 2808
rect 8628 2836 8634 2848
rect 9861 2839 9919 2845
rect 9861 2836 9873 2839
rect 8628 2808 9873 2836
rect 8628 2796 8634 2808
rect 9861 2805 9873 2808
rect 9907 2805 9919 2839
rect 9861 2799 9919 2805
rect 10321 2839 10379 2845
rect 10321 2805 10333 2839
rect 10367 2836 10379 2839
rect 11808 2836 11836 2876
rect 14001 2873 14013 2876
rect 14047 2873 14059 2907
rect 14734 2904 14740 2916
rect 14695 2876 14740 2904
rect 14001 2867 14059 2873
rect 14734 2864 14740 2876
rect 14792 2864 14798 2916
rect 15010 2864 15016 2916
rect 15068 2904 15074 2916
rect 15473 2907 15531 2913
rect 15473 2904 15485 2907
rect 15068 2876 15485 2904
rect 15068 2864 15074 2876
rect 15473 2873 15485 2876
rect 15519 2873 15531 2907
rect 15473 2867 15531 2873
rect 16022 2864 16028 2916
rect 16080 2913 16086 2916
rect 16080 2907 16144 2913
rect 16080 2873 16098 2907
rect 16132 2873 16144 2907
rect 16080 2867 16144 2873
rect 16080 2864 16086 2867
rect 16206 2864 16212 2916
rect 16264 2904 16270 2916
rect 20548 2904 20576 2935
rect 16264 2876 20576 2904
rect 20809 2907 20867 2913
rect 16264 2864 16270 2876
rect 20809 2873 20821 2907
rect 20855 2904 20867 2907
rect 22186 2904 22192 2916
rect 20855 2876 22192 2904
rect 20855 2873 20867 2876
rect 20809 2867 20867 2873
rect 22186 2864 22192 2876
rect 22244 2864 22250 2916
rect 10367 2808 11836 2836
rect 14369 2839 14427 2845
rect 10367 2805 10379 2808
rect 10321 2799 10379 2805
rect 14369 2805 14381 2839
rect 14415 2836 14427 2839
rect 14458 2836 14464 2848
rect 14415 2808 14464 2836
rect 14415 2805 14427 2808
rect 14369 2799 14427 2805
rect 14458 2796 14464 2808
rect 14516 2796 14522 2848
rect 14829 2839 14887 2845
rect 14829 2805 14841 2839
rect 14875 2836 14887 2839
rect 16482 2836 16488 2848
rect 14875 2808 16488 2836
rect 14875 2805 14887 2808
rect 14829 2799 14887 2805
rect 16482 2796 16488 2808
rect 16540 2796 16546 2848
rect 17954 2796 17960 2848
rect 18012 2836 18018 2848
rect 18601 2839 18659 2845
rect 18601 2836 18613 2839
rect 18012 2808 18613 2836
rect 18012 2796 18018 2808
rect 18601 2805 18613 2808
rect 18647 2805 18659 2839
rect 18601 2799 18659 2805
rect 18693 2839 18751 2845
rect 18693 2805 18705 2839
rect 18739 2836 18751 2839
rect 19150 2836 19156 2848
rect 18739 2808 19156 2836
rect 18739 2805 18751 2808
rect 18693 2799 18751 2805
rect 19150 2796 19156 2808
rect 19208 2796 19214 2848
rect 20622 2796 20628 2848
rect 20680 2836 20686 2848
rect 22554 2836 22560 2848
rect 20680 2808 22560 2836
rect 20680 2796 20686 2808
rect 22554 2796 22560 2808
rect 22612 2796 22618 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 2038 2632 2044 2644
rect 1995 2604 2044 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 2038 2592 2044 2604
rect 2096 2592 2102 2644
rect 2317 2635 2375 2641
rect 2317 2601 2329 2635
rect 2363 2632 2375 2635
rect 2682 2632 2688 2644
rect 2363 2604 2688 2632
rect 2363 2601 2375 2604
rect 2317 2595 2375 2601
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 3326 2632 3332 2644
rect 3068 2604 3332 2632
rect 2590 2524 2596 2576
rect 2648 2564 2654 2576
rect 3068 2564 3096 2604
rect 3326 2592 3332 2604
rect 3384 2632 3390 2644
rect 5258 2632 5264 2644
rect 3384 2604 5264 2632
rect 3384 2592 3390 2604
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 5810 2592 5816 2644
rect 5868 2632 5874 2644
rect 5905 2635 5963 2641
rect 5905 2632 5917 2635
rect 5868 2604 5917 2632
rect 5868 2592 5874 2604
rect 5905 2601 5917 2604
rect 5951 2601 5963 2635
rect 5905 2595 5963 2601
rect 6178 2592 6184 2644
rect 6236 2632 6242 2644
rect 6917 2635 6975 2641
rect 6917 2632 6929 2635
rect 6236 2604 6929 2632
rect 6236 2592 6242 2604
rect 6917 2601 6929 2604
rect 6963 2601 6975 2635
rect 6917 2595 6975 2601
rect 7742 2592 7748 2644
rect 7800 2632 7806 2644
rect 8294 2632 8300 2644
rect 7800 2604 8300 2632
rect 7800 2592 7806 2604
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 8662 2592 8668 2644
rect 8720 2632 8726 2644
rect 10229 2635 10287 2641
rect 8720 2604 10180 2632
rect 8720 2592 8726 2604
rect 2648 2536 3096 2564
rect 2648 2524 2654 2536
rect 3142 2524 3148 2576
rect 3200 2564 3206 2576
rect 4678 2567 4736 2573
rect 4678 2564 4690 2567
rect 3200 2536 4690 2564
rect 3200 2524 3206 2536
rect 4678 2533 4690 2536
rect 4724 2533 4736 2567
rect 4678 2527 4736 2533
rect 5442 2524 5448 2576
rect 5500 2564 5506 2576
rect 6086 2564 6092 2576
rect 5500 2536 6092 2564
rect 5500 2524 5506 2536
rect 6086 2524 6092 2536
rect 6144 2564 6150 2576
rect 6365 2567 6423 2573
rect 6365 2564 6377 2567
rect 6144 2536 6377 2564
rect 6144 2524 6150 2536
rect 6365 2533 6377 2536
rect 6411 2533 6423 2567
rect 6365 2527 6423 2533
rect 6638 2524 6644 2576
rect 6696 2564 6702 2576
rect 7650 2564 7656 2576
rect 6696 2536 7656 2564
rect 6696 2524 6702 2536
rect 7650 2524 7656 2536
rect 7708 2524 7714 2576
rect 10152 2564 10180 2604
rect 10229 2601 10241 2635
rect 10275 2632 10287 2635
rect 10318 2632 10324 2644
rect 10275 2604 10324 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 10318 2592 10324 2604
rect 10376 2592 10382 2644
rect 10502 2592 10508 2644
rect 10560 2632 10566 2644
rect 11149 2635 11207 2641
rect 11149 2632 11161 2635
rect 10560 2604 11161 2632
rect 10560 2592 10566 2604
rect 11149 2601 11161 2604
rect 11195 2601 11207 2635
rect 11149 2595 11207 2601
rect 12621 2635 12679 2641
rect 12621 2601 12633 2635
rect 12667 2632 12679 2635
rect 12802 2632 12808 2644
rect 12667 2604 12808 2632
rect 12667 2601 12679 2604
rect 12621 2595 12679 2601
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 12986 2632 12992 2644
rect 12947 2604 12992 2632
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 14829 2635 14887 2641
rect 14829 2601 14841 2635
rect 14875 2632 14887 2635
rect 15930 2632 15936 2644
rect 14875 2604 15936 2632
rect 14875 2601 14887 2604
rect 14829 2595 14887 2601
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 16669 2635 16727 2641
rect 16669 2601 16681 2635
rect 16715 2632 16727 2635
rect 17126 2632 17132 2644
rect 16715 2604 17132 2632
rect 16715 2601 16727 2604
rect 16669 2595 16727 2601
rect 17126 2592 17132 2604
rect 17184 2592 17190 2644
rect 17221 2635 17279 2641
rect 17221 2601 17233 2635
rect 17267 2632 17279 2635
rect 17494 2632 17500 2644
rect 17267 2604 17500 2632
rect 17267 2601 17279 2604
rect 17221 2595 17279 2601
rect 17494 2592 17500 2604
rect 17552 2592 17558 2644
rect 18693 2635 18751 2641
rect 18693 2632 18705 2635
rect 18432 2604 18705 2632
rect 10689 2567 10747 2573
rect 10689 2564 10701 2567
rect 10152 2536 10701 2564
rect 10689 2533 10701 2536
rect 10735 2533 10747 2567
rect 13909 2567 13967 2573
rect 13909 2564 13921 2567
rect 10689 2527 10747 2533
rect 11900 2536 13921 2564
rect 1946 2456 1952 2508
rect 2004 2496 2010 2508
rect 2409 2499 2467 2505
rect 2409 2496 2421 2499
rect 2004 2468 2421 2496
rect 2004 2456 2010 2468
rect 2409 2465 2421 2468
rect 2455 2496 2467 2499
rect 3418 2496 3424 2508
rect 2455 2468 3424 2496
rect 2455 2465 2467 2468
rect 2409 2459 2467 2465
rect 3418 2456 3424 2468
rect 3476 2456 3482 2508
rect 3513 2499 3571 2505
rect 3513 2465 3525 2499
rect 3559 2496 3571 2499
rect 4430 2496 4436 2508
rect 3559 2468 4016 2496
rect 4391 2468 4436 2496
rect 3559 2465 3571 2468
rect 3513 2459 3571 2465
rect 2590 2428 2596 2440
rect 2551 2400 2596 2428
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 3605 2431 3663 2437
rect 3605 2428 3617 2431
rect 3099 2400 3617 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 3605 2397 3617 2400
rect 3651 2428 3663 2431
rect 3694 2428 3700 2440
rect 3651 2400 3700 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 3694 2388 3700 2400
rect 3752 2388 3758 2440
rect 3786 2388 3792 2440
rect 3844 2428 3850 2440
rect 3988 2428 4016 2468
rect 4430 2456 4436 2468
rect 4488 2456 4494 2508
rect 4982 2456 4988 2508
rect 5040 2496 5046 2508
rect 6273 2499 6331 2505
rect 6273 2496 6285 2499
rect 5040 2468 6285 2496
rect 5040 2456 5046 2468
rect 6273 2465 6285 2468
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 7190 2456 7196 2508
rect 7248 2496 7254 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 7248 2468 7297 2496
rect 7248 2456 7254 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 9122 2496 9128 2508
rect 7285 2459 7343 2465
rect 7576 2468 8616 2496
rect 9035 2468 9128 2496
rect 3844 2400 3889 2428
rect 3988 2400 4384 2428
rect 3844 2388 3850 2400
rect 4356 2372 4384 2400
rect 5534 2388 5540 2440
rect 5592 2428 5598 2440
rect 6457 2431 6515 2437
rect 6457 2428 6469 2431
rect 5592 2400 6469 2428
rect 5592 2388 5598 2400
rect 6457 2397 6469 2400
rect 6503 2397 6515 2431
rect 7374 2428 7380 2440
rect 7335 2400 7380 2428
rect 6457 2391 6515 2397
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 7576 2437 7604 2468
rect 8588 2440 8616 2468
rect 9122 2456 9128 2468
rect 9180 2496 9186 2508
rect 9950 2496 9956 2508
rect 9180 2468 9956 2496
rect 9180 2456 9186 2468
rect 9950 2456 9956 2468
rect 10008 2456 10014 2508
rect 10134 2496 10140 2508
rect 10095 2468 10140 2496
rect 10134 2456 10140 2468
rect 10192 2456 10198 2508
rect 10318 2456 10324 2508
rect 10376 2496 10382 2508
rect 10376 2468 11468 2496
rect 10376 2456 10382 2468
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2397 7619 2431
rect 7561 2391 7619 2397
rect 8294 2388 8300 2440
rect 8352 2428 8358 2440
rect 8389 2431 8447 2437
rect 8389 2428 8401 2431
rect 8352 2400 8401 2428
rect 8352 2388 8358 2400
rect 8389 2397 8401 2400
rect 8435 2397 8447 2431
rect 8570 2428 8576 2440
rect 8531 2400 8576 2428
rect 8389 2391 8447 2397
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 10410 2428 10416 2440
rect 10371 2400 10416 2428
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 11241 2431 11299 2437
rect 11241 2397 11253 2431
rect 11287 2397 11299 2431
rect 11241 2391 11299 2397
rect 11333 2431 11391 2437
rect 11333 2397 11345 2431
rect 11379 2397 11391 2431
rect 11440 2428 11468 2468
rect 11606 2456 11612 2508
rect 11664 2496 11670 2508
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 11664 2468 11805 2496
rect 11664 2456 11670 2468
rect 11793 2465 11805 2468
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 11900 2428 11928 2536
rect 13909 2533 13921 2536
rect 13955 2533 13967 2567
rect 13909 2527 13967 2533
rect 14737 2567 14795 2573
rect 14737 2533 14749 2567
rect 14783 2564 14795 2567
rect 16390 2564 16396 2576
rect 14783 2536 16396 2564
rect 14783 2533 14795 2536
rect 14737 2527 14795 2533
rect 16390 2524 16396 2536
rect 16448 2524 16454 2576
rect 16577 2567 16635 2573
rect 16577 2533 16589 2567
rect 16623 2564 16635 2567
rect 16850 2564 16856 2576
rect 16623 2536 16856 2564
rect 16623 2533 16635 2536
rect 16577 2527 16635 2533
rect 16850 2524 16856 2536
rect 16908 2524 16914 2576
rect 17586 2564 17592 2576
rect 17547 2536 17592 2564
rect 17586 2524 17592 2536
rect 17644 2524 17650 2576
rect 12250 2456 12256 2508
rect 12308 2496 12314 2508
rect 13633 2499 13691 2505
rect 13633 2496 13645 2499
rect 12308 2468 13645 2496
rect 12308 2456 12314 2468
rect 13633 2465 13645 2468
rect 13679 2465 13691 2499
rect 15194 2496 15200 2508
rect 13633 2459 13691 2465
rect 13740 2468 15200 2496
rect 11440 2400 11928 2428
rect 11333 2391 11391 2397
rect 3145 2363 3203 2369
rect 3145 2329 3157 2363
rect 3191 2360 3203 2363
rect 4154 2360 4160 2372
rect 3191 2332 4160 2360
rect 3191 2329 3203 2332
rect 3145 2323 3203 2329
rect 4154 2320 4160 2332
rect 4212 2320 4218 2372
rect 4338 2360 4344 2372
rect 4299 2332 4344 2360
rect 4338 2320 4344 2332
rect 4396 2320 4402 2372
rect 5813 2363 5871 2369
rect 5813 2329 5825 2363
rect 5859 2360 5871 2363
rect 5902 2360 5908 2372
rect 5859 2332 5908 2360
rect 5859 2329 5871 2332
rect 5813 2323 5871 2329
rect 5902 2320 5908 2332
rect 5960 2320 5966 2372
rect 7929 2363 7987 2369
rect 7929 2329 7941 2363
rect 7975 2360 7987 2363
rect 11256 2360 11284 2391
rect 7975 2332 11284 2360
rect 7975 2329 7987 2332
rect 7929 2323 7987 2329
rect 3786 2252 3792 2304
rect 3844 2292 3850 2304
rect 7834 2292 7840 2304
rect 3844 2264 7840 2292
rect 3844 2252 3850 2264
rect 7834 2252 7840 2264
rect 7892 2252 7898 2304
rect 9306 2292 9312 2304
rect 9267 2264 9312 2292
rect 9306 2252 9312 2264
rect 9364 2252 9370 2304
rect 9766 2292 9772 2304
rect 9727 2264 9772 2292
rect 9766 2252 9772 2264
rect 9824 2252 9830 2304
rect 10689 2295 10747 2301
rect 10689 2261 10701 2295
rect 10735 2292 10747 2295
rect 10781 2295 10839 2301
rect 10781 2292 10793 2295
rect 10735 2264 10793 2292
rect 10735 2261 10747 2264
rect 10689 2255 10747 2261
rect 10781 2261 10793 2264
rect 10827 2261 10839 2295
rect 10781 2255 10839 2261
rect 10870 2252 10876 2304
rect 10928 2292 10934 2304
rect 11348 2292 11376 2391
rect 11974 2388 11980 2440
rect 12032 2428 12038 2440
rect 12032 2400 12077 2428
rect 12032 2388 12038 2400
rect 12342 2388 12348 2440
rect 12400 2428 12406 2440
rect 13078 2428 13084 2440
rect 12400 2400 13084 2428
rect 12400 2388 12406 2400
rect 13078 2388 13084 2400
rect 13136 2388 13142 2440
rect 13170 2388 13176 2440
rect 13228 2428 13234 2440
rect 13228 2400 13273 2428
rect 13228 2388 13234 2400
rect 12434 2320 12440 2372
rect 12492 2360 12498 2372
rect 13740 2360 13768 2468
rect 15194 2456 15200 2468
rect 15252 2456 15258 2508
rect 15562 2456 15568 2508
rect 15620 2496 15626 2508
rect 15657 2499 15715 2505
rect 15657 2496 15669 2499
rect 15620 2468 15669 2496
rect 15620 2456 15626 2468
rect 15657 2465 15669 2468
rect 15703 2465 15715 2499
rect 17034 2496 17040 2508
rect 15657 2459 15715 2465
rect 16776 2468 17040 2496
rect 15013 2431 15071 2437
rect 15013 2397 15025 2431
rect 15059 2428 15071 2431
rect 16776 2428 16804 2468
rect 17034 2456 17040 2468
rect 17092 2456 17098 2508
rect 17678 2496 17684 2508
rect 17639 2468 17684 2496
rect 17678 2456 17684 2468
rect 17736 2456 17742 2508
rect 17954 2456 17960 2508
rect 18012 2496 18018 2508
rect 18432 2496 18460 2604
rect 18693 2601 18705 2604
rect 18739 2601 18751 2635
rect 18693 2595 18751 2601
rect 19337 2635 19395 2641
rect 19337 2601 19349 2635
rect 19383 2632 19395 2635
rect 19702 2632 19708 2644
rect 19383 2604 19564 2632
rect 19663 2604 19708 2632
rect 19383 2601 19395 2604
rect 19337 2595 19395 2601
rect 18782 2564 18788 2576
rect 18743 2536 18788 2564
rect 18782 2524 18788 2536
rect 18840 2524 18846 2576
rect 19536 2564 19564 2604
rect 19702 2592 19708 2604
rect 19760 2592 19766 2644
rect 20530 2632 20536 2644
rect 19812 2604 20536 2632
rect 19812 2564 19840 2604
rect 20530 2592 20536 2604
rect 20588 2592 20594 2644
rect 20622 2564 20628 2576
rect 19536 2536 19840 2564
rect 20583 2536 20628 2564
rect 20622 2524 20628 2536
rect 20680 2524 20686 2576
rect 18012 2468 18460 2496
rect 18012 2456 18018 2468
rect 19886 2456 19892 2508
rect 19944 2496 19950 2508
rect 20349 2499 20407 2505
rect 20349 2496 20361 2499
rect 19944 2468 20361 2496
rect 19944 2456 19950 2468
rect 20349 2465 20361 2468
rect 20395 2465 20407 2499
rect 20349 2459 20407 2465
rect 15059 2400 16804 2428
rect 16853 2431 16911 2437
rect 15059 2397 15071 2400
rect 15013 2391 15071 2397
rect 16853 2397 16865 2431
rect 16899 2428 16911 2431
rect 17773 2431 17831 2437
rect 17773 2428 17785 2431
rect 16899 2400 17785 2428
rect 16899 2397 16911 2400
rect 16853 2391 16911 2397
rect 17773 2397 17785 2400
rect 17819 2428 17831 2431
rect 18598 2428 18604 2440
rect 17819 2400 18604 2428
rect 17819 2397 17831 2400
rect 17773 2391 17831 2397
rect 18598 2388 18604 2400
rect 18656 2388 18662 2440
rect 18690 2388 18696 2440
rect 18748 2428 18754 2440
rect 18877 2431 18935 2437
rect 18877 2428 18889 2431
rect 18748 2400 18889 2428
rect 18748 2388 18754 2400
rect 18877 2397 18889 2400
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 19797 2431 19855 2437
rect 19797 2397 19809 2431
rect 19843 2397 19855 2431
rect 19978 2428 19984 2440
rect 19939 2400 19984 2428
rect 19797 2391 19855 2397
rect 12492 2332 13768 2360
rect 14369 2363 14427 2369
rect 12492 2320 12498 2332
rect 14369 2329 14381 2363
rect 14415 2360 14427 2363
rect 14458 2360 14464 2372
rect 14415 2332 14464 2360
rect 14415 2329 14427 2332
rect 14369 2323 14427 2329
rect 14458 2320 14464 2332
rect 14516 2320 14522 2372
rect 15841 2363 15899 2369
rect 15841 2329 15853 2363
rect 15887 2360 15899 2363
rect 17954 2360 17960 2372
rect 15887 2332 17960 2360
rect 15887 2329 15899 2332
rect 15841 2323 15899 2329
rect 17954 2320 17960 2332
rect 18012 2320 18018 2372
rect 18325 2363 18383 2369
rect 18325 2329 18337 2363
rect 18371 2360 18383 2363
rect 18966 2360 18972 2372
rect 18371 2332 18972 2360
rect 18371 2329 18383 2332
rect 18325 2323 18383 2329
rect 18966 2320 18972 2332
rect 19024 2320 19030 2372
rect 10928 2264 11376 2292
rect 16209 2295 16267 2301
rect 10928 2252 10934 2264
rect 16209 2261 16221 2295
rect 16255 2292 16267 2295
rect 16298 2292 16304 2304
rect 16255 2264 16304 2292
rect 16255 2261 16267 2264
rect 16209 2255 16267 2261
rect 16298 2252 16304 2264
rect 16356 2252 16362 2304
rect 17310 2252 17316 2304
rect 17368 2292 17374 2304
rect 19812 2292 19840 2391
rect 19978 2388 19984 2400
rect 20036 2388 20042 2440
rect 17368 2264 19840 2292
rect 17368 2252 17374 2264
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20438 2292 20444 2304
rect 20036 2264 20444 2292
rect 20036 2252 20042 2264
rect 20438 2252 20444 2264
rect 20496 2252 20502 2304
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 4154 2048 4160 2100
rect 4212 2088 4218 2100
rect 4982 2088 4988 2100
rect 4212 2060 4988 2088
rect 4212 2048 4218 2060
rect 4982 2048 4988 2060
rect 5040 2048 5046 2100
rect 9950 2048 9956 2100
rect 10008 2088 10014 2100
rect 16206 2088 16212 2100
rect 10008 2060 16212 2088
rect 10008 2048 10014 2060
rect 16206 2048 16212 2060
rect 16264 2048 16270 2100
rect 16574 2048 16580 2100
rect 16632 2088 16638 2100
rect 18598 2088 18604 2100
rect 16632 2060 18604 2088
rect 16632 2048 16638 2060
rect 18598 2048 18604 2060
rect 18656 2048 18662 2100
rect 18782 2048 18788 2100
rect 18840 2088 18846 2100
rect 19426 2088 19432 2100
rect 18840 2060 19432 2088
rect 18840 2048 18846 2060
rect 19426 2048 19432 2060
rect 19484 2048 19490 2100
rect 2774 1980 2780 2032
rect 2832 2020 2838 2032
rect 7006 2020 7012 2032
rect 2832 1992 7012 2020
rect 2832 1980 2838 1992
rect 7006 1980 7012 1992
rect 7064 1980 7070 2032
rect 8202 1980 8208 2032
rect 8260 2020 8266 2032
rect 10870 2020 10876 2032
rect 8260 1992 10876 2020
rect 8260 1980 8266 1992
rect 10870 1980 10876 1992
rect 10928 1980 10934 2032
rect 198 1912 204 1964
rect 256 1952 262 1964
rect 8294 1952 8300 1964
rect 256 1924 8300 1952
rect 256 1912 262 1924
rect 8294 1912 8300 1924
rect 8352 1952 8358 1964
rect 9030 1952 9036 1964
rect 8352 1924 9036 1952
rect 8352 1912 8358 1924
rect 9030 1912 9036 1924
rect 9088 1912 9094 1964
rect 9306 1912 9312 1964
rect 9364 1952 9370 1964
rect 21450 1952 21456 1964
rect 9364 1924 21456 1952
rect 9364 1912 9370 1924
rect 21450 1912 21456 1924
rect 21508 1912 21514 1964
rect 6546 1844 6552 1896
rect 6604 1884 6610 1896
rect 10318 1884 10324 1896
rect 6604 1856 10324 1884
rect 6604 1844 6610 1856
rect 10318 1844 10324 1856
rect 10376 1844 10382 1896
rect 11054 1844 11060 1896
rect 11112 1884 11118 1896
rect 19886 1884 19892 1896
rect 11112 1856 19892 1884
rect 11112 1844 11118 1856
rect 19886 1844 19892 1856
rect 19944 1844 19950 1896
rect 4890 1776 4896 1828
rect 4948 1816 4954 1828
rect 9766 1816 9772 1828
rect 4948 1788 9772 1816
rect 4948 1776 4954 1788
rect 9766 1776 9772 1788
rect 9824 1776 9830 1828
rect 10134 1776 10140 1828
rect 10192 1816 10198 1828
rect 10962 1816 10968 1828
rect 10192 1788 10968 1816
rect 10192 1776 10198 1788
rect 10962 1776 10968 1788
rect 11020 1776 11026 1828
rect 11149 1819 11207 1825
rect 11149 1785 11161 1819
rect 11195 1816 11207 1819
rect 11974 1816 11980 1828
rect 11195 1788 11980 1816
rect 11195 1785 11207 1788
rect 11149 1779 11207 1785
rect 11974 1776 11980 1788
rect 12032 1776 12038 1828
rect 18874 1776 18880 1828
rect 18932 1816 18938 1828
rect 20714 1816 20720 1828
rect 18932 1788 20720 1816
rect 18932 1776 18938 1788
rect 20714 1776 20720 1788
rect 20772 1776 20778 1828
rect 566 1708 572 1760
rect 624 1748 630 1760
rect 7742 1748 7748 1760
rect 624 1720 7748 1748
rect 624 1708 630 1720
rect 7742 1708 7748 1720
rect 7800 1708 7806 1760
rect 7834 1708 7840 1760
rect 7892 1748 7898 1760
rect 13538 1748 13544 1760
rect 7892 1720 13544 1748
rect 7892 1708 7898 1720
rect 13538 1708 13544 1720
rect 13596 1708 13602 1760
rect 5718 1640 5724 1692
rect 5776 1680 5782 1692
rect 11149 1683 11207 1689
rect 11149 1680 11161 1683
rect 5776 1652 11161 1680
rect 5776 1640 5782 1652
rect 11149 1649 11161 1652
rect 11195 1649 11207 1683
rect 17862 1680 17868 1692
rect 11149 1643 11207 1649
rect 11256 1652 17868 1680
rect 1302 1572 1308 1624
rect 1360 1612 1366 1624
rect 7558 1612 7564 1624
rect 1360 1584 7564 1612
rect 1360 1572 1366 1584
rect 7558 1572 7564 1584
rect 7616 1572 7622 1624
rect 8754 1612 8760 1624
rect 8667 1584 8760 1612
rect 8754 1572 8760 1584
rect 8812 1612 8818 1624
rect 11256 1612 11284 1652
rect 17862 1640 17868 1652
rect 17920 1640 17926 1692
rect 8812 1584 11284 1612
rect 8812 1572 8818 1584
rect 13814 1572 13820 1624
rect 13872 1612 13878 1624
rect 16206 1612 16212 1624
rect 13872 1584 16212 1612
rect 13872 1572 13878 1584
rect 16206 1572 16212 1584
rect 16264 1572 16270 1624
rect 17218 1572 17224 1624
rect 17276 1612 17282 1624
rect 19610 1612 19616 1624
rect 17276 1584 19616 1612
rect 17276 1572 17282 1584
rect 19610 1572 19616 1584
rect 19668 1572 19674 1624
rect 3970 1504 3976 1556
rect 4028 1544 4034 1556
rect 17586 1544 17592 1556
rect 4028 1516 17592 1544
rect 4028 1504 4034 1516
rect 17586 1504 17592 1516
rect 17644 1504 17650 1556
rect 7190 1436 7196 1488
rect 7248 1476 7254 1488
rect 11698 1476 11704 1488
rect 7248 1448 11704 1476
rect 7248 1436 7254 1448
rect 11698 1436 11704 1448
rect 11756 1436 11762 1488
rect 5350 1368 5356 1420
rect 5408 1408 5414 1420
rect 8757 1411 8815 1417
rect 8757 1408 8769 1411
rect 5408 1380 8769 1408
rect 5408 1368 5414 1380
rect 8757 1377 8769 1380
rect 8803 1377 8815 1411
rect 8757 1371 8815 1377
rect 9674 1368 9680 1420
rect 9732 1408 9738 1420
rect 14366 1408 14372 1420
rect 9732 1380 14372 1408
rect 9732 1368 9738 1380
rect 14366 1368 14372 1380
rect 14424 1368 14430 1420
rect 10778 1232 10784 1284
rect 10836 1272 10842 1284
rect 15102 1272 15108 1284
rect 10836 1244 15108 1272
rect 10836 1232 10842 1244
rect 15102 1232 15108 1244
rect 15160 1232 15166 1284
rect 2038 1164 2044 1216
rect 2096 1204 2102 1216
rect 7190 1204 7196 1216
rect 2096 1176 7196 1204
rect 2096 1164 2102 1176
rect 7190 1164 7196 1176
rect 7248 1164 7254 1216
rect 1670 1096 1676 1148
rect 1728 1136 1734 1148
rect 7374 1136 7380 1148
rect 1728 1108 7380 1136
rect 1728 1096 1734 1108
rect 7374 1096 7380 1108
rect 7432 1096 7438 1148
<< via1 >>
rect 4068 21360 4120 21412
rect 10508 21360 10560 21412
rect 3700 21088 3752 21140
rect 8760 21088 8812 21140
rect 14464 20680 14516 20732
rect 18144 20680 18196 20732
rect 1676 20476 1728 20528
rect 4252 20476 4304 20528
rect 2596 20408 2648 20460
rect 8576 20408 8628 20460
rect 4712 20340 4764 20392
rect 5172 20340 5224 20392
rect 9404 20340 9456 20392
rect 10784 20340 10836 20392
rect 14372 20340 14424 20392
rect 21456 20340 21508 20392
rect 3792 20272 3844 20324
rect 10876 20272 10928 20324
rect 19616 20272 19668 20324
rect 20352 20272 20404 20324
rect 4068 20204 4120 20256
rect 13176 20204 13228 20256
rect 13728 20204 13780 20256
rect 19064 20204 19116 20256
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 3792 20000 3844 20052
rect 6644 20000 6696 20052
rect 10232 20043 10284 20052
rect 10232 20009 10241 20043
rect 10241 20009 10275 20043
rect 10275 20009 10284 20043
rect 10232 20000 10284 20009
rect 2504 19932 2556 19984
rect 2596 19864 2648 19916
rect 3240 19907 3292 19916
rect 3240 19873 3249 19907
rect 3249 19873 3283 19907
rect 3283 19873 3292 19907
rect 3240 19864 3292 19873
rect 4988 19864 5040 19916
rect 5448 19907 5500 19916
rect 1860 19839 1912 19848
rect 1860 19805 1869 19839
rect 1869 19805 1903 19839
rect 1903 19805 1912 19839
rect 1860 19796 1912 19805
rect 2780 19796 2832 19848
rect 4252 19796 4304 19848
rect 4712 19839 4764 19848
rect 4712 19805 4721 19839
rect 4721 19805 4755 19839
rect 4755 19805 4764 19839
rect 4712 19796 4764 19805
rect 4160 19728 4212 19780
rect 5448 19873 5457 19907
rect 5457 19873 5491 19907
rect 5491 19873 5500 19907
rect 5448 19864 5500 19873
rect 6092 19907 6144 19916
rect 6092 19873 6101 19907
rect 6101 19873 6135 19907
rect 6135 19873 6144 19907
rect 6092 19864 6144 19873
rect 6920 19932 6972 19984
rect 7104 19932 7156 19984
rect 7472 19932 7524 19984
rect 9680 19932 9732 19984
rect 10968 19932 11020 19984
rect 14372 20000 14424 20052
rect 18052 20000 18104 20052
rect 22560 20000 22612 20052
rect 12992 19932 13044 19984
rect 16948 19932 17000 19984
rect 17960 19932 18012 19984
rect 19892 19975 19944 19984
rect 6736 19864 6788 19916
rect 5264 19796 5316 19848
rect 8392 19864 8444 19916
rect 10140 19907 10192 19916
rect 10140 19873 10149 19907
rect 10149 19873 10183 19907
rect 10183 19873 10192 19907
rect 10140 19864 10192 19873
rect 5356 19728 5408 19780
rect 6184 19660 6236 19712
rect 9036 19839 9088 19848
rect 9036 19805 9045 19839
rect 9045 19805 9079 19839
rect 9079 19805 9088 19839
rect 9036 19796 9088 19805
rect 8392 19728 8444 19780
rect 9220 19728 9272 19780
rect 10324 19864 10376 19916
rect 10876 19864 10928 19916
rect 12624 19907 12676 19916
rect 12624 19873 12633 19907
rect 12633 19873 12667 19907
rect 12667 19873 12676 19907
rect 12624 19864 12676 19873
rect 12072 19839 12124 19848
rect 12072 19805 12081 19839
rect 12081 19805 12115 19839
rect 12115 19805 12124 19839
rect 12072 19796 12124 19805
rect 13452 19796 13504 19848
rect 14188 19839 14240 19848
rect 14188 19805 14197 19839
rect 14197 19805 14231 19839
rect 14231 19805 14240 19839
rect 14188 19796 14240 19805
rect 15108 19796 15160 19848
rect 13728 19771 13780 19780
rect 13728 19737 13737 19771
rect 13737 19737 13771 19771
rect 13771 19737 13780 19771
rect 13728 19728 13780 19737
rect 9680 19660 9732 19712
rect 9772 19703 9824 19712
rect 9772 19669 9781 19703
rect 9781 19669 9815 19703
rect 9815 19669 9824 19703
rect 9772 19660 9824 19669
rect 10048 19660 10100 19712
rect 10600 19660 10652 19712
rect 12808 19660 12860 19712
rect 12900 19660 12952 19712
rect 15200 19660 15252 19712
rect 16580 19864 16632 19916
rect 16764 19907 16816 19916
rect 16764 19873 16773 19907
rect 16773 19873 16807 19907
rect 16807 19873 16816 19907
rect 16764 19864 16816 19873
rect 17500 19907 17552 19916
rect 17500 19873 17509 19907
rect 17509 19873 17543 19907
rect 17543 19873 17552 19907
rect 17500 19864 17552 19873
rect 18880 19907 18932 19916
rect 15936 19839 15988 19848
rect 15936 19805 15945 19839
rect 15945 19805 15979 19839
rect 15979 19805 15988 19839
rect 15936 19796 15988 19805
rect 16120 19839 16172 19848
rect 16120 19805 16129 19839
rect 16129 19805 16163 19839
rect 16163 19805 16172 19839
rect 16120 19796 16172 19805
rect 16212 19728 16264 19780
rect 18880 19873 18889 19907
rect 18889 19873 18923 19907
rect 18923 19873 18932 19907
rect 18880 19864 18932 19873
rect 19616 19907 19668 19916
rect 19616 19873 19625 19907
rect 19625 19873 19659 19907
rect 19659 19873 19668 19907
rect 19616 19864 19668 19873
rect 19892 19941 19901 19975
rect 19901 19941 19935 19975
rect 19935 19941 19944 19975
rect 19892 19932 19944 19941
rect 20628 19975 20680 19984
rect 20628 19941 20637 19975
rect 20637 19941 20671 19975
rect 20671 19941 20680 19975
rect 20628 19932 20680 19941
rect 20352 19907 20404 19916
rect 20352 19873 20361 19907
rect 20361 19873 20395 19907
rect 20395 19873 20404 19907
rect 20352 19864 20404 19873
rect 22192 19796 22244 19848
rect 17132 19660 17184 19712
rect 18604 19660 18656 19712
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 3332 19431 3384 19440
rect 3332 19397 3341 19431
rect 3341 19397 3375 19431
rect 3375 19397 3384 19431
rect 3332 19388 3384 19397
rect 3792 19431 3844 19440
rect 3792 19397 3801 19431
rect 3801 19397 3835 19431
rect 3835 19397 3844 19431
rect 3792 19388 3844 19397
rect 1952 19295 2004 19304
rect 940 19184 992 19236
rect 1584 19184 1636 19236
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 2412 19295 2464 19304
rect 2412 19261 2421 19295
rect 2421 19261 2455 19295
rect 2455 19261 2464 19295
rect 2412 19252 2464 19261
rect 2504 19184 2556 19236
rect 1308 19116 1360 19168
rect 2872 19252 2924 19304
rect 3056 19252 3108 19304
rect 4068 19320 4120 19372
rect 4344 19320 4396 19372
rect 5816 19456 5868 19508
rect 7196 19456 7248 19508
rect 8392 19499 8444 19508
rect 8392 19465 8401 19499
rect 8401 19465 8435 19499
rect 8435 19465 8444 19499
rect 8392 19456 8444 19465
rect 9496 19456 9548 19508
rect 11612 19456 11664 19508
rect 12440 19499 12492 19508
rect 12440 19465 12449 19499
rect 12449 19465 12483 19499
rect 12483 19465 12492 19499
rect 12440 19456 12492 19465
rect 14280 19456 14332 19508
rect 10324 19388 10376 19440
rect 4252 19252 4304 19304
rect 4804 19295 4856 19304
rect 4804 19261 4813 19295
rect 4813 19261 4847 19295
rect 4847 19261 4856 19295
rect 4804 19252 4856 19261
rect 5356 19252 5408 19304
rect 5632 19252 5684 19304
rect 6552 19252 6604 19304
rect 7104 19252 7156 19304
rect 2688 19116 2740 19168
rect 4160 19116 4212 19168
rect 5448 19184 5500 19236
rect 5540 19184 5592 19236
rect 8668 19252 8720 19304
rect 12072 19320 12124 19372
rect 13728 19320 13780 19372
rect 9680 19252 9732 19304
rect 12440 19252 12492 19304
rect 13452 19295 13504 19304
rect 13452 19261 13461 19295
rect 13461 19261 13495 19295
rect 13495 19261 13504 19295
rect 13452 19252 13504 19261
rect 14004 19252 14056 19304
rect 17960 19456 18012 19508
rect 18880 19456 18932 19508
rect 16948 19320 17000 19372
rect 17408 19320 17460 19372
rect 20444 19320 20496 19372
rect 7748 19184 7800 19236
rect 8300 19184 8352 19236
rect 9588 19184 9640 19236
rect 9956 19184 10008 19236
rect 4896 19116 4948 19168
rect 5816 19116 5868 19168
rect 6368 19116 6420 19168
rect 8392 19116 8444 19168
rect 10048 19116 10100 19168
rect 10324 19116 10376 19168
rect 10508 19116 10560 19168
rect 11888 19184 11940 19236
rect 11704 19159 11756 19168
rect 11704 19125 11713 19159
rect 11713 19125 11747 19159
rect 11747 19125 11756 19159
rect 11704 19116 11756 19125
rect 11796 19116 11848 19168
rect 13084 19184 13136 19236
rect 12164 19116 12216 19168
rect 13820 19116 13872 19168
rect 16856 19184 16908 19236
rect 17040 19252 17092 19304
rect 17500 19295 17552 19304
rect 17500 19261 17509 19295
rect 17509 19261 17543 19295
rect 17543 19261 17552 19295
rect 17500 19252 17552 19261
rect 18696 19252 18748 19304
rect 19800 19252 19852 19304
rect 17776 19184 17828 19236
rect 18144 19184 18196 19236
rect 19616 19184 19668 19236
rect 16396 19116 16448 19168
rect 17868 19116 17920 19168
rect 18880 19116 18932 19168
rect 20168 19159 20220 19168
rect 20168 19125 20177 19159
rect 20177 19125 20211 19159
rect 20211 19125 20220 19159
rect 20168 19116 20220 19125
rect 20536 19159 20588 19168
rect 20536 19125 20545 19159
rect 20545 19125 20579 19159
rect 20579 19125 20588 19159
rect 20536 19116 20588 19125
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 2320 18955 2372 18964
rect 2320 18921 2329 18955
rect 2329 18921 2363 18955
rect 2363 18921 2372 18955
rect 2320 18912 2372 18921
rect 3240 18912 3292 18964
rect 5080 18912 5132 18964
rect 6184 18955 6236 18964
rect 6184 18921 6193 18955
rect 6193 18921 6227 18955
rect 6227 18921 6236 18955
rect 6184 18912 6236 18921
rect 9496 18912 9548 18964
rect 572 18844 624 18896
rect 2688 18844 2740 18896
rect 2136 18776 2188 18828
rect 4804 18844 4856 18896
rect 4896 18844 4948 18896
rect 8392 18844 8444 18896
rect 9588 18844 9640 18896
rect 10048 18955 10100 18964
rect 10048 18921 10057 18955
rect 10057 18921 10091 18955
rect 10091 18921 10100 18955
rect 10048 18912 10100 18921
rect 12164 18912 12216 18964
rect 14372 18912 14424 18964
rect 17224 18912 17276 18964
rect 17316 18912 17368 18964
rect 4712 18776 4764 18828
rect 6368 18776 6420 18828
rect 6736 18819 6788 18828
rect 6736 18785 6745 18819
rect 6745 18785 6779 18819
rect 6779 18785 6788 18819
rect 6736 18776 6788 18785
rect 7104 18776 7156 18828
rect 2044 18708 2096 18760
rect 2412 18751 2464 18760
rect 2412 18717 2421 18751
rect 2421 18717 2455 18751
rect 2455 18717 2464 18751
rect 2412 18708 2464 18717
rect 2688 18708 2740 18760
rect 3424 18751 3476 18760
rect 3424 18717 3433 18751
rect 3433 18717 3467 18751
rect 3467 18717 3476 18751
rect 3424 18708 3476 18717
rect 1584 18615 1636 18624
rect 1584 18581 1593 18615
rect 1593 18581 1627 18615
rect 1627 18581 1636 18615
rect 1584 18572 1636 18581
rect 2872 18572 2924 18624
rect 5816 18708 5868 18760
rect 8668 18776 8720 18828
rect 10232 18844 10284 18896
rect 9128 18708 9180 18760
rect 9864 18776 9916 18828
rect 9956 18776 10008 18828
rect 12716 18844 12768 18896
rect 13084 18844 13136 18896
rect 13544 18844 13596 18896
rect 15476 18844 15528 18896
rect 17592 18844 17644 18896
rect 18788 18844 18840 18896
rect 19340 18844 19392 18896
rect 12072 18776 12124 18828
rect 10784 18708 10836 18760
rect 11152 18708 11204 18760
rect 13636 18776 13688 18828
rect 13820 18776 13872 18828
rect 15292 18819 15344 18828
rect 15292 18785 15301 18819
rect 15301 18785 15335 18819
rect 15335 18785 15344 18819
rect 15292 18776 15344 18785
rect 16120 18819 16172 18828
rect 16120 18785 16154 18819
rect 16154 18785 16172 18819
rect 16120 18776 16172 18785
rect 16948 18776 17000 18828
rect 17500 18819 17552 18828
rect 17500 18785 17509 18819
rect 17509 18785 17543 18819
rect 17543 18785 17552 18819
rect 17500 18776 17552 18785
rect 10508 18640 10560 18692
rect 15476 18708 15528 18760
rect 17040 18708 17092 18760
rect 18972 18776 19024 18828
rect 19156 18819 19208 18828
rect 19156 18785 19165 18819
rect 19165 18785 19199 18819
rect 19199 18785 19208 18819
rect 19156 18776 19208 18785
rect 18788 18708 18840 18760
rect 19800 18708 19852 18760
rect 20444 18751 20496 18760
rect 20444 18717 20453 18751
rect 20453 18717 20487 18751
rect 20487 18717 20496 18751
rect 20444 18708 20496 18717
rect 14280 18640 14332 18692
rect 5356 18572 5408 18624
rect 5724 18615 5776 18624
rect 5724 18581 5733 18615
rect 5733 18581 5767 18615
rect 5767 18581 5776 18615
rect 5724 18572 5776 18581
rect 5908 18572 5960 18624
rect 7380 18572 7432 18624
rect 8024 18572 8076 18624
rect 11612 18572 11664 18624
rect 11704 18572 11756 18624
rect 14096 18572 14148 18624
rect 14188 18572 14240 18624
rect 16856 18640 16908 18692
rect 20536 18640 20588 18692
rect 16764 18572 16816 18624
rect 17224 18615 17276 18624
rect 17224 18581 17233 18615
rect 17233 18581 17267 18615
rect 17267 18581 17276 18615
rect 17224 18572 17276 18581
rect 18972 18572 19024 18624
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 2412 18368 2464 18420
rect 4804 18368 4856 18420
rect 5724 18368 5776 18420
rect 7472 18411 7524 18420
rect 7472 18377 7481 18411
rect 7481 18377 7515 18411
rect 7515 18377 7524 18411
rect 7472 18368 7524 18377
rect 9036 18368 9088 18420
rect 10140 18368 10192 18420
rect 12072 18411 12124 18420
rect 12072 18377 12081 18411
rect 12081 18377 12115 18411
rect 12115 18377 12124 18411
rect 12072 18368 12124 18377
rect 12624 18368 12676 18420
rect 12716 18368 12768 18420
rect 13268 18368 13320 18420
rect 14096 18368 14148 18420
rect 1952 18164 2004 18216
rect 2044 18164 2096 18216
rect 3056 18164 3108 18216
rect 4804 18232 4856 18284
rect 7288 18300 7340 18352
rect 7748 18300 7800 18352
rect 3792 18164 3844 18216
rect 6276 18232 6328 18284
rect 7564 18232 7616 18284
rect 6920 18207 6972 18216
rect 2964 18096 3016 18148
rect 2780 18028 2832 18080
rect 4712 18096 4764 18148
rect 5347 18139 5399 18148
rect 5347 18105 5356 18139
rect 5356 18105 5390 18139
rect 5390 18105 5399 18139
rect 5347 18096 5399 18105
rect 6920 18173 6929 18207
rect 6929 18173 6963 18207
rect 6963 18173 6972 18207
rect 6920 18164 6972 18173
rect 8116 18275 8168 18284
rect 8116 18241 8125 18275
rect 8125 18241 8159 18275
rect 8159 18241 8168 18275
rect 8116 18232 8168 18241
rect 9588 18232 9640 18284
rect 4344 18028 4396 18080
rect 4896 18028 4948 18080
rect 5448 18028 5500 18080
rect 5816 18028 5868 18080
rect 6276 18028 6328 18080
rect 6828 18028 6880 18080
rect 7104 18096 7156 18148
rect 7748 18096 7800 18148
rect 8576 18096 8628 18148
rect 9404 18164 9456 18216
rect 11888 18300 11940 18352
rect 10416 18232 10468 18284
rect 10324 18164 10376 18216
rect 10508 18164 10560 18216
rect 12256 18232 12308 18284
rect 14556 18300 14608 18352
rect 17224 18368 17276 18420
rect 19156 18368 19208 18420
rect 12716 18164 12768 18216
rect 13084 18275 13136 18284
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 14188 18232 14240 18284
rect 14280 18232 14332 18284
rect 15200 18275 15252 18284
rect 15200 18241 15209 18275
rect 15209 18241 15243 18275
rect 15243 18241 15252 18275
rect 15200 18232 15252 18241
rect 17960 18300 18012 18352
rect 18604 18300 18656 18352
rect 21824 18300 21876 18352
rect 16120 18207 16172 18216
rect 10416 18096 10468 18148
rect 11888 18096 11940 18148
rect 11980 18096 12032 18148
rect 8300 18028 8352 18080
rect 8852 18071 8904 18080
rect 8852 18037 8861 18071
rect 8861 18037 8895 18071
rect 8895 18037 8904 18071
rect 8852 18028 8904 18037
rect 9036 18028 9088 18080
rect 9864 18071 9916 18080
rect 9864 18037 9873 18071
rect 9873 18037 9907 18071
rect 9907 18037 9916 18071
rect 9864 18028 9916 18037
rect 12808 18071 12860 18080
rect 12808 18037 12817 18071
rect 12817 18037 12851 18071
rect 12851 18037 12860 18071
rect 12808 18028 12860 18037
rect 13084 18028 13136 18080
rect 14464 18028 14516 18080
rect 15384 18096 15436 18148
rect 16120 18173 16129 18207
rect 16129 18173 16163 18207
rect 16163 18173 16172 18207
rect 16120 18164 16172 18173
rect 16764 18164 16816 18216
rect 17316 18232 17368 18284
rect 18512 18232 18564 18284
rect 17224 18207 17276 18216
rect 17224 18173 17233 18207
rect 17233 18173 17267 18207
rect 17267 18173 17276 18207
rect 17224 18164 17276 18173
rect 16304 18096 16356 18148
rect 17960 18096 18012 18148
rect 19248 18232 19300 18284
rect 20536 18232 20588 18284
rect 19156 18164 19208 18216
rect 19892 18096 19944 18148
rect 16396 18028 16448 18080
rect 17684 18028 17736 18080
rect 18236 18071 18288 18080
rect 18236 18037 18245 18071
rect 18245 18037 18279 18071
rect 18279 18037 18288 18071
rect 18236 18028 18288 18037
rect 18420 18071 18472 18080
rect 18420 18037 18429 18071
rect 18429 18037 18463 18071
rect 18463 18037 18472 18071
rect 18420 18028 18472 18037
rect 19156 18028 19208 18080
rect 20628 18071 20680 18080
rect 20628 18037 20637 18071
rect 20637 18037 20671 18071
rect 20671 18037 20680 18071
rect 20628 18028 20680 18037
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1676 17824 1728 17876
rect 2872 17867 2924 17876
rect 204 17756 256 17808
rect 1860 17799 1912 17808
rect 1860 17765 1869 17799
rect 1869 17765 1903 17799
rect 1903 17765 1912 17799
rect 1860 17756 1912 17765
rect 2872 17833 2881 17867
rect 2881 17833 2915 17867
rect 2915 17833 2924 17867
rect 2872 17824 2924 17833
rect 3424 17824 3476 17876
rect 4344 17824 4396 17876
rect 5080 17867 5132 17876
rect 5080 17833 5089 17867
rect 5089 17833 5123 17867
rect 5123 17833 5132 17867
rect 5080 17824 5132 17833
rect 6000 17824 6052 17876
rect 6092 17824 6144 17876
rect 8576 17867 8628 17876
rect 8576 17833 8585 17867
rect 8585 17833 8619 17867
rect 8619 17833 8628 17867
rect 8576 17824 8628 17833
rect 9220 17824 9272 17876
rect 2596 17688 2648 17740
rect 3056 17688 3108 17740
rect 3332 17688 3384 17740
rect 5264 17756 5316 17808
rect 7932 17756 7984 17808
rect 5448 17731 5500 17740
rect 5448 17697 5457 17731
rect 5457 17697 5491 17731
rect 5491 17697 5500 17731
rect 5448 17688 5500 17697
rect 5816 17688 5868 17740
rect 6736 17731 6788 17740
rect 6736 17697 6745 17731
rect 6745 17697 6779 17731
rect 6779 17697 6788 17731
rect 6736 17688 6788 17697
rect 7840 17688 7892 17740
rect 9220 17688 9272 17740
rect 9772 17756 9824 17808
rect 12348 17824 12400 17876
rect 13360 17824 13412 17876
rect 14556 17824 14608 17876
rect 11980 17756 12032 17808
rect 12256 17756 12308 17808
rect 13176 17756 13228 17808
rect 10048 17688 10100 17740
rect 10324 17731 10376 17740
rect 10324 17697 10333 17731
rect 10333 17697 10367 17731
rect 10367 17697 10376 17731
rect 10324 17688 10376 17697
rect 11152 17731 11204 17740
rect 2228 17620 2280 17672
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 3240 17620 3292 17672
rect 4712 17663 4764 17672
rect 4712 17629 4721 17663
rect 4721 17629 4755 17663
rect 4755 17629 4764 17663
rect 4712 17620 4764 17629
rect 5540 17663 5592 17672
rect 5540 17629 5549 17663
rect 5549 17629 5583 17663
rect 5583 17629 5592 17663
rect 5540 17620 5592 17629
rect 3608 17595 3660 17604
rect 3608 17561 3617 17595
rect 3617 17561 3651 17595
rect 3651 17561 3660 17595
rect 3608 17552 3660 17561
rect 6276 17620 6328 17672
rect 7472 17620 7524 17672
rect 8300 17620 8352 17672
rect 9128 17663 9180 17672
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 6000 17552 6052 17604
rect 11152 17697 11161 17731
rect 11161 17697 11195 17731
rect 11195 17697 11204 17731
rect 11152 17688 11204 17697
rect 13452 17731 13504 17740
rect 12164 17663 12216 17672
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 11796 17552 11848 17604
rect 12348 17620 12400 17672
rect 13452 17697 13461 17731
rect 13461 17697 13495 17731
rect 13495 17697 13504 17731
rect 15200 17756 15252 17808
rect 15660 17824 15712 17876
rect 17868 17824 17920 17876
rect 18052 17756 18104 17808
rect 19708 17756 19760 17808
rect 20352 17756 20404 17808
rect 13452 17688 13504 17697
rect 15568 17688 15620 17740
rect 14188 17620 14240 17672
rect 14372 17620 14424 17672
rect 14832 17663 14884 17672
rect 14832 17629 14841 17663
rect 14841 17629 14875 17663
rect 14875 17629 14884 17663
rect 14832 17620 14884 17629
rect 15292 17620 15344 17672
rect 16488 17688 16540 17740
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 16028 17620 16080 17672
rect 17040 17688 17092 17740
rect 20260 17688 20312 17740
rect 4988 17484 5040 17536
rect 9864 17484 9916 17536
rect 11152 17484 11204 17536
rect 15384 17552 15436 17604
rect 17500 17620 17552 17672
rect 17592 17620 17644 17672
rect 15936 17484 15988 17536
rect 17592 17484 17644 17536
rect 17868 17484 17920 17536
rect 19064 17663 19116 17672
rect 19064 17629 19073 17663
rect 19073 17629 19107 17663
rect 19107 17629 19116 17663
rect 19064 17620 19116 17629
rect 20536 17620 20588 17672
rect 19524 17527 19576 17536
rect 19524 17493 19533 17527
rect 19533 17493 19567 17527
rect 19567 17493 19576 17527
rect 19524 17484 19576 17493
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 3424 17280 3476 17332
rect 3608 17280 3660 17332
rect 5816 17280 5868 17332
rect 6552 17280 6604 17332
rect 7932 17280 7984 17332
rect 8852 17280 8904 17332
rect 9772 17280 9824 17332
rect 10876 17280 10928 17332
rect 12440 17323 12492 17332
rect 12440 17289 12449 17323
rect 12449 17289 12483 17323
rect 12483 17289 12492 17323
rect 12440 17280 12492 17289
rect 14832 17280 14884 17332
rect 15660 17280 15712 17332
rect 16304 17280 16356 17332
rect 16672 17280 16724 17332
rect 17316 17280 17368 17332
rect 17500 17280 17552 17332
rect 19984 17280 20036 17332
rect 20720 17280 20772 17332
rect 21272 17280 21324 17332
rect 3792 17144 3844 17196
rect 4252 17212 4304 17264
rect 5908 17212 5960 17264
rect 4712 17187 4764 17196
rect 4712 17153 4721 17187
rect 4721 17153 4755 17187
rect 4755 17153 4764 17187
rect 4712 17144 4764 17153
rect 5724 17144 5776 17196
rect 7840 17212 7892 17264
rect 8024 17255 8076 17264
rect 8024 17221 8033 17255
rect 8033 17221 8067 17255
rect 8067 17221 8076 17255
rect 8024 17212 8076 17221
rect 7196 17144 7248 17196
rect 8392 17144 8444 17196
rect 8852 17144 8904 17196
rect 9128 17144 9180 17196
rect 9588 17144 9640 17196
rect 12532 17212 12584 17264
rect 12624 17212 12676 17264
rect 1216 17076 1268 17128
rect 1768 17076 1820 17128
rect 2044 17076 2096 17128
rect 2688 17076 2740 17128
rect 3148 17076 3200 17128
rect 3976 17076 4028 17128
rect 4988 17076 5040 17128
rect 10784 17076 10836 17128
rect 11152 17144 11204 17196
rect 13084 17187 13136 17196
rect 13084 17153 13093 17187
rect 13093 17153 13127 17187
rect 13127 17153 13136 17187
rect 13084 17144 13136 17153
rect 15384 17187 15436 17196
rect 11888 17076 11940 17128
rect 13636 17076 13688 17128
rect 15384 17153 15393 17187
rect 15393 17153 15427 17187
rect 15427 17153 15436 17187
rect 15384 17144 15436 17153
rect 16672 17144 16724 17196
rect 18880 17144 18932 17196
rect 19708 17187 19760 17196
rect 19708 17153 19717 17187
rect 19717 17153 19751 17187
rect 19751 17153 19760 17187
rect 19708 17144 19760 17153
rect 20536 17144 20588 17196
rect 21548 17144 21600 17196
rect 17040 17076 17092 17128
rect 17592 17076 17644 17128
rect 2504 17008 2556 17060
rect 5080 16940 5132 16992
rect 6644 17008 6696 17060
rect 5632 16983 5684 16992
rect 5632 16949 5641 16983
rect 5641 16949 5675 16983
rect 5675 16949 5684 16983
rect 5632 16940 5684 16949
rect 5816 16940 5868 16992
rect 6828 16983 6880 16992
rect 6828 16949 6837 16983
rect 6837 16949 6871 16983
rect 6871 16949 6880 16983
rect 6828 16940 6880 16949
rect 8852 16983 8904 16992
rect 8852 16949 8861 16983
rect 8861 16949 8895 16983
rect 8895 16949 8904 16983
rect 8852 16940 8904 16949
rect 9680 17008 9732 17060
rect 11152 17008 11204 17060
rect 12532 17008 12584 17060
rect 13820 17008 13872 17060
rect 14004 17051 14056 17060
rect 14004 17017 14038 17051
rect 14038 17017 14056 17051
rect 14004 17008 14056 17017
rect 15200 17008 15252 17060
rect 9496 16940 9548 16992
rect 10416 16983 10468 16992
rect 10416 16949 10425 16983
rect 10425 16949 10459 16983
rect 10459 16949 10468 16983
rect 10416 16940 10468 16949
rect 11980 16940 12032 16992
rect 12808 16983 12860 16992
rect 12808 16949 12817 16983
rect 12817 16949 12851 16983
rect 12851 16949 12860 16983
rect 12808 16940 12860 16949
rect 13084 16940 13136 16992
rect 18328 17008 18380 17060
rect 19156 17008 19208 17060
rect 19248 17008 19300 17060
rect 21088 17008 21140 17060
rect 16948 16940 17000 16992
rect 17040 16940 17092 16992
rect 17960 16940 18012 16992
rect 18420 16983 18472 16992
rect 18420 16949 18429 16983
rect 18429 16949 18463 16983
rect 18463 16949 18472 16983
rect 18420 16940 18472 16949
rect 18880 16940 18932 16992
rect 20076 16983 20128 16992
rect 20076 16949 20085 16983
rect 20085 16949 20119 16983
rect 20119 16949 20128 16983
rect 20076 16940 20128 16949
rect 20536 16983 20588 16992
rect 20536 16949 20545 16983
rect 20545 16949 20579 16983
rect 20579 16949 20588 16983
rect 20536 16940 20588 16949
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 2504 16736 2556 16788
rect 4252 16736 4304 16788
rect 4528 16779 4580 16788
rect 4528 16745 4537 16779
rect 4537 16745 4571 16779
rect 4571 16745 4580 16779
rect 4528 16736 4580 16745
rect 5080 16736 5132 16788
rect 5356 16736 5408 16788
rect 6368 16736 6420 16788
rect 6644 16736 6696 16788
rect 6828 16736 6880 16788
rect 9588 16736 9640 16788
rect 11060 16736 11112 16788
rect 11888 16779 11940 16788
rect 11888 16745 11897 16779
rect 11897 16745 11931 16779
rect 11931 16745 11940 16779
rect 11888 16736 11940 16745
rect 2320 16711 2372 16720
rect 2320 16677 2329 16711
rect 2329 16677 2363 16711
rect 2363 16677 2372 16711
rect 2320 16668 2372 16677
rect 2412 16711 2464 16720
rect 2412 16677 2421 16711
rect 2421 16677 2455 16711
rect 2455 16677 2464 16711
rect 2412 16668 2464 16677
rect 3700 16668 3752 16720
rect 4988 16668 5040 16720
rect 3332 16643 3384 16652
rect 3332 16609 3341 16643
rect 3341 16609 3375 16643
rect 3375 16609 3384 16643
rect 3332 16600 3384 16609
rect 3424 16643 3476 16652
rect 3424 16609 3433 16643
rect 3433 16609 3467 16643
rect 3467 16609 3476 16643
rect 3424 16600 3476 16609
rect 4804 16600 4856 16652
rect 4896 16600 4948 16652
rect 5080 16600 5132 16652
rect 2688 16532 2740 16584
rect 5724 16668 5776 16720
rect 6920 16668 6972 16720
rect 7472 16668 7524 16720
rect 8300 16668 8352 16720
rect 8668 16668 8720 16720
rect 9496 16668 9548 16720
rect 13084 16736 13136 16788
rect 13728 16736 13780 16788
rect 15568 16779 15620 16788
rect 15568 16745 15577 16779
rect 15577 16745 15611 16779
rect 15611 16745 15620 16779
rect 15568 16736 15620 16745
rect 15936 16779 15988 16788
rect 15936 16745 15945 16779
rect 15945 16745 15979 16779
rect 15979 16745 15988 16779
rect 15936 16736 15988 16745
rect 16304 16736 16356 16788
rect 16580 16779 16632 16788
rect 16580 16745 16589 16779
rect 16589 16745 16623 16779
rect 16623 16745 16632 16779
rect 16580 16736 16632 16745
rect 17132 16736 17184 16788
rect 17592 16779 17644 16788
rect 5908 16600 5960 16652
rect 6000 16600 6052 16652
rect 6828 16600 6880 16652
rect 8576 16600 8628 16652
rect 9036 16600 9088 16652
rect 9312 16600 9364 16652
rect 9956 16643 10008 16652
rect 9956 16609 9965 16643
rect 9965 16609 9999 16643
rect 9999 16609 10008 16643
rect 9956 16600 10008 16609
rect 11796 16600 11848 16652
rect 11980 16600 12032 16652
rect 12716 16668 12768 16720
rect 12440 16600 12492 16652
rect 13084 16600 13136 16652
rect 14280 16668 14332 16720
rect 7472 16575 7524 16584
rect 4528 16464 4580 16516
rect 5080 16464 5132 16516
rect 3976 16396 4028 16448
rect 4896 16439 4948 16448
rect 4896 16405 4905 16439
rect 4905 16405 4939 16439
rect 4939 16405 4948 16439
rect 4896 16396 4948 16405
rect 5540 16396 5592 16448
rect 6920 16507 6972 16516
rect 6920 16473 6929 16507
rect 6929 16473 6963 16507
rect 6963 16473 6972 16507
rect 6920 16464 6972 16473
rect 7196 16396 7248 16448
rect 7472 16541 7481 16575
rect 7481 16541 7515 16575
rect 7515 16541 7524 16575
rect 7472 16532 7524 16541
rect 7748 16532 7800 16584
rect 10508 16575 10560 16584
rect 10508 16541 10517 16575
rect 10517 16541 10551 16575
rect 10551 16541 10560 16575
rect 10508 16532 10560 16541
rect 12072 16532 12124 16584
rect 10692 16396 10744 16448
rect 12532 16396 12584 16448
rect 14096 16532 14148 16584
rect 17316 16668 17368 16720
rect 17592 16745 17601 16779
rect 17601 16745 17635 16779
rect 17635 16745 17644 16779
rect 17592 16736 17644 16745
rect 19248 16736 19300 16788
rect 19616 16736 19668 16788
rect 20168 16736 20220 16788
rect 15200 16600 15252 16652
rect 15476 16600 15528 16652
rect 16028 16532 16080 16584
rect 14004 16464 14056 16516
rect 16396 16532 16448 16584
rect 16580 16464 16632 16516
rect 16856 16464 16908 16516
rect 13636 16396 13688 16448
rect 15844 16396 15896 16448
rect 17776 16532 17828 16584
rect 18328 16600 18380 16652
rect 17868 16464 17920 16516
rect 19248 16532 19300 16584
rect 18420 16464 18472 16516
rect 18604 16507 18656 16516
rect 18604 16473 18613 16507
rect 18613 16473 18647 16507
rect 18647 16473 18656 16507
rect 18604 16464 18656 16473
rect 18788 16464 18840 16516
rect 17592 16396 17644 16448
rect 19616 16439 19668 16448
rect 19616 16405 19625 16439
rect 19625 16405 19659 16439
rect 19659 16405 19668 16439
rect 19616 16396 19668 16405
rect 20168 16396 20220 16448
rect 20628 16396 20680 16448
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 1492 16192 1544 16244
rect 2596 16235 2648 16244
rect 2596 16201 2605 16235
rect 2605 16201 2639 16235
rect 2639 16201 2648 16235
rect 2596 16192 2648 16201
rect 5448 16192 5500 16244
rect 7748 16192 7800 16244
rect 8852 16192 8904 16244
rect 2688 16056 2740 16108
rect 3976 16056 4028 16108
rect 4252 16099 4304 16108
rect 4252 16065 4261 16099
rect 4261 16065 4295 16099
rect 4295 16065 4304 16099
rect 4252 16056 4304 16065
rect 4620 16124 4672 16176
rect 4804 16099 4856 16108
rect 4804 16065 4813 16099
rect 4813 16065 4847 16099
rect 4847 16065 4856 16099
rect 6184 16124 6236 16176
rect 4804 16056 4856 16065
rect 1676 15988 1728 16040
rect 2044 15988 2096 16040
rect 2136 16031 2188 16040
rect 2136 15997 2145 16031
rect 2145 15997 2179 16031
rect 2179 15997 2188 16031
rect 2136 15988 2188 15997
rect 2780 15988 2832 16040
rect 8760 16056 8812 16108
rect 9312 16056 9364 16108
rect 8944 15988 8996 16040
rect 9588 16056 9640 16108
rect 10508 15988 10560 16040
rect 12900 16192 12952 16244
rect 12992 16192 13044 16244
rect 14188 16192 14240 16244
rect 15108 16192 15160 16244
rect 15844 16235 15896 16244
rect 15844 16201 15853 16235
rect 15853 16201 15887 16235
rect 15887 16201 15896 16235
rect 15844 16192 15896 16201
rect 17960 16192 18012 16244
rect 18512 16192 18564 16244
rect 18788 16192 18840 16244
rect 13268 16056 13320 16108
rect 15108 16056 15160 16108
rect 15476 16099 15528 16108
rect 15476 16065 15485 16099
rect 15485 16065 15519 16099
rect 15519 16065 15528 16099
rect 15476 16056 15528 16065
rect 4620 15920 4672 15972
rect 5540 15920 5592 15972
rect 6920 15920 6972 15972
rect 7196 15920 7248 15972
rect 9128 15920 9180 15972
rect 10048 15920 10100 15972
rect 11612 15920 11664 15972
rect 13268 15920 13320 15972
rect 2412 15852 2464 15904
rect 4712 15852 4764 15904
rect 5632 15895 5684 15904
rect 5632 15861 5641 15895
rect 5641 15861 5675 15895
rect 5675 15861 5684 15895
rect 5632 15852 5684 15861
rect 6276 15895 6328 15904
rect 6276 15861 6285 15895
rect 6285 15861 6319 15895
rect 6319 15861 6328 15895
rect 6276 15852 6328 15861
rect 6368 15852 6420 15904
rect 7288 15852 7340 15904
rect 7472 15852 7524 15904
rect 8852 15895 8904 15904
rect 8852 15861 8861 15895
rect 8861 15861 8895 15895
rect 8895 15861 8904 15895
rect 8852 15852 8904 15861
rect 9680 15852 9732 15904
rect 10968 15852 11020 15904
rect 11796 15895 11848 15904
rect 11796 15861 11805 15895
rect 11805 15861 11839 15895
rect 11839 15861 11848 15895
rect 11796 15852 11848 15861
rect 12716 15852 12768 15904
rect 12900 15895 12952 15904
rect 12900 15861 12909 15895
rect 12909 15861 12943 15895
rect 12943 15861 12952 15895
rect 12900 15852 12952 15861
rect 13820 15895 13872 15904
rect 13820 15861 13829 15895
rect 13829 15861 13863 15895
rect 13863 15861 13872 15895
rect 13820 15852 13872 15861
rect 16396 16099 16448 16108
rect 16396 16065 16405 16099
rect 16405 16065 16439 16099
rect 16439 16065 16448 16099
rect 16396 16056 16448 16065
rect 16212 15988 16264 16040
rect 16764 16124 16816 16176
rect 17132 16124 17184 16176
rect 16948 16056 17000 16108
rect 17684 16056 17736 16108
rect 18972 16124 19024 16176
rect 20444 16124 20496 16176
rect 19708 16099 19760 16108
rect 19708 16065 19717 16099
rect 19717 16065 19751 16099
rect 19751 16065 19760 16099
rect 19708 16056 19760 16065
rect 20628 16099 20680 16108
rect 20628 16065 20637 16099
rect 20637 16065 20671 16099
rect 20671 16065 20680 16099
rect 20628 16056 20680 16065
rect 19248 15988 19300 16040
rect 16028 15852 16080 15904
rect 16120 15852 16172 15904
rect 16304 15852 16356 15904
rect 17132 15852 17184 15904
rect 17316 15895 17368 15904
rect 17316 15861 17325 15895
rect 17325 15861 17359 15895
rect 17359 15861 17368 15895
rect 17316 15852 17368 15861
rect 18604 15895 18656 15904
rect 18604 15861 18613 15895
rect 18613 15861 18647 15895
rect 18647 15861 18656 15895
rect 18604 15852 18656 15861
rect 19432 15895 19484 15904
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 19432 15852 19484 15861
rect 19524 15895 19576 15904
rect 19524 15861 19533 15895
rect 19533 15861 19567 15895
rect 19567 15861 19576 15895
rect 19524 15852 19576 15861
rect 19984 15852 20036 15904
rect 20536 15895 20588 15904
rect 20536 15861 20545 15895
rect 20545 15861 20579 15895
rect 20579 15861 20588 15895
rect 20536 15852 20588 15861
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 2320 15691 2372 15700
rect 2320 15657 2329 15691
rect 2329 15657 2363 15691
rect 2363 15657 2372 15691
rect 2320 15648 2372 15657
rect 4068 15648 4120 15700
rect 6092 15648 6144 15700
rect 6276 15648 6328 15700
rect 9680 15691 9732 15700
rect 9680 15657 9689 15691
rect 9689 15657 9723 15691
rect 9723 15657 9732 15691
rect 9680 15648 9732 15657
rect 13820 15648 13872 15700
rect 4620 15580 4672 15632
rect 2228 15512 2280 15564
rect 1492 15444 1544 15496
rect 2596 15512 2648 15564
rect 4804 15512 4856 15564
rect 5448 15512 5500 15564
rect 6460 15512 6512 15564
rect 2780 15444 2832 15496
rect 3792 15444 3844 15496
rect 6000 15487 6052 15496
rect 4896 15376 4948 15428
rect 6000 15453 6009 15487
rect 6009 15453 6043 15487
rect 6043 15453 6052 15487
rect 6000 15444 6052 15453
rect 6184 15487 6236 15496
rect 6184 15453 6193 15487
rect 6193 15453 6227 15487
rect 6227 15453 6236 15487
rect 6184 15444 6236 15453
rect 6276 15376 6328 15428
rect 7196 15555 7248 15564
rect 7196 15521 7230 15555
rect 7230 15521 7248 15555
rect 7196 15512 7248 15521
rect 7472 15512 7524 15564
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 2412 15308 2464 15360
rect 2964 15351 3016 15360
rect 2964 15317 2973 15351
rect 2973 15317 3007 15351
rect 3007 15317 3016 15351
rect 2964 15308 3016 15317
rect 5264 15308 5316 15360
rect 5540 15351 5592 15360
rect 5540 15317 5549 15351
rect 5549 15317 5583 15351
rect 5583 15317 5592 15351
rect 5540 15308 5592 15317
rect 6368 15308 6420 15360
rect 6644 15308 6696 15360
rect 8300 15419 8352 15428
rect 8300 15385 8309 15419
rect 8309 15385 8343 15419
rect 8343 15385 8352 15419
rect 8300 15376 8352 15385
rect 7840 15308 7892 15360
rect 8116 15308 8168 15360
rect 10508 15580 10560 15632
rect 9588 15512 9640 15564
rect 10692 15512 10744 15564
rect 12072 15580 12124 15632
rect 13544 15580 13596 15632
rect 16304 15648 16356 15700
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 9956 15444 10008 15496
rect 13636 15512 13688 15564
rect 14096 15512 14148 15564
rect 9496 15376 9548 15428
rect 14280 15444 14332 15496
rect 17316 15580 17368 15632
rect 18972 15580 19024 15632
rect 19616 15648 19668 15700
rect 20536 15580 20588 15632
rect 15200 15512 15252 15564
rect 15568 15444 15620 15496
rect 16764 15555 16816 15564
rect 16764 15521 16773 15555
rect 16773 15521 16807 15555
rect 16807 15521 16816 15555
rect 16764 15512 16816 15521
rect 16856 15487 16908 15496
rect 15476 15376 15528 15428
rect 16856 15453 16865 15487
rect 16865 15453 16899 15487
rect 16899 15453 16908 15487
rect 16856 15444 16908 15453
rect 8760 15308 8812 15360
rect 12256 15308 12308 15360
rect 14648 15308 14700 15360
rect 16672 15376 16724 15428
rect 16028 15308 16080 15360
rect 17500 15512 17552 15564
rect 18604 15555 18656 15564
rect 17316 15444 17368 15496
rect 17960 15487 18012 15496
rect 17960 15453 17969 15487
rect 17969 15453 18003 15487
rect 18003 15453 18012 15487
rect 18604 15521 18613 15555
rect 18613 15521 18647 15555
rect 18647 15521 18656 15555
rect 18604 15512 18656 15521
rect 18880 15487 18932 15496
rect 17960 15444 18012 15453
rect 18880 15453 18889 15487
rect 18889 15453 18923 15487
rect 18923 15453 18932 15487
rect 18880 15444 18932 15453
rect 20444 15512 20496 15564
rect 17408 15351 17460 15360
rect 17408 15317 17417 15351
rect 17417 15317 17451 15351
rect 17451 15317 17460 15351
rect 17408 15308 17460 15317
rect 17960 15308 18012 15360
rect 19616 15444 19668 15496
rect 21364 15308 21416 15360
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 2412 15104 2464 15156
rect 5264 15104 5316 15156
rect 5632 15104 5684 15156
rect 7196 15104 7248 15156
rect 6092 15036 6144 15088
rect 8116 15036 8168 15088
rect 6460 14968 6512 15020
rect 6644 14968 6696 15020
rect 11612 15104 11664 15156
rect 12808 15104 12860 15156
rect 15016 15104 15068 15156
rect 1768 14900 1820 14952
rect 2412 14900 2464 14952
rect 5080 14900 5132 14952
rect 6368 14900 6420 14952
rect 2780 14832 2832 14884
rect 3516 14832 3568 14884
rect 5264 14875 5316 14884
rect 4620 14764 4672 14816
rect 5264 14841 5298 14875
rect 5298 14841 5316 14875
rect 5264 14832 5316 14841
rect 6276 14832 6328 14884
rect 7748 14900 7800 14952
rect 7932 14900 7984 14952
rect 12164 14968 12216 15020
rect 12348 14968 12400 15020
rect 12716 14968 12768 15020
rect 17500 15036 17552 15088
rect 19432 15104 19484 15156
rect 14096 15011 14148 15020
rect 12440 14900 12492 14952
rect 13084 14900 13136 14952
rect 13728 14900 13780 14952
rect 14096 14977 14105 15011
rect 14105 14977 14139 15011
rect 14139 14977 14148 15011
rect 14096 14968 14148 14977
rect 15384 14968 15436 15020
rect 15476 14900 15528 14952
rect 18236 14968 18288 15020
rect 19708 15011 19760 15020
rect 19708 14977 19717 15011
rect 19717 14977 19751 15011
rect 19751 14977 19760 15011
rect 19708 14968 19760 14977
rect 20536 15011 20588 15020
rect 20536 14977 20545 15011
rect 20545 14977 20579 15011
rect 20579 14977 20588 15011
rect 20536 14968 20588 14977
rect 17040 14900 17092 14952
rect 6184 14764 6236 14816
rect 9680 14832 9732 14884
rect 11428 14832 11480 14884
rect 14648 14832 14700 14884
rect 9404 14764 9456 14816
rect 10876 14764 10928 14816
rect 12164 14764 12216 14816
rect 12808 14764 12860 14816
rect 15844 14832 15896 14884
rect 16672 14832 16724 14884
rect 16948 14832 17000 14884
rect 15476 14807 15528 14816
rect 15476 14773 15485 14807
rect 15485 14773 15519 14807
rect 15519 14773 15528 14807
rect 15752 14807 15804 14816
rect 15476 14764 15528 14773
rect 15752 14773 15761 14807
rect 15761 14773 15795 14807
rect 15795 14773 15804 14807
rect 15752 14764 15804 14773
rect 17316 14764 17368 14816
rect 18420 14832 18472 14884
rect 20076 14832 20128 14884
rect 18512 14764 18564 14816
rect 19064 14807 19116 14816
rect 19064 14773 19073 14807
rect 19073 14773 19107 14807
rect 19107 14773 19116 14807
rect 19064 14764 19116 14773
rect 19340 14764 19392 14816
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 5540 14560 5592 14612
rect 6920 14560 6972 14612
rect 8576 14603 8628 14612
rect 8576 14569 8585 14603
rect 8585 14569 8619 14603
rect 8619 14569 8628 14603
rect 8576 14560 8628 14569
rect 8852 14560 8904 14612
rect 9496 14560 9548 14612
rect 10232 14560 10284 14612
rect 3608 14492 3660 14544
rect 4528 14492 4580 14544
rect 2872 14424 2924 14476
rect 4712 14467 4764 14476
rect 4712 14433 4721 14467
rect 4721 14433 4755 14467
rect 4755 14433 4764 14467
rect 4712 14424 4764 14433
rect 5356 14424 5408 14476
rect 7288 14492 7340 14544
rect 7748 14492 7800 14544
rect 6920 14424 6972 14476
rect 7656 14424 7708 14476
rect 7932 14467 7984 14476
rect 7932 14433 7941 14467
rect 7941 14433 7975 14467
rect 7975 14433 7984 14467
rect 7932 14424 7984 14433
rect 8484 14492 8536 14544
rect 11888 14492 11940 14544
rect 16764 14560 16816 14612
rect 17776 14560 17828 14612
rect 20076 14603 20128 14612
rect 20076 14569 20085 14603
rect 20085 14569 20119 14603
rect 20119 14569 20128 14603
rect 20076 14560 20128 14569
rect 20812 14560 20864 14612
rect 12716 14535 12768 14544
rect 12716 14501 12725 14535
rect 12725 14501 12759 14535
rect 12759 14501 12768 14535
rect 12716 14492 12768 14501
rect 9772 14424 9824 14476
rect 11060 14424 11112 14476
rect 11612 14424 11664 14476
rect 2780 14356 2832 14408
rect 4620 14356 4672 14408
rect 3332 14288 3384 14340
rect 3608 14288 3660 14340
rect 4988 14356 5040 14408
rect 2780 14220 2832 14272
rect 5356 14220 5408 14272
rect 7380 14356 7432 14408
rect 8116 14399 8168 14408
rect 8116 14365 8125 14399
rect 8125 14365 8159 14399
rect 8159 14365 8168 14399
rect 8116 14356 8168 14365
rect 8576 14356 8628 14408
rect 8760 14356 8812 14408
rect 9128 14399 9180 14408
rect 9128 14365 9137 14399
rect 9137 14365 9171 14399
rect 9171 14365 9180 14399
rect 9128 14356 9180 14365
rect 9864 14356 9916 14408
rect 10876 14399 10928 14408
rect 10876 14365 10885 14399
rect 10885 14365 10919 14399
rect 10919 14365 10928 14399
rect 10876 14356 10928 14365
rect 11520 14356 11572 14408
rect 5540 14220 5592 14272
rect 7472 14220 7524 14272
rect 8300 14220 8352 14272
rect 13084 14356 13136 14408
rect 17960 14492 18012 14544
rect 18052 14492 18104 14544
rect 15844 14424 15896 14476
rect 16028 14424 16080 14476
rect 17040 14467 17092 14476
rect 17040 14433 17049 14467
rect 17049 14433 17083 14467
rect 17083 14433 17092 14467
rect 17040 14424 17092 14433
rect 17316 14467 17368 14476
rect 17316 14433 17350 14467
rect 17350 14433 17368 14467
rect 17316 14424 17368 14433
rect 17592 14424 17644 14476
rect 15200 14356 15252 14408
rect 13360 14331 13412 14340
rect 13360 14297 13369 14331
rect 13369 14297 13403 14331
rect 13403 14297 13412 14331
rect 13360 14288 13412 14297
rect 13544 14288 13596 14340
rect 14924 14288 14976 14340
rect 16488 14399 16540 14408
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16672 14399 16724 14408
rect 16488 14356 16540 14365
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 16672 14356 16724 14365
rect 18236 14424 18288 14476
rect 21364 14492 21416 14544
rect 16764 14288 16816 14340
rect 18144 14288 18196 14340
rect 19708 14356 19760 14408
rect 20812 14356 20864 14408
rect 19340 14288 19392 14340
rect 11152 14220 11204 14272
rect 11612 14220 11664 14272
rect 13452 14220 13504 14272
rect 15936 14220 15988 14272
rect 16028 14220 16080 14272
rect 17684 14220 17736 14272
rect 17776 14220 17828 14272
rect 19708 14263 19760 14272
rect 19708 14229 19717 14263
rect 19717 14229 19751 14263
rect 19751 14229 19760 14263
rect 19708 14220 19760 14229
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 5540 14016 5592 14068
rect 6000 14016 6052 14068
rect 6736 14016 6788 14068
rect 2872 13991 2924 14000
rect 2872 13957 2881 13991
rect 2881 13957 2915 13991
rect 2915 13957 2924 13991
rect 2872 13948 2924 13957
rect 4896 13948 4948 14000
rect 2596 13880 2648 13932
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 6092 13880 6144 13932
rect 2964 13812 3016 13864
rect 2780 13744 2832 13796
rect 3516 13744 3568 13796
rect 3700 13744 3752 13796
rect 1400 13719 1452 13728
rect 1400 13685 1409 13719
rect 1409 13685 1443 13719
rect 1443 13685 1452 13719
rect 1400 13676 1452 13685
rect 1860 13676 1912 13728
rect 2596 13676 2648 13728
rect 3976 13676 4028 13728
rect 4988 13812 5040 13864
rect 5264 13812 5316 13864
rect 5356 13812 5408 13864
rect 6736 13880 6788 13932
rect 9680 14016 9732 14068
rect 12716 14016 12768 14068
rect 12808 14016 12860 14068
rect 13176 14016 13228 14068
rect 13728 14016 13780 14068
rect 14372 14016 14424 14068
rect 16304 14016 16356 14068
rect 16856 14016 16908 14068
rect 17040 14016 17092 14068
rect 17500 14016 17552 14068
rect 20904 14059 20956 14068
rect 12532 13948 12584 14000
rect 7288 13812 7340 13864
rect 8852 13812 8904 13864
rect 6552 13744 6604 13796
rect 9496 13812 9548 13864
rect 9680 13880 9732 13932
rect 10232 13880 10284 13932
rect 10876 13880 10928 13932
rect 14280 13880 14332 13932
rect 12072 13812 12124 13864
rect 6000 13676 6052 13728
rect 6276 13676 6328 13728
rect 8852 13676 8904 13728
rect 12256 13744 12308 13796
rect 14188 13812 14240 13864
rect 14648 13812 14700 13864
rect 15016 13812 15068 13864
rect 16672 13880 16724 13932
rect 13544 13744 13596 13796
rect 15200 13744 15252 13796
rect 16856 13744 16908 13796
rect 10324 13719 10376 13728
rect 10324 13685 10333 13719
rect 10333 13685 10367 13719
rect 10367 13685 10376 13719
rect 10324 13676 10376 13685
rect 11428 13719 11480 13728
rect 11428 13685 11437 13719
rect 11437 13685 11471 13719
rect 11471 13685 11480 13719
rect 11428 13676 11480 13685
rect 11704 13676 11756 13728
rect 15476 13676 15528 13728
rect 17132 13719 17184 13728
rect 17132 13685 17141 13719
rect 17141 13685 17175 13719
rect 17175 13685 17184 13719
rect 17132 13676 17184 13685
rect 17960 13880 18012 13932
rect 20904 14025 20913 14059
rect 20913 14025 20947 14059
rect 20947 14025 20956 14059
rect 20904 14016 20956 14025
rect 19432 13948 19484 14000
rect 19340 13880 19392 13932
rect 20168 13855 20220 13864
rect 17868 13744 17920 13796
rect 17592 13676 17644 13728
rect 17960 13676 18012 13728
rect 19248 13676 19300 13728
rect 20168 13821 20177 13855
rect 20177 13821 20211 13855
rect 20211 13821 20220 13855
rect 20168 13812 20220 13821
rect 20720 13855 20772 13864
rect 20720 13821 20729 13855
rect 20729 13821 20763 13855
rect 20763 13821 20772 13855
rect 20720 13812 20772 13821
rect 20076 13719 20128 13728
rect 20076 13685 20085 13719
rect 20085 13685 20119 13719
rect 20119 13685 20128 13719
rect 20076 13676 20128 13685
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 2412 13472 2464 13524
rect 3516 13472 3568 13524
rect 5448 13472 5500 13524
rect 7380 13472 7432 13524
rect 5080 13404 5132 13456
rect 6276 13404 6328 13456
rect 7288 13404 7340 13456
rect 7840 13404 7892 13456
rect 9864 13404 9916 13456
rect 10876 13404 10928 13456
rect 11060 13472 11112 13524
rect 11520 13472 11572 13524
rect 12072 13472 12124 13524
rect 11704 13404 11756 13456
rect 1584 13379 1636 13388
rect 1584 13345 1593 13379
rect 1593 13345 1627 13379
rect 1627 13345 1636 13379
rect 1584 13336 1636 13345
rect 2412 13336 2464 13388
rect 2596 13379 2648 13388
rect 2596 13345 2630 13379
rect 2630 13345 2648 13379
rect 2596 13336 2648 13345
rect 5448 13336 5500 13388
rect 4068 13268 4120 13320
rect 5632 13311 5684 13320
rect 5632 13277 5641 13311
rect 5641 13277 5675 13311
rect 5675 13277 5684 13311
rect 5632 13268 5684 13277
rect 5724 13311 5776 13320
rect 5724 13277 5733 13311
rect 5733 13277 5767 13311
rect 5767 13277 5776 13311
rect 5724 13268 5776 13277
rect 1952 13132 2004 13184
rect 6092 13200 6144 13252
rect 7748 13336 7800 13388
rect 8760 13336 8812 13388
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 8300 13268 8352 13320
rect 8484 13311 8536 13320
rect 8484 13277 8493 13311
rect 8493 13277 8527 13311
rect 8527 13277 8536 13311
rect 8484 13268 8536 13277
rect 9312 13336 9364 13388
rect 11428 13336 11480 13388
rect 11796 13336 11848 13388
rect 9496 13268 9548 13320
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 10232 13268 10284 13277
rect 10600 13268 10652 13320
rect 11704 13311 11756 13320
rect 11704 13277 11713 13311
rect 11713 13277 11747 13311
rect 11747 13277 11756 13311
rect 11704 13268 11756 13277
rect 14096 13404 14148 13456
rect 14556 13404 14608 13456
rect 15476 13472 15528 13524
rect 17132 13472 17184 13524
rect 17408 13472 17460 13524
rect 17868 13472 17920 13524
rect 19708 13472 19760 13524
rect 16856 13404 16908 13456
rect 18696 13404 18748 13456
rect 19064 13404 19116 13456
rect 12992 13311 13044 13320
rect 12992 13277 13001 13311
rect 13001 13277 13035 13311
rect 13035 13277 13044 13311
rect 12992 13268 13044 13277
rect 13636 13336 13688 13388
rect 14280 13336 14332 13388
rect 14648 13336 14700 13388
rect 16580 13336 16632 13388
rect 17776 13336 17828 13388
rect 18052 13336 18104 13388
rect 20352 13336 20404 13388
rect 13544 13311 13596 13320
rect 13544 13277 13553 13311
rect 13553 13277 13587 13311
rect 13587 13277 13596 13311
rect 13544 13268 13596 13277
rect 15200 13268 15252 13320
rect 15936 13311 15988 13320
rect 15936 13277 15945 13311
rect 15945 13277 15979 13311
rect 15979 13277 15988 13311
rect 15936 13268 15988 13277
rect 16856 13311 16908 13320
rect 16856 13277 16865 13311
rect 16865 13277 16899 13311
rect 16899 13277 16908 13311
rect 16856 13268 16908 13277
rect 16948 13311 17000 13320
rect 16948 13277 16957 13311
rect 16957 13277 16991 13311
rect 16991 13277 17000 13311
rect 16948 13268 17000 13277
rect 17316 13268 17368 13320
rect 18236 13268 18288 13320
rect 19064 13311 19116 13320
rect 19064 13277 19073 13311
rect 19073 13277 19107 13311
rect 19107 13277 19116 13311
rect 19064 13268 19116 13277
rect 19340 13268 19392 13320
rect 19708 13268 19760 13320
rect 19892 13268 19944 13320
rect 10324 13200 10376 13252
rect 3700 13175 3752 13184
rect 3700 13141 3709 13175
rect 3709 13141 3743 13175
rect 3743 13141 3752 13175
rect 3700 13132 3752 13141
rect 4160 13175 4212 13184
rect 4160 13141 4169 13175
rect 4169 13141 4203 13175
rect 4203 13141 4212 13175
rect 4160 13132 4212 13141
rect 4988 13132 5040 13184
rect 7656 13132 7708 13184
rect 9404 13132 9456 13184
rect 11060 13132 11112 13184
rect 18788 13200 18840 13252
rect 15384 13132 15436 13184
rect 15568 13132 15620 13184
rect 19340 13132 19392 13184
rect 19892 13132 19944 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 4160 12928 4212 12980
rect 5448 12971 5500 12980
rect 5448 12937 5457 12971
rect 5457 12937 5491 12971
rect 5491 12937 5500 12971
rect 5448 12928 5500 12937
rect 6460 12971 6512 12980
rect 6460 12937 6469 12971
rect 6469 12937 6503 12971
rect 6503 12937 6512 12971
rect 6460 12928 6512 12937
rect 6828 12928 6880 12980
rect 7196 12971 7248 12980
rect 7196 12937 7205 12971
rect 7205 12937 7239 12971
rect 7239 12937 7248 12971
rect 7196 12928 7248 12937
rect 7472 12928 7524 12980
rect 4068 12860 4120 12912
rect 6092 12860 6144 12912
rect 2412 12724 2464 12776
rect 3700 12724 3752 12776
rect 3608 12656 3660 12708
rect 5724 12792 5776 12844
rect 8760 12928 8812 12980
rect 10508 12928 10560 12980
rect 8484 12860 8536 12912
rect 9036 12860 9088 12912
rect 6552 12724 6604 12776
rect 7196 12724 7248 12776
rect 10508 12835 10560 12844
rect 10508 12801 10517 12835
rect 10517 12801 10551 12835
rect 10551 12801 10560 12835
rect 10508 12792 10560 12801
rect 6368 12656 6420 12708
rect 6828 12699 6880 12708
rect 6828 12665 6837 12699
rect 6837 12665 6871 12699
rect 6871 12665 6880 12699
rect 6828 12656 6880 12665
rect 7472 12656 7524 12708
rect 7840 12656 7892 12708
rect 9404 12724 9456 12776
rect 10324 12767 10376 12776
rect 10324 12733 10333 12767
rect 10333 12733 10367 12767
rect 10367 12733 10376 12767
rect 10324 12724 10376 12733
rect 11612 12928 11664 12980
rect 12072 12928 12124 12980
rect 12256 12928 12308 12980
rect 14832 12928 14884 12980
rect 14924 12928 14976 12980
rect 11060 12792 11112 12844
rect 11980 12860 12032 12912
rect 11888 12835 11940 12844
rect 11888 12801 11897 12835
rect 11897 12801 11931 12835
rect 11931 12801 11940 12835
rect 11888 12792 11940 12801
rect 11152 12724 11204 12776
rect 1952 12631 2004 12640
rect 1952 12597 1961 12631
rect 1961 12597 1995 12631
rect 1995 12597 2004 12631
rect 1952 12588 2004 12597
rect 3424 12588 3476 12640
rect 3700 12588 3752 12640
rect 4252 12631 4304 12640
rect 4252 12597 4261 12631
rect 4261 12597 4295 12631
rect 4295 12597 4304 12631
rect 4252 12588 4304 12597
rect 5264 12588 5316 12640
rect 5908 12631 5960 12640
rect 5908 12597 5917 12631
rect 5917 12597 5951 12631
rect 5951 12597 5960 12631
rect 5908 12588 5960 12597
rect 6092 12588 6144 12640
rect 6644 12588 6696 12640
rect 7288 12588 7340 12640
rect 8300 12588 8352 12640
rect 8944 12631 8996 12640
rect 8944 12597 8953 12631
rect 8953 12597 8987 12631
rect 8987 12597 8996 12631
rect 8944 12588 8996 12597
rect 10876 12656 10928 12708
rect 12716 12860 12768 12912
rect 14188 12860 14240 12912
rect 15200 12860 15252 12912
rect 15476 12860 15528 12912
rect 13820 12792 13872 12844
rect 16028 12928 16080 12980
rect 16488 12928 16540 12980
rect 15936 12860 15988 12912
rect 17316 12860 17368 12912
rect 19892 12928 19944 12980
rect 19248 12860 19300 12912
rect 19340 12860 19392 12912
rect 16948 12835 17000 12844
rect 12164 12724 12216 12776
rect 12440 12724 12492 12776
rect 13452 12724 13504 12776
rect 14280 12724 14332 12776
rect 16304 12724 16356 12776
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 16764 12724 16816 12776
rect 13360 12656 13412 12708
rect 13544 12656 13596 12708
rect 13912 12656 13964 12708
rect 14004 12656 14056 12708
rect 14924 12656 14976 12708
rect 18604 12792 18656 12844
rect 18788 12792 18840 12844
rect 18880 12724 18932 12776
rect 19064 12724 19116 12776
rect 19340 12724 19392 12776
rect 20444 12835 20496 12844
rect 20444 12801 20453 12835
rect 20453 12801 20487 12835
rect 20487 12801 20496 12835
rect 20444 12792 20496 12801
rect 18420 12699 18472 12708
rect 13268 12588 13320 12640
rect 13636 12588 13688 12640
rect 14556 12588 14608 12640
rect 16580 12588 16632 12640
rect 18420 12665 18429 12699
rect 18429 12665 18463 12699
rect 18463 12665 18472 12699
rect 18420 12656 18472 12665
rect 17960 12588 18012 12640
rect 19340 12631 19392 12640
rect 19340 12597 19349 12631
rect 19349 12597 19383 12631
rect 19383 12597 19392 12631
rect 19340 12588 19392 12597
rect 20812 12588 20864 12640
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 1124 12384 1176 12436
rect 1952 12427 2004 12436
rect 1952 12393 1961 12427
rect 1961 12393 1995 12427
rect 1995 12393 2004 12427
rect 1952 12384 2004 12393
rect 1492 12248 1544 12300
rect 3516 12248 3568 12300
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 3608 12223 3660 12232
rect 3608 12189 3617 12223
rect 3617 12189 3651 12223
rect 3651 12189 3660 12223
rect 3608 12180 3660 12189
rect 3884 12384 3936 12436
rect 5724 12384 5776 12436
rect 7104 12384 7156 12436
rect 7380 12427 7432 12436
rect 7380 12393 7389 12427
rect 7389 12393 7423 12427
rect 7423 12393 7432 12427
rect 7380 12384 7432 12393
rect 7656 12384 7708 12436
rect 8944 12384 8996 12436
rect 10324 12384 10376 12436
rect 10600 12384 10652 12436
rect 10876 12384 10928 12436
rect 11980 12384 12032 12436
rect 12992 12384 13044 12436
rect 14096 12427 14148 12436
rect 14096 12393 14105 12427
rect 14105 12393 14139 12427
rect 14139 12393 14148 12427
rect 14096 12384 14148 12393
rect 15752 12384 15804 12436
rect 15936 12384 15988 12436
rect 17040 12384 17092 12436
rect 6552 12316 6604 12368
rect 8116 12316 8168 12368
rect 8300 12316 8352 12368
rect 4804 12248 4856 12300
rect 6092 12248 6144 12300
rect 7564 12248 7616 12300
rect 8668 12248 8720 12300
rect 9496 12316 9548 12368
rect 13544 12316 13596 12368
rect 14188 12316 14240 12368
rect 18880 12384 18932 12436
rect 18972 12384 19024 12436
rect 19340 12384 19392 12436
rect 4252 12180 4304 12232
rect 4344 12180 4396 12232
rect 6920 12223 6972 12232
rect 6920 12189 6929 12223
rect 6929 12189 6963 12223
rect 6963 12189 6972 12223
rect 7840 12223 7892 12232
rect 6920 12180 6972 12189
rect 7840 12189 7849 12223
rect 7849 12189 7883 12223
rect 7883 12189 7892 12223
rect 7840 12180 7892 12189
rect 11060 12248 11112 12300
rect 5908 12112 5960 12164
rect 7104 12112 7156 12164
rect 8852 12180 8904 12232
rect 9036 12223 9088 12232
rect 9036 12189 9045 12223
rect 9045 12189 9079 12223
rect 9079 12189 9088 12223
rect 9036 12180 9088 12189
rect 4712 12044 4764 12096
rect 9772 12112 9824 12164
rect 12716 12248 12768 12300
rect 13820 12248 13872 12300
rect 13912 12248 13964 12300
rect 13544 12223 13596 12232
rect 8208 12044 8260 12096
rect 8576 12044 8628 12096
rect 10968 12044 11020 12096
rect 13544 12189 13553 12223
rect 13553 12189 13587 12223
rect 13587 12189 13596 12223
rect 13544 12180 13596 12189
rect 14372 12180 14424 12232
rect 13084 12112 13136 12164
rect 13636 12112 13688 12164
rect 14188 12112 14240 12164
rect 14832 12180 14884 12232
rect 15384 12180 15436 12232
rect 17500 12248 17552 12300
rect 17960 12316 18012 12368
rect 17776 12248 17828 12300
rect 19248 12316 19300 12368
rect 20904 12316 20956 12368
rect 18972 12248 19024 12300
rect 14924 12112 14976 12164
rect 15108 12112 15160 12164
rect 12440 12044 12492 12096
rect 12624 12044 12676 12096
rect 12992 12044 13044 12096
rect 15568 12112 15620 12164
rect 20536 12248 20588 12300
rect 20444 12180 20496 12232
rect 15844 12112 15896 12164
rect 16212 12044 16264 12096
rect 19248 12044 19300 12096
rect 19708 12044 19760 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 3240 11840 3292 11892
rect 3608 11840 3660 11892
rect 4160 11840 4212 11892
rect 5632 11840 5684 11892
rect 6368 11840 6420 11892
rect 7380 11840 7432 11892
rect 7840 11883 7892 11892
rect 7840 11849 7849 11883
rect 7849 11849 7883 11883
rect 7883 11849 7892 11883
rect 7840 11840 7892 11849
rect 8392 11840 8444 11892
rect 8576 11840 8628 11892
rect 9036 11883 9088 11892
rect 9036 11849 9045 11883
rect 9045 11849 9079 11883
rect 9079 11849 9088 11883
rect 9036 11840 9088 11849
rect 9864 11883 9916 11892
rect 9864 11849 9873 11883
rect 9873 11849 9907 11883
rect 9907 11849 9916 11883
rect 9864 11840 9916 11849
rect 4804 11772 4856 11824
rect 5356 11704 5408 11756
rect 7932 11772 7984 11824
rect 1676 11611 1728 11620
rect 1676 11577 1685 11611
rect 1685 11577 1719 11611
rect 1719 11577 1728 11611
rect 1676 11568 1728 11577
rect 1860 11568 1912 11620
rect 2412 11568 2464 11620
rect 3332 11636 3384 11688
rect 4896 11679 4948 11688
rect 4896 11645 4905 11679
rect 4905 11645 4939 11679
rect 4939 11645 4948 11679
rect 4896 11636 4948 11645
rect 6920 11704 6972 11756
rect 8116 11704 8168 11756
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 9312 11772 9364 11824
rect 12256 11840 12308 11892
rect 12716 11840 12768 11892
rect 8392 11704 8444 11713
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 10968 11704 11020 11756
rect 11980 11772 12032 11824
rect 13912 11772 13964 11824
rect 14280 11772 14332 11824
rect 15844 11840 15896 11892
rect 15936 11840 15988 11892
rect 16212 11840 16264 11892
rect 17684 11840 17736 11892
rect 17776 11840 17828 11892
rect 17316 11772 17368 11824
rect 20444 11840 20496 11892
rect 21180 11840 21232 11892
rect 19708 11815 19760 11824
rect 19708 11781 19717 11815
rect 19717 11781 19751 11815
rect 19751 11781 19760 11815
rect 19708 11772 19760 11781
rect 7840 11636 7892 11688
rect 8208 11679 8260 11688
rect 8208 11645 8217 11679
rect 8217 11645 8251 11679
rect 8251 11645 8260 11679
rect 8208 11636 8260 11645
rect 10692 11636 10744 11688
rect 4252 11568 4304 11620
rect 5724 11568 5776 11620
rect 10784 11568 10836 11620
rect 11152 11636 11204 11688
rect 11704 11704 11756 11756
rect 11888 11704 11940 11756
rect 12440 11747 12492 11756
rect 12440 11713 12449 11747
rect 12449 11713 12483 11747
rect 12483 11713 12492 11747
rect 12440 11704 12492 11713
rect 12716 11679 12768 11688
rect 12716 11645 12750 11679
rect 12750 11645 12768 11679
rect 12716 11636 12768 11645
rect 12992 11636 13044 11688
rect 14188 11704 14240 11756
rect 15384 11704 15436 11756
rect 15844 11704 15896 11756
rect 1952 11500 2004 11552
rect 4068 11500 4120 11552
rect 5908 11500 5960 11552
rect 6184 11500 6236 11552
rect 6828 11500 6880 11552
rect 9128 11500 9180 11552
rect 10048 11500 10100 11552
rect 10876 11500 10928 11552
rect 13728 11568 13780 11620
rect 14188 11568 14240 11620
rect 15936 11636 15988 11688
rect 16028 11636 16080 11688
rect 16396 11679 16448 11688
rect 16396 11645 16405 11679
rect 16405 11645 16439 11679
rect 16439 11645 16448 11679
rect 16396 11636 16448 11645
rect 17224 11636 17276 11688
rect 17960 11636 18012 11688
rect 19248 11704 19300 11756
rect 18880 11636 18932 11688
rect 20812 11772 20864 11824
rect 20812 11636 20864 11688
rect 14648 11611 14700 11620
rect 14648 11577 14671 11611
rect 14671 11577 14700 11611
rect 14648 11568 14700 11577
rect 14832 11568 14884 11620
rect 18420 11568 18472 11620
rect 11796 11500 11848 11552
rect 15108 11500 15160 11552
rect 16764 11500 16816 11552
rect 17132 11500 17184 11552
rect 17316 11543 17368 11552
rect 17316 11509 17325 11543
rect 17325 11509 17359 11543
rect 17359 11509 17368 11543
rect 17316 11500 17368 11509
rect 17408 11500 17460 11552
rect 19432 11500 19484 11552
rect 20536 11500 20588 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 3332 11296 3384 11348
rect 3516 11339 3568 11348
rect 3516 11305 3525 11339
rect 3525 11305 3559 11339
rect 3559 11305 3568 11339
rect 3516 11296 3568 11305
rect 4068 11339 4120 11348
rect 4068 11305 4077 11339
rect 4077 11305 4111 11339
rect 4111 11305 4120 11339
rect 4068 11296 4120 11305
rect 4160 11296 4212 11348
rect 3884 11228 3936 11280
rect 4712 11228 4764 11280
rect 1860 11203 1912 11212
rect 1860 11169 1869 11203
rect 1869 11169 1903 11203
rect 1903 11169 1912 11203
rect 1860 11160 1912 11169
rect 2688 11160 2740 11212
rect 4160 11160 4212 11212
rect 5080 11203 5132 11212
rect 5080 11169 5089 11203
rect 5089 11169 5123 11203
rect 5123 11169 5132 11203
rect 5080 11160 5132 11169
rect 4252 11092 4304 11144
rect 3240 11024 3292 11076
rect 5080 11024 5132 11076
rect 5356 11024 5408 11076
rect 8300 11296 8352 11348
rect 8392 11228 8444 11280
rect 9496 11296 9548 11348
rect 9772 11296 9824 11348
rect 9312 11228 9364 11280
rect 12624 11296 12676 11348
rect 12808 11296 12860 11348
rect 13176 11296 13228 11348
rect 13544 11296 13596 11348
rect 15660 11339 15712 11348
rect 5724 11203 5776 11212
rect 5724 11169 5733 11203
rect 5733 11169 5767 11203
rect 5767 11169 5776 11203
rect 5724 11160 5776 11169
rect 5540 11092 5592 11144
rect 6368 11160 6420 11212
rect 7288 11160 7340 11212
rect 8484 11160 8536 11212
rect 11796 11160 11848 11212
rect 12072 11160 12124 11212
rect 8392 11092 8444 11144
rect 11152 11092 11204 11144
rect 7104 11067 7156 11076
rect 7104 11033 7113 11067
rect 7113 11033 7147 11067
rect 7147 11033 7156 11067
rect 7104 11024 7156 11033
rect 7380 11024 7432 11076
rect 14096 11228 14148 11280
rect 14740 11228 14792 11280
rect 15660 11305 15669 11339
rect 15669 11305 15703 11339
rect 15703 11305 15712 11339
rect 15660 11296 15712 11305
rect 18512 11296 18564 11348
rect 18972 11296 19024 11348
rect 20536 11339 20588 11348
rect 20536 11305 20545 11339
rect 20545 11305 20579 11339
rect 20579 11305 20588 11339
rect 20536 11296 20588 11305
rect 15844 11228 15896 11280
rect 12440 11203 12492 11212
rect 12440 11169 12449 11203
rect 12449 11169 12483 11203
rect 12483 11169 12492 11203
rect 12440 11160 12492 11169
rect 13636 11160 13688 11212
rect 14372 11160 14424 11212
rect 13912 11092 13964 11144
rect 14004 11092 14056 11144
rect 7748 10956 7800 11008
rect 13636 11024 13688 11076
rect 14096 11067 14148 11076
rect 14096 11033 14105 11067
rect 14105 11033 14139 11067
rect 14139 11033 14148 11067
rect 14096 11024 14148 11033
rect 15476 11092 15528 11144
rect 17132 11228 17184 11280
rect 18144 11228 18196 11280
rect 19708 11228 19760 11280
rect 17408 11160 17460 11212
rect 17592 11160 17644 11212
rect 18972 11160 19024 11212
rect 20628 11160 20680 11212
rect 15844 11135 15896 11144
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 17040 11135 17092 11144
rect 17040 11101 17049 11135
rect 17049 11101 17083 11135
rect 17083 11101 17092 11135
rect 17040 11092 17092 11101
rect 17224 11135 17276 11144
rect 17224 11101 17233 11135
rect 17233 11101 17267 11135
rect 17267 11101 17276 11135
rect 17224 11092 17276 11101
rect 17868 11092 17920 11144
rect 20536 11092 20588 11144
rect 21548 11092 21600 11144
rect 18420 11024 18472 11076
rect 8852 10956 8904 11008
rect 12808 10956 12860 11008
rect 14556 10956 14608 11008
rect 15200 10956 15252 11008
rect 15936 10956 15988 11008
rect 17132 10956 17184 11008
rect 20444 10956 20496 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 3240 10795 3292 10804
rect 3240 10761 3249 10795
rect 3249 10761 3283 10795
rect 3283 10761 3292 10795
rect 3240 10752 3292 10761
rect 3700 10795 3752 10804
rect 3700 10761 3709 10795
rect 3709 10761 3743 10795
rect 3743 10761 3752 10795
rect 3700 10752 3752 10761
rect 4160 10752 4212 10804
rect 4712 10752 4764 10804
rect 7472 10752 7524 10804
rect 4068 10684 4120 10736
rect 4528 10659 4580 10668
rect 3516 10591 3568 10600
rect 3516 10557 3525 10591
rect 3525 10557 3559 10591
rect 3559 10557 3568 10591
rect 3516 10548 3568 10557
rect 2596 10480 2648 10532
rect 4528 10625 4537 10659
rect 4537 10625 4571 10659
rect 4571 10625 4580 10659
rect 4528 10616 4580 10625
rect 5448 10616 5500 10668
rect 7288 10616 7340 10668
rect 4896 10548 4948 10600
rect 5632 10548 5684 10600
rect 6184 10591 6236 10600
rect 6184 10557 6193 10591
rect 6193 10557 6227 10591
rect 6227 10557 6236 10591
rect 6184 10548 6236 10557
rect 6920 10548 6972 10600
rect 8668 10752 8720 10804
rect 9312 10752 9364 10804
rect 9036 10616 9088 10668
rect 8852 10548 8904 10600
rect 10416 10752 10468 10804
rect 10692 10752 10744 10804
rect 11060 10752 11112 10804
rect 13452 10752 13504 10804
rect 9772 10591 9824 10600
rect 9772 10557 9781 10591
rect 9781 10557 9815 10591
rect 9815 10557 9824 10591
rect 9772 10548 9824 10557
rect 12440 10684 12492 10736
rect 14188 10752 14240 10804
rect 17316 10752 17368 10804
rect 19064 10752 19116 10804
rect 13636 10616 13688 10668
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 15200 10616 15252 10668
rect 19432 10684 19484 10736
rect 2228 10412 2280 10464
rect 4712 10412 4764 10464
rect 6092 10480 6144 10532
rect 5908 10412 5960 10464
rect 10140 10480 10192 10532
rect 8300 10455 8352 10464
rect 8300 10421 8309 10455
rect 8309 10421 8343 10455
rect 8343 10421 8352 10455
rect 8300 10412 8352 10421
rect 10692 10412 10744 10464
rect 11336 10480 11388 10532
rect 13452 10548 13504 10600
rect 13820 10548 13872 10600
rect 12072 10480 12124 10532
rect 15384 10548 15436 10600
rect 17132 10616 17184 10668
rect 17500 10659 17552 10668
rect 17500 10625 17509 10659
rect 17509 10625 17543 10659
rect 17543 10625 17552 10659
rect 17500 10616 17552 10625
rect 15844 10548 15896 10600
rect 12164 10412 12216 10464
rect 14832 10480 14884 10532
rect 16304 10523 16356 10532
rect 12808 10455 12860 10464
rect 12808 10421 12817 10455
rect 12817 10421 12851 10455
rect 12851 10421 12860 10455
rect 12808 10412 12860 10421
rect 13820 10455 13872 10464
rect 13820 10421 13829 10455
rect 13829 10421 13863 10455
rect 13863 10421 13872 10455
rect 13820 10412 13872 10421
rect 14372 10412 14424 10464
rect 15108 10412 15160 10464
rect 15660 10412 15712 10464
rect 16304 10489 16313 10523
rect 16313 10489 16347 10523
rect 16347 10489 16356 10523
rect 16304 10480 16356 10489
rect 17132 10480 17184 10532
rect 17316 10523 17368 10532
rect 17316 10489 17325 10523
rect 17325 10489 17359 10523
rect 17359 10489 17368 10523
rect 17316 10480 17368 10489
rect 16212 10455 16264 10464
rect 16212 10421 16221 10455
rect 16221 10421 16255 10455
rect 16255 10421 16264 10455
rect 16212 10412 16264 10421
rect 16580 10412 16632 10464
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 18144 10548 18196 10600
rect 19248 10548 19300 10600
rect 19892 10616 19944 10668
rect 20444 10548 20496 10600
rect 17868 10480 17920 10532
rect 18880 10412 18932 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 1768 10208 1820 10260
rect 1860 10208 1912 10260
rect 2044 10208 2096 10260
rect 2872 10208 2924 10260
rect 4528 10208 4580 10260
rect 5632 10208 5684 10260
rect 6184 10208 6236 10260
rect 2780 10140 2832 10192
rect 6644 10208 6696 10260
rect 7196 10208 7248 10260
rect 8208 10251 8260 10260
rect 8208 10217 8217 10251
rect 8217 10217 8251 10251
rect 8251 10217 8260 10251
rect 8208 10208 8260 10217
rect 8300 10208 8352 10260
rect 9036 10208 9088 10260
rect 10508 10208 10560 10260
rect 10692 10251 10744 10260
rect 10692 10217 10701 10251
rect 10701 10217 10735 10251
rect 10735 10217 10744 10251
rect 10692 10208 10744 10217
rect 11060 10208 11112 10260
rect 12624 10208 12676 10260
rect 14464 10208 14516 10260
rect 16120 10208 16172 10260
rect 16212 10208 16264 10260
rect 17040 10208 17092 10260
rect 17500 10208 17552 10260
rect 18236 10208 18288 10260
rect 20168 10208 20220 10260
rect 20628 10208 20680 10260
rect 2320 10072 2372 10124
rect 2504 10115 2556 10124
rect 2504 10081 2513 10115
rect 2513 10081 2547 10115
rect 2547 10081 2556 10115
rect 2504 10072 2556 10081
rect 12532 10140 12584 10192
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 4160 10072 4212 10124
rect 4712 10072 4764 10124
rect 4896 10072 4948 10124
rect 7012 10072 7064 10124
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 6092 10004 6144 10056
rect 6644 10004 6696 10056
rect 7748 10072 7800 10124
rect 8024 10115 8076 10124
rect 8024 10081 8033 10115
rect 8033 10081 8067 10115
rect 8067 10081 8076 10115
rect 8024 10072 8076 10081
rect 8300 10072 8352 10124
rect 8668 10072 8720 10124
rect 9864 10072 9916 10124
rect 3884 9936 3936 9988
rect 2320 9868 2372 9920
rect 3516 9868 3568 9920
rect 6000 9911 6052 9920
rect 6000 9877 6009 9911
rect 6009 9877 6043 9911
rect 6043 9877 6052 9911
rect 6000 9868 6052 9877
rect 6828 9911 6880 9920
rect 6828 9877 6837 9911
rect 6837 9877 6871 9911
rect 6871 9877 6880 9911
rect 6828 9868 6880 9877
rect 7288 9936 7340 9988
rect 8760 10004 8812 10056
rect 8852 10004 8904 10056
rect 9036 10047 9088 10056
rect 9036 10013 9045 10047
rect 9045 10013 9079 10047
rect 9079 10013 9088 10047
rect 9036 10004 9088 10013
rect 9128 10047 9180 10056
rect 9128 10013 9137 10047
rect 9137 10013 9171 10047
rect 9171 10013 9180 10047
rect 9128 10004 9180 10013
rect 7472 9936 7524 9988
rect 7840 9936 7892 9988
rect 8116 9936 8168 9988
rect 8392 9936 8444 9988
rect 9956 10004 10008 10056
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 10508 10072 10560 10124
rect 11060 10115 11112 10124
rect 10600 10004 10652 10056
rect 11060 10081 11069 10115
rect 11069 10081 11103 10115
rect 11103 10081 11112 10115
rect 11060 10072 11112 10081
rect 11796 10072 11848 10124
rect 13452 10072 13504 10124
rect 14556 10072 14608 10124
rect 17132 10072 17184 10124
rect 18236 10072 18288 10124
rect 18420 10072 18472 10124
rect 19064 10115 19116 10124
rect 19064 10081 19073 10115
rect 19073 10081 19107 10115
rect 19107 10081 19116 10115
rect 19064 10072 19116 10081
rect 19616 10140 19668 10192
rect 19892 10072 19944 10124
rect 10508 9979 10560 9988
rect 10508 9945 10517 9979
rect 10517 9945 10551 9979
rect 10551 9945 10560 9979
rect 10508 9936 10560 9945
rect 11060 9936 11112 9988
rect 9680 9911 9732 9920
rect 9680 9877 9689 9911
rect 9689 9877 9723 9911
rect 9723 9877 9732 9911
rect 9680 9868 9732 9877
rect 9864 9868 9916 9920
rect 11704 10004 11756 10056
rect 12992 10047 13044 10056
rect 12992 10013 13001 10047
rect 13001 10013 13035 10047
rect 13035 10013 13044 10047
rect 12992 10004 13044 10013
rect 11612 9936 11664 9988
rect 12164 9936 12216 9988
rect 12072 9911 12124 9920
rect 12072 9877 12081 9911
rect 12081 9877 12115 9911
rect 12115 9877 12124 9911
rect 12072 9868 12124 9877
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 13452 9911 13504 9920
rect 12440 9868 12492 9877
rect 13452 9877 13461 9911
rect 13461 9877 13495 9911
rect 13495 9877 13504 9911
rect 13452 9868 13504 9877
rect 13544 9868 13596 9920
rect 14188 10004 14240 10056
rect 14924 10004 14976 10056
rect 17224 10047 17276 10056
rect 17224 10013 17233 10047
rect 17233 10013 17267 10047
rect 17267 10013 17276 10047
rect 17224 10004 17276 10013
rect 17500 10004 17552 10056
rect 17592 10004 17644 10056
rect 18328 10004 18380 10056
rect 14464 9868 14516 9920
rect 17040 9868 17092 9920
rect 18788 9936 18840 9988
rect 19064 9868 19116 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 2504 9664 2556 9716
rect 3884 9664 3936 9716
rect 4252 9596 4304 9648
rect 2596 9528 2648 9580
rect 1768 9460 1820 9512
rect 2412 9392 2464 9444
rect 3148 9528 3200 9580
rect 3332 9528 3384 9580
rect 3608 9528 3660 9580
rect 4160 9528 4212 9580
rect 3516 9503 3568 9512
rect 3516 9469 3525 9503
rect 3525 9469 3559 9503
rect 3559 9469 3568 9503
rect 3516 9460 3568 9469
rect 5448 9571 5500 9580
rect 5448 9537 5457 9571
rect 5457 9537 5491 9571
rect 5491 9537 5500 9571
rect 5448 9528 5500 9537
rect 8668 9664 8720 9716
rect 9128 9664 9180 9716
rect 10140 9707 10192 9716
rect 10140 9673 10149 9707
rect 10149 9673 10183 9707
rect 10183 9673 10192 9707
rect 10140 9664 10192 9673
rect 11888 9664 11940 9716
rect 13084 9664 13136 9716
rect 15108 9664 15160 9716
rect 16580 9664 16632 9716
rect 16764 9664 16816 9716
rect 11980 9639 12032 9648
rect 6460 9460 6512 9512
rect 6644 9460 6696 9512
rect 9772 9528 9824 9580
rect 11980 9605 11989 9639
rect 11989 9605 12023 9639
rect 12023 9605 12032 9639
rect 11980 9596 12032 9605
rect 15660 9596 15712 9648
rect 16856 9596 16908 9648
rect 17500 9596 17552 9648
rect 18144 9596 18196 9648
rect 19156 9596 19208 9648
rect 19892 9596 19944 9648
rect 11152 9528 11204 9580
rect 12256 9528 12308 9580
rect 14188 9528 14240 9580
rect 15292 9528 15344 9580
rect 5080 9392 5132 9444
rect 6368 9392 6420 9444
rect 9312 9460 9364 9512
rect 9864 9460 9916 9512
rect 10600 9460 10652 9512
rect 12348 9460 12400 9512
rect 13636 9460 13688 9512
rect 14280 9503 14332 9512
rect 14280 9469 14289 9503
rect 14289 9469 14323 9503
rect 14323 9469 14332 9503
rect 14280 9460 14332 9469
rect 15752 9528 15804 9580
rect 15844 9571 15896 9580
rect 15844 9537 15853 9571
rect 15853 9537 15887 9571
rect 15887 9537 15896 9571
rect 15844 9528 15896 9537
rect 17040 9528 17092 9580
rect 7196 9392 7248 9444
rect 7288 9392 7340 9444
rect 2504 9367 2556 9376
rect 2504 9333 2513 9367
rect 2513 9333 2547 9367
rect 2547 9333 2556 9367
rect 2504 9324 2556 9333
rect 3424 9324 3476 9376
rect 3608 9367 3660 9376
rect 3608 9333 3617 9367
rect 3617 9333 3651 9367
rect 3651 9333 3660 9367
rect 4528 9367 4580 9376
rect 3608 9324 3660 9333
rect 4528 9333 4537 9367
rect 4537 9333 4571 9367
rect 4571 9333 4580 9367
rect 4528 9324 4580 9333
rect 4620 9324 4672 9376
rect 4896 9367 4948 9376
rect 4896 9333 4905 9367
rect 4905 9333 4939 9367
rect 4939 9333 4948 9367
rect 4896 9324 4948 9333
rect 5264 9367 5316 9376
rect 5264 9333 5273 9367
rect 5273 9333 5307 9367
rect 5307 9333 5316 9367
rect 5264 9324 5316 9333
rect 5356 9367 5408 9376
rect 5356 9333 5365 9367
rect 5365 9333 5399 9367
rect 5399 9333 5408 9367
rect 5356 9324 5408 9333
rect 6276 9324 6328 9376
rect 8392 9324 8444 9376
rect 8852 9392 8904 9444
rect 9220 9392 9272 9444
rect 9772 9392 9824 9444
rect 11060 9392 11112 9444
rect 11980 9392 12032 9444
rect 12164 9392 12216 9444
rect 17592 9460 17644 9512
rect 18144 9460 18196 9512
rect 18788 9528 18840 9580
rect 19432 9528 19484 9580
rect 20444 9528 20496 9580
rect 20168 9460 20220 9512
rect 20536 9460 20588 9512
rect 16304 9392 16356 9444
rect 10416 9367 10468 9376
rect 10416 9333 10425 9367
rect 10425 9333 10459 9367
rect 10459 9333 10468 9367
rect 10416 9324 10468 9333
rect 10600 9324 10652 9376
rect 13084 9324 13136 9376
rect 14556 9324 14608 9376
rect 17868 9324 17920 9376
rect 19432 9367 19484 9376
rect 19432 9333 19441 9367
rect 19441 9333 19475 9367
rect 19475 9333 19484 9367
rect 19432 9324 19484 9333
rect 20444 9367 20496 9376
rect 20444 9333 20453 9367
rect 20453 9333 20487 9367
rect 20487 9333 20496 9367
rect 20444 9324 20496 9333
rect 20536 9367 20588 9376
rect 20536 9333 20545 9367
rect 20545 9333 20579 9367
rect 20579 9333 20588 9367
rect 20536 9324 20588 9333
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 2412 9163 2464 9172
rect 2412 9129 2421 9163
rect 2421 9129 2455 9163
rect 2455 9129 2464 9163
rect 2412 9120 2464 9129
rect 2780 9120 2832 9172
rect 3424 9120 3476 9172
rect 4528 9120 4580 9172
rect 5172 9120 5224 9172
rect 2320 9095 2372 9104
rect 2320 9061 2329 9095
rect 2329 9061 2363 9095
rect 2363 9061 2372 9095
rect 2320 9052 2372 9061
rect 3792 9052 3844 9104
rect 3884 9052 3936 9104
rect 6184 9120 6236 9172
rect 6460 9163 6512 9172
rect 6460 9129 6469 9163
rect 6469 9129 6503 9163
rect 6503 9129 6512 9163
rect 6460 9120 6512 9129
rect 7472 9120 7524 9172
rect 7748 9120 7800 9172
rect 9220 9163 9272 9172
rect 5448 9052 5500 9104
rect 1676 8984 1728 9036
rect 2688 8916 2740 8968
rect 3424 8959 3476 8968
rect 3424 8925 3433 8959
rect 3433 8925 3467 8959
rect 3467 8925 3476 8959
rect 3424 8916 3476 8925
rect 3056 8848 3108 8900
rect 3240 8848 3292 8900
rect 4160 8916 4212 8968
rect 4620 8959 4672 8968
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 4896 8984 4948 9036
rect 6184 8984 6236 9036
rect 6368 9052 6420 9104
rect 7748 8984 7800 9036
rect 8852 9052 8904 9104
rect 9220 9129 9229 9163
rect 9229 9129 9263 9163
rect 9263 9129 9272 9163
rect 9220 9120 9272 9129
rect 10416 9120 10468 9172
rect 10692 9120 10744 9172
rect 11796 9120 11848 9172
rect 12440 9120 12492 9172
rect 9312 9052 9364 9104
rect 9956 9052 10008 9104
rect 8392 8984 8444 9036
rect 9864 8984 9916 9036
rect 10600 8984 10652 9036
rect 12348 9052 12400 9104
rect 14096 9120 14148 9172
rect 15200 9120 15252 9172
rect 15844 9120 15896 9172
rect 16488 9120 16540 9172
rect 18144 9120 18196 9172
rect 19616 9163 19668 9172
rect 15292 9052 15344 9104
rect 15568 9052 15620 9104
rect 18604 9052 18656 9104
rect 19616 9129 19625 9163
rect 19625 9129 19659 9163
rect 19659 9129 19668 9163
rect 19616 9120 19668 9129
rect 20904 9052 20956 9104
rect 12992 8984 13044 9036
rect 14464 8984 14516 9036
rect 15016 8984 15068 9036
rect 16580 8984 16632 9036
rect 16948 8984 17000 9036
rect 17500 9027 17552 9036
rect 17500 8993 17509 9027
rect 17509 8993 17543 9027
rect 17543 8993 17552 9027
rect 17500 8984 17552 8993
rect 8852 8916 8904 8968
rect 10140 8916 10192 8968
rect 14004 8916 14056 8968
rect 14280 8916 14332 8968
rect 17132 8916 17184 8968
rect 6368 8848 6420 8900
rect 4988 8780 5040 8832
rect 5356 8780 5408 8832
rect 6644 8780 6696 8832
rect 8944 8848 8996 8900
rect 9220 8848 9272 8900
rect 8576 8780 8628 8832
rect 8852 8780 8904 8832
rect 9864 8780 9916 8832
rect 13912 8848 13964 8900
rect 12164 8780 12216 8832
rect 12624 8780 12676 8832
rect 13452 8780 13504 8832
rect 13636 8780 13688 8832
rect 16304 8848 16356 8900
rect 14924 8780 14976 8832
rect 15844 8780 15896 8832
rect 16028 8780 16080 8832
rect 17960 8984 18012 9036
rect 18328 8984 18380 9036
rect 19984 8984 20036 9036
rect 19340 8916 19392 8968
rect 18144 8848 18196 8900
rect 19156 8780 19208 8832
rect 19892 8780 19944 8832
rect 20720 8780 20772 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2504 8576 2556 8628
rect 3976 8576 4028 8628
rect 5172 8576 5224 8628
rect 6184 8576 6236 8628
rect 6552 8576 6604 8628
rect 6644 8576 6696 8628
rect 3424 8508 3476 8560
rect 3792 8508 3844 8560
rect 5448 8551 5500 8560
rect 5448 8517 5457 8551
rect 5457 8517 5491 8551
rect 5491 8517 5500 8551
rect 5448 8508 5500 8517
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 3240 8440 3292 8492
rect 7748 8576 7800 8628
rect 8208 8576 8260 8628
rect 12532 8576 12584 8628
rect 7840 8508 7892 8560
rect 9864 8508 9916 8560
rect 1400 8372 1452 8424
rect 3056 8372 3108 8424
rect 3332 8372 3384 8424
rect 3700 8372 3752 8424
rect 4068 8415 4120 8424
rect 4068 8381 4077 8415
rect 4077 8381 4111 8415
rect 4111 8381 4120 8415
rect 4068 8372 4120 8381
rect 4896 8372 4948 8424
rect 5080 8372 5132 8424
rect 8208 8440 8260 8492
rect 8392 8440 8444 8492
rect 8576 8440 8628 8492
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 10140 8483 10192 8492
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 11060 8483 11112 8492
rect 11060 8449 11069 8483
rect 11069 8449 11103 8483
rect 11103 8449 11112 8483
rect 11060 8440 11112 8449
rect 11980 8551 12032 8560
rect 11980 8517 11989 8551
rect 11989 8517 12023 8551
rect 12023 8517 12032 8551
rect 11980 8508 12032 8517
rect 13636 8576 13688 8628
rect 13912 8576 13964 8628
rect 18512 8576 18564 8628
rect 19064 8619 19116 8628
rect 19064 8585 19073 8619
rect 19073 8585 19107 8619
rect 19107 8585 19116 8619
rect 19064 8576 19116 8585
rect 19708 8576 19760 8628
rect 20444 8576 20496 8628
rect 12808 8508 12860 8560
rect 14464 8551 14516 8560
rect 14464 8517 14473 8551
rect 14473 8517 14507 8551
rect 14507 8517 14516 8551
rect 14464 8508 14516 8517
rect 17132 8508 17184 8560
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 13544 8440 13596 8492
rect 14096 8483 14148 8492
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 14280 8440 14332 8492
rect 14372 8440 14424 8492
rect 15016 8483 15068 8492
rect 15016 8449 15025 8483
rect 15025 8449 15059 8483
rect 15059 8449 15068 8483
rect 15016 8440 15068 8449
rect 15752 8440 15804 8492
rect 19432 8508 19484 8560
rect 6460 8372 6512 8424
rect 8852 8415 8904 8424
rect 4160 8304 4212 8356
rect 4344 8347 4396 8356
rect 4344 8313 4378 8347
rect 4378 8313 4396 8347
rect 4344 8304 4396 8313
rect 7104 8347 7156 8356
rect 7104 8313 7138 8347
rect 7138 8313 7156 8347
rect 8852 8381 8861 8415
rect 8861 8381 8895 8415
rect 8895 8381 8904 8415
rect 8852 8372 8904 8381
rect 9128 8372 9180 8424
rect 11796 8415 11848 8424
rect 11796 8381 11805 8415
rect 11805 8381 11839 8415
rect 11839 8381 11848 8415
rect 11796 8372 11848 8381
rect 13728 8372 13780 8424
rect 13912 8415 13964 8424
rect 13912 8381 13921 8415
rect 13921 8381 13955 8415
rect 13955 8381 13964 8415
rect 13912 8372 13964 8381
rect 15108 8372 15160 8424
rect 15568 8415 15620 8424
rect 15568 8381 15577 8415
rect 15577 8381 15611 8415
rect 15611 8381 15620 8415
rect 15568 8372 15620 8381
rect 16028 8372 16080 8424
rect 18420 8440 18472 8492
rect 18788 8440 18840 8492
rect 18880 8440 18932 8492
rect 20352 8440 20404 8492
rect 7104 8304 7156 8313
rect 1400 8279 1452 8288
rect 1400 8245 1409 8279
rect 1409 8245 1443 8279
rect 1443 8245 1452 8279
rect 1400 8236 1452 8245
rect 3976 8236 4028 8288
rect 5632 8236 5684 8288
rect 6368 8236 6420 8288
rect 6552 8236 6604 8288
rect 8484 8279 8536 8288
rect 8484 8245 8493 8279
rect 8493 8245 8527 8279
rect 8527 8245 8536 8279
rect 8484 8236 8536 8245
rect 8668 8236 8720 8288
rect 8852 8236 8904 8288
rect 9956 8279 10008 8288
rect 9956 8245 9965 8279
rect 9965 8245 9999 8279
rect 9999 8245 10008 8279
rect 9956 8236 10008 8245
rect 10692 8304 10744 8356
rect 11980 8236 12032 8288
rect 16212 8304 16264 8356
rect 16856 8372 16908 8424
rect 18696 8372 18748 8424
rect 19156 8372 19208 8424
rect 20720 8372 20772 8424
rect 14464 8236 14516 8288
rect 15200 8236 15252 8288
rect 15844 8236 15896 8288
rect 16396 8236 16448 8288
rect 17592 8236 17644 8288
rect 20260 8304 20312 8356
rect 21364 8236 21416 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 3976 8032 4028 8084
rect 6000 8032 6052 8084
rect 6184 8032 6236 8084
rect 6460 8032 6512 8084
rect 8300 8032 8352 8084
rect 2596 7939 2648 7948
rect 2596 7905 2630 7939
rect 2630 7905 2648 7939
rect 2596 7896 2648 7905
rect 4252 7896 4304 7948
rect 5448 7939 5500 7948
rect 1768 7692 1820 7744
rect 3976 7828 4028 7880
rect 5448 7905 5457 7939
rect 5457 7905 5491 7939
rect 5491 7905 5500 7939
rect 5448 7896 5500 7905
rect 6276 7939 6328 7948
rect 6276 7905 6285 7939
rect 6285 7905 6319 7939
rect 6319 7905 6328 7939
rect 6276 7896 6328 7905
rect 9128 8032 9180 8084
rect 9956 8032 10008 8084
rect 10048 8032 10100 8084
rect 9680 7964 9732 8016
rect 4344 7760 4396 7812
rect 4804 7760 4856 7812
rect 7472 7896 7524 7948
rect 7656 7896 7708 7948
rect 7840 7896 7892 7948
rect 8208 7939 8260 7948
rect 8208 7905 8242 7939
rect 8242 7905 8260 7939
rect 10324 7964 10376 8016
rect 9956 7939 10008 7948
rect 8208 7896 8260 7905
rect 9956 7905 9965 7939
rect 9965 7905 9999 7939
rect 9999 7905 10008 7939
rect 9956 7896 10008 7905
rect 10600 7939 10652 7948
rect 10600 7905 10609 7939
rect 10609 7905 10643 7939
rect 10643 7905 10652 7939
rect 10600 7896 10652 7905
rect 12164 7964 12216 8016
rect 12348 8032 12400 8084
rect 13820 8032 13872 8084
rect 14372 8032 14424 8084
rect 15016 8032 15068 8084
rect 15292 8075 15344 8084
rect 15292 8041 15301 8075
rect 15301 8041 15335 8075
rect 15335 8041 15344 8075
rect 15292 8032 15344 8041
rect 15660 8032 15712 8084
rect 17684 8032 17736 8084
rect 18880 8032 18932 8084
rect 20076 8032 20128 8084
rect 4068 7692 4120 7744
rect 6000 7692 6052 7744
rect 7288 7692 7340 7744
rect 7380 7692 7432 7744
rect 7748 7828 7800 7880
rect 9496 7828 9548 7880
rect 10508 7828 10560 7880
rect 11980 7896 12032 7948
rect 12440 7896 12492 7948
rect 14648 7964 14700 8016
rect 15108 7964 15160 8016
rect 9220 7760 9272 7812
rect 10416 7760 10468 7812
rect 14096 7896 14148 7948
rect 15476 7896 15528 7948
rect 17592 7896 17644 7948
rect 18052 7896 18104 7948
rect 20076 7939 20128 7948
rect 20076 7905 20085 7939
rect 20085 7905 20119 7939
rect 20119 7905 20128 7939
rect 20076 7896 20128 7905
rect 15016 7828 15068 7880
rect 16028 7828 16080 7880
rect 17040 7871 17092 7880
rect 17040 7837 17049 7871
rect 17049 7837 17083 7871
rect 17083 7837 17092 7871
rect 17040 7828 17092 7837
rect 19708 7828 19760 7880
rect 20168 7871 20220 7880
rect 20168 7837 20177 7871
rect 20177 7837 20211 7871
rect 20211 7837 20220 7871
rect 20168 7828 20220 7837
rect 9128 7692 9180 7744
rect 9312 7692 9364 7744
rect 11980 7735 12032 7744
rect 11980 7701 11989 7735
rect 11989 7701 12023 7735
rect 12023 7701 12032 7735
rect 11980 7692 12032 7701
rect 12716 7692 12768 7744
rect 14188 7692 14240 7744
rect 14924 7735 14976 7744
rect 14924 7701 14933 7735
rect 14933 7701 14967 7735
rect 14967 7701 14976 7735
rect 14924 7692 14976 7701
rect 19064 7760 19116 7812
rect 19616 7760 19668 7812
rect 18604 7692 18656 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 2688 7488 2740 7540
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 4068 7488 4120 7540
rect 5448 7531 5500 7540
rect 5448 7497 5457 7531
rect 5457 7497 5491 7531
rect 5491 7497 5500 7531
rect 5448 7488 5500 7497
rect 6460 7488 6512 7540
rect 7840 7488 7892 7540
rect 8208 7488 8260 7540
rect 8668 7488 8720 7540
rect 9220 7488 9272 7540
rect 9496 7488 9548 7540
rect 9588 7488 9640 7540
rect 11612 7488 11664 7540
rect 5080 7352 5132 7404
rect 13728 7420 13780 7472
rect 14096 7463 14148 7472
rect 6092 7395 6144 7404
rect 6092 7361 6101 7395
rect 6101 7361 6135 7395
rect 6135 7361 6144 7395
rect 6092 7352 6144 7361
rect 8208 7352 8260 7404
rect 8300 7352 8352 7404
rect 9220 7352 9272 7404
rect 9404 7395 9456 7404
rect 9404 7361 9413 7395
rect 9413 7361 9447 7395
rect 9447 7361 9456 7395
rect 9404 7352 9456 7361
rect 10416 7352 10468 7404
rect 10968 7352 11020 7404
rect 6828 7284 6880 7336
rect 7196 7284 7248 7336
rect 7748 7284 7800 7336
rect 7840 7284 7892 7336
rect 8116 7284 8168 7336
rect 2044 7259 2096 7268
rect 2044 7225 2078 7259
rect 2078 7225 2096 7259
rect 4068 7259 4120 7268
rect 2044 7216 2096 7225
rect 4068 7225 4102 7259
rect 4102 7225 4120 7259
rect 4068 7216 4120 7225
rect 5080 7148 5132 7200
rect 6920 7216 6972 7268
rect 8576 7284 8628 7336
rect 11612 7352 11664 7404
rect 12072 7352 12124 7404
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 12440 7352 12492 7361
rect 14096 7429 14105 7463
rect 14105 7429 14139 7463
rect 14139 7429 14148 7463
rect 14096 7420 14148 7429
rect 14372 7352 14424 7404
rect 16028 7488 16080 7540
rect 16212 7488 16264 7540
rect 16856 7488 16908 7540
rect 14924 7420 14976 7472
rect 17776 7488 17828 7540
rect 17868 7488 17920 7540
rect 18512 7488 18564 7540
rect 15200 7352 15252 7404
rect 15384 7352 15436 7404
rect 16488 7352 16540 7404
rect 16856 7395 16908 7404
rect 16856 7361 16865 7395
rect 16865 7361 16899 7395
rect 16899 7361 16908 7395
rect 16856 7352 16908 7361
rect 17960 7420 18012 7472
rect 17684 7352 17736 7404
rect 20168 7488 20220 7540
rect 20536 7420 20588 7472
rect 18880 7352 18932 7404
rect 19708 7395 19760 7404
rect 6000 7148 6052 7200
rect 6368 7148 6420 7200
rect 9036 7216 9088 7268
rect 9404 7216 9456 7268
rect 8852 7148 8904 7200
rect 10508 7216 10560 7268
rect 10416 7148 10468 7200
rect 10876 7191 10928 7200
rect 10876 7157 10885 7191
rect 10885 7157 10919 7191
rect 10919 7157 10928 7191
rect 10876 7148 10928 7157
rect 11060 7216 11112 7268
rect 11428 7216 11480 7268
rect 14648 7284 14700 7336
rect 14188 7216 14240 7268
rect 14372 7216 14424 7268
rect 14556 7259 14608 7268
rect 14556 7225 14565 7259
rect 14565 7225 14599 7259
rect 14599 7225 14608 7259
rect 14556 7216 14608 7225
rect 15108 7216 15160 7268
rect 15476 7216 15528 7268
rect 19340 7284 19392 7336
rect 19708 7361 19717 7395
rect 19717 7361 19751 7395
rect 19751 7361 19760 7395
rect 19708 7352 19760 7361
rect 12164 7148 12216 7200
rect 15292 7148 15344 7200
rect 15660 7148 15712 7200
rect 16212 7148 16264 7200
rect 16580 7148 16632 7200
rect 17224 7148 17276 7200
rect 18696 7148 18748 7200
rect 20628 7216 20680 7268
rect 20444 7191 20496 7200
rect 20444 7157 20453 7191
rect 20453 7157 20487 7191
rect 20487 7157 20496 7191
rect 20444 7148 20496 7157
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 1400 6944 1452 6996
rect 5908 6944 5960 6996
rect 6368 6944 6420 6996
rect 6460 6944 6512 6996
rect 7196 6944 7248 6996
rect 7380 6944 7432 6996
rect 7656 6944 7708 6996
rect 8576 6987 8628 6996
rect 8576 6953 8585 6987
rect 8585 6953 8619 6987
rect 8619 6953 8628 6987
rect 8576 6944 8628 6953
rect 9036 6987 9088 6996
rect 9036 6953 9045 6987
rect 9045 6953 9079 6987
rect 9079 6953 9088 6987
rect 9036 6944 9088 6953
rect 9588 6944 9640 6996
rect 10876 6944 10928 6996
rect 11244 6987 11296 6996
rect 11244 6953 11253 6987
rect 11253 6953 11287 6987
rect 11287 6953 11296 6987
rect 11244 6944 11296 6953
rect 2964 6876 3016 6928
rect 3608 6876 3660 6928
rect 6184 6876 6236 6928
rect 6276 6876 6328 6928
rect 1768 6808 1820 6860
rect 3700 6808 3752 6860
rect 5816 6808 5868 6860
rect 6736 6851 6788 6860
rect 6736 6817 6745 6851
rect 6745 6817 6779 6851
rect 6779 6817 6788 6851
rect 7748 6876 7800 6928
rect 8116 6876 8168 6928
rect 6736 6808 6788 6817
rect 2688 6783 2740 6792
rect 2688 6749 2697 6783
rect 2697 6749 2731 6783
rect 2731 6749 2740 6783
rect 2688 6740 2740 6749
rect 4252 6740 4304 6792
rect 5080 6740 5132 6792
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 5908 6740 5960 6792
rect 6828 6783 6880 6792
rect 6828 6749 6837 6783
rect 6837 6749 6871 6783
rect 6871 6749 6880 6783
rect 6828 6740 6880 6749
rect 7564 6740 7616 6792
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 8668 6876 8720 6928
rect 11520 6876 11572 6928
rect 12164 6944 12216 6996
rect 12808 6944 12860 6996
rect 13176 6944 13228 6996
rect 15476 6944 15528 6996
rect 15660 6987 15712 6996
rect 15660 6953 15669 6987
rect 15669 6953 15703 6987
rect 15703 6953 15712 6987
rect 15660 6944 15712 6953
rect 16856 6944 16908 6996
rect 17040 6944 17092 6996
rect 17868 6987 17920 6996
rect 12072 6876 12124 6928
rect 9496 6808 9548 6860
rect 9588 6740 9640 6792
rect 10416 6783 10468 6792
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 10416 6740 10468 6749
rect 1768 6715 1820 6724
rect 1768 6681 1777 6715
rect 1777 6681 1811 6715
rect 1811 6681 1820 6715
rect 1768 6672 1820 6681
rect 3608 6647 3660 6656
rect 3608 6613 3617 6647
rect 3617 6613 3651 6647
rect 3651 6613 3660 6647
rect 3608 6604 3660 6613
rect 3976 6604 4028 6656
rect 11060 6672 11112 6724
rect 11428 6740 11480 6792
rect 11612 6808 11664 6860
rect 11888 6808 11940 6860
rect 12900 6876 12952 6928
rect 13084 6876 13136 6928
rect 14188 6876 14240 6928
rect 14372 6876 14424 6928
rect 15108 6876 15160 6928
rect 15752 6876 15804 6928
rect 17224 6919 17276 6928
rect 12532 6808 12584 6860
rect 13912 6808 13964 6860
rect 17224 6885 17233 6919
rect 17233 6885 17267 6919
rect 17267 6885 17276 6919
rect 17224 6876 17276 6885
rect 17868 6953 17877 6987
rect 17877 6953 17911 6987
rect 17911 6953 17920 6987
rect 17868 6944 17920 6953
rect 18236 6987 18288 6996
rect 18236 6953 18245 6987
rect 18245 6953 18279 6987
rect 18279 6953 18288 6987
rect 18236 6944 18288 6953
rect 18328 6987 18380 6996
rect 18328 6953 18337 6987
rect 18337 6953 18371 6987
rect 18371 6953 18380 6987
rect 18328 6944 18380 6953
rect 18512 6944 18564 6996
rect 18696 6944 18748 6996
rect 18788 6944 18840 6996
rect 19340 6944 19392 6996
rect 11980 6740 12032 6792
rect 13176 6740 13228 6792
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 14096 6783 14148 6792
rect 14096 6749 14105 6783
rect 14105 6749 14139 6783
rect 14139 6749 14148 6783
rect 14096 6740 14148 6749
rect 15384 6740 15436 6792
rect 6000 6604 6052 6656
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 8024 6604 8076 6656
rect 9220 6604 9272 6656
rect 9312 6604 9364 6656
rect 9772 6604 9824 6656
rect 10692 6604 10744 6656
rect 11612 6604 11664 6656
rect 13360 6604 13412 6656
rect 13544 6604 13596 6656
rect 16028 6740 16080 6792
rect 17684 6808 17736 6860
rect 19524 6876 19576 6928
rect 18328 6740 18380 6792
rect 19248 6808 19300 6860
rect 21088 6808 21140 6860
rect 19156 6783 19208 6792
rect 19156 6749 19165 6783
rect 19165 6749 19199 6783
rect 19199 6749 19208 6783
rect 19156 6740 19208 6749
rect 15108 6604 15160 6656
rect 17684 6672 17736 6724
rect 16764 6604 16816 6656
rect 17408 6604 17460 6656
rect 17592 6604 17644 6656
rect 20260 6604 20312 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 2136 6400 2188 6452
rect 4252 6400 4304 6452
rect 13268 6400 13320 6452
rect 13360 6400 13412 6452
rect 14004 6443 14056 6452
rect 1768 6332 1820 6384
rect 2320 6332 2372 6384
rect 3608 6332 3660 6384
rect 4068 6332 4120 6384
rect 2228 6264 2280 6316
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 3792 6264 3844 6316
rect 4712 6307 4764 6316
rect 4712 6273 4721 6307
rect 4721 6273 4755 6307
rect 4755 6273 4764 6307
rect 4712 6264 4764 6273
rect 6276 6332 6328 6384
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 6644 6332 6696 6384
rect 7656 6375 7708 6384
rect 7656 6341 7665 6375
rect 7665 6341 7699 6375
rect 7699 6341 7708 6375
rect 7656 6332 7708 6341
rect 8024 6332 8076 6384
rect 8116 6332 8168 6384
rect 5724 6264 5776 6273
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 6828 6264 6880 6316
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 7932 6196 7984 6248
rect 9036 6332 9088 6384
rect 8576 6264 8628 6316
rect 11060 6332 11112 6384
rect 11888 6332 11940 6384
rect 8392 6196 8444 6248
rect 9220 6239 9272 6248
rect 9220 6205 9229 6239
rect 9229 6205 9263 6239
rect 9263 6205 9272 6239
rect 9220 6196 9272 6205
rect 11980 6264 12032 6316
rect 14004 6409 14013 6443
rect 14013 6409 14047 6443
rect 14047 6409 14056 6443
rect 14004 6400 14056 6409
rect 17500 6400 17552 6452
rect 19248 6400 19300 6452
rect 13912 6332 13964 6384
rect 14372 6332 14424 6384
rect 16028 6332 16080 6384
rect 17408 6307 17460 6316
rect 17408 6273 17417 6307
rect 17417 6273 17451 6307
rect 17451 6273 17460 6307
rect 17408 6264 17460 6273
rect 17960 6264 18012 6316
rect 18328 6264 18380 6316
rect 6092 6128 6144 6180
rect 1952 6103 2004 6112
rect 1952 6069 1961 6103
rect 1961 6069 1995 6103
rect 1995 6069 2004 6103
rect 1952 6060 2004 6069
rect 2320 6103 2372 6112
rect 2320 6069 2329 6103
rect 2329 6069 2363 6103
rect 2363 6069 2372 6103
rect 2320 6060 2372 6069
rect 2412 6103 2464 6112
rect 2412 6069 2421 6103
rect 2421 6069 2455 6103
rect 2455 6069 2464 6103
rect 3240 6103 3292 6112
rect 2412 6060 2464 6069
rect 3240 6069 3249 6103
rect 3249 6069 3283 6103
rect 3283 6069 3292 6103
rect 3240 6060 3292 6069
rect 4068 6103 4120 6112
rect 4068 6069 4077 6103
rect 4077 6069 4111 6103
rect 4111 6069 4120 6103
rect 4068 6060 4120 6069
rect 6644 6060 6696 6112
rect 7380 6060 7432 6112
rect 7748 6060 7800 6112
rect 8024 6128 8076 6180
rect 8576 6128 8628 6180
rect 9496 6128 9548 6180
rect 9312 6060 9364 6112
rect 11888 6128 11940 6180
rect 12532 6196 12584 6248
rect 13820 6196 13872 6248
rect 14464 6239 14516 6248
rect 14464 6205 14473 6239
rect 14473 6205 14507 6239
rect 14507 6205 14516 6239
rect 14464 6196 14516 6205
rect 11060 6060 11112 6112
rect 12808 6060 12860 6112
rect 12992 6128 13044 6180
rect 15384 6128 15436 6180
rect 17592 6196 17644 6248
rect 17960 6128 18012 6180
rect 18880 6196 18932 6248
rect 19156 6196 19208 6248
rect 20444 6196 20496 6248
rect 20260 6128 20312 6180
rect 14096 6060 14148 6112
rect 15200 6060 15252 6112
rect 17776 6060 17828 6112
rect 18052 6103 18104 6112
rect 18052 6069 18061 6103
rect 18061 6069 18095 6103
rect 18095 6069 18104 6103
rect 18052 6060 18104 6069
rect 18328 6060 18380 6112
rect 20812 6060 20864 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 3700 5856 3752 5908
rect 1400 5788 1452 5840
rect 1952 5720 2004 5772
rect 1860 5652 1912 5704
rect 3884 5720 3936 5772
rect 4712 5788 4764 5840
rect 6092 5856 6144 5908
rect 6184 5856 6236 5908
rect 7288 5856 7340 5908
rect 8576 5899 8628 5908
rect 5540 5788 5592 5840
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 9312 5856 9364 5908
rect 6460 5720 6512 5772
rect 5724 5652 5776 5704
rect 5540 5584 5592 5636
rect 6092 5584 6144 5636
rect 7288 5720 7340 5772
rect 7380 5720 7432 5772
rect 6736 5695 6788 5704
rect 6736 5661 6745 5695
rect 6745 5661 6779 5695
rect 6779 5661 6788 5695
rect 6736 5652 6788 5661
rect 7012 5652 7064 5704
rect 8392 5652 8444 5704
rect 9036 5720 9088 5772
rect 11060 5788 11112 5840
rect 12348 5856 12400 5908
rect 12808 5856 12860 5908
rect 12992 5788 13044 5840
rect 13360 5831 13412 5840
rect 13360 5797 13394 5831
rect 13394 5797 13412 5831
rect 14096 5856 14148 5908
rect 15016 5856 15068 5908
rect 16120 5856 16172 5908
rect 18052 5856 18104 5908
rect 19800 5899 19852 5908
rect 19800 5865 19809 5899
rect 19809 5865 19843 5899
rect 19843 5865 19852 5899
rect 19800 5856 19852 5865
rect 20628 5856 20680 5908
rect 13360 5788 13412 5797
rect 11612 5720 11664 5772
rect 12348 5720 12400 5772
rect 12624 5720 12676 5772
rect 13176 5720 13228 5772
rect 14188 5720 14240 5772
rect 15108 5720 15160 5772
rect 19892 5831 19944 5840
rect 19892 5797 19901 5831
rect 19901 5797 19935 5831
rect 19935 5797 19944 5831
rect 19892 5788 19944 5797
rect 21272 5788 21324 5840
rect 15752 5720 15804 5772
rect 16856 5720 16908 5772
rect 17040 5763 17092 5772
rect 17040 5729 17074 5763
rect 17074 5729 17092 5763
rect 17040 5720 17092 5729
rect 18328 5720 18380 5772
rect 20444 5720 20496 5772
rect 8116 5584 8168 5636
rect 3516 5516 3568 5568
rect 3884 5516 3936 5568
rect 5080 5516 5132 5568
rect 7012 5516 7064 5568
rect 7840 5516 7892 5568
rect 12164 5652 12216 5704
rect 10692 5584 10744 5636
rect 12624 5584 12676 5636
rect 13084 5584 13136 5636
rect 14464 5627 14516 5636
rect 14464 5593 14473 5627
rect 14473 5593 14507 5627
rect 14507 5593 14516 5627
rect 14464 5584 14516 5593
rect 15200 5652 15252 5704
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 16028 5652 16080 5661
rect 18144 5652 18196 5704
rect 19524 5652 19576 5704
rect 16580 5584 16632 5636
rect 17776 5584 17828 5636
rect 9588 5516 9640 5568
rect 10416 5516 10468 5568
rect 11152 5516 11204 5568
rect 12164 5516 12216 5568
rect 12992 5516 13044 5568
rect 13728 5516 13780 5568
rect 17500 5516 17552 5568
rect 17684 5516 17736 5568
rect 18696 5516 18748 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 1584 5355 1636 5364
rect 1584 5321 1593 5355
rect 1593 5321 1627 5355
rect 1627 5321 1636 5355
rect 1584 5312 1636 5321
rect 3240 5312 3292 5364
rect 4896 5312 4948 5364
rect 5264 5312 5316 5364
rect 7196 5312 7248 5364
rect 8208 5355 8260 5364
rect 8208 5321 8217 5355
rect 8217 5321 8251 5355
rect 8251 5321 8260 5355
rect 8208 5312 8260 5321
rect 3332 5244 3384 5296
rect 6276 5244 6328 5296
rect 1860 5176 1912 5228
rect 3884 5176 3936 5228
rect 4712 5176 4764 5228
rect 3700 5108 3752 5160
rect 4068 5108 4120 5160
rect 4252 5108 4304 5160
rect 5080 5108 5132 5160
rect 6000 5108 6052 5160
rect 6184 5151 6236 5160
rect 6184 5117 6193 5151
rect 6193 5117 6227 5151
rect 6227 5117 6236 5151
rect 6184 5108 6236 5117
rect 2228 5083 2280 5092
rect 2228 5049 2262 5083
rect 2262 5049 2280 5083
rect 2228 5040 2280 5049
rect 4344 5040 4396 5092
rect 5540 5040 5592 5092
rect 8116 5176 8168 5228
rect 8668 5176 8720 5228
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 9036 5312 9088 5364
rect 9128 5312 9180 5364
rect 10692 5312 10744 5364
rect 12440 5312 12492 5364
rect 14556 5312 14608 5364
rect 12164 5176 12216 5228
rect 12992 5176 13044 5228
rect 13360 5176 13412 5228
rect 14556 5176 14608 5228
rect 14648 5176 14700 5228
rect 15384 5219 15436 5228
rect 15384 5185 15393 5219
rect 15393 5185 15427 5219
rect 15427 5185 15436 5219
rect 16856 5312 16908 5364
rect 17040 5312 17092 5364
rect 17960 5312 18012 5364
rect 19064 5312 19116 5364
rect 20260 5355 20312 5364
rect 15384 5176 15436 5185
rect 20260 5321 20269 5355
rect 20269 5321 20303 5355
rect 20303 5321 20312 5355
rect 20260 5312 20312 5321
rect 6828 5108 6880 5117
rect 9588 5108 9640 5160
rect 10140 5108 10192 5160
rect 6736 5040 6788 5092
rect 7104 5083 7156 5092
rect 7104 5049 7138 5083
rect 7138 5049 7156 5083
rect 7104 5040 7156 5049
rect 7472 5040 7524 5092
rect 8852 5040 8904 5092
rect 3608 4972 3660 5024
rect 9404 5040 9456 5092
rect 11612 5040 11664 5092
rect 18880 5151 18932 5160
rect 15844 5040 15896 5092
rect 16028 5040 16080 5092
rect 18880 5117 18889 5151
rect 18889 5117 18923 5151
rect 18923 5117 18932 5151
rect 18880 5108 18932 5117
rect 20076 5108 20128 5160
rect 20536 5151 20588 5160
rect 20536 5117 20545 5151
rect 20545 5117 20579 5151
rect 20579 5117 20588 5151
rect 20536 5108 20588 5117
rect 18788 5040 18840 5092
rect 19708 5040 19760 5092
rect 9036 4972 9088 5024
rect 10048 4972 10100 5024
rect 10416 4972 10468 5024
rect 10784 4972 10836 5024
rect 10876 4972 10928 5024
rect 11428 5015 11480 5024
rect 11428 4981 11437 5015
rect 11437 4981 11471 5015
rect 11471 4981 11480 5015
rect 11428 4972 11480 4981
rect 12440 5015 12492 5024
rect 12440 4981 12449 5015
rect 12449 4981 12483 5015
rect 12483 4981 12492 5015
rect 12440 4972 12492 4981
rect 13268 5015 13320 5024
rect 13268 4981 13277 5015
rect 13277 4981 13311 5015
rect 13311 4981 13320 5015
rect 13268 4972 13320 4981
rect 13912 4972 13964 5024
rect 14096 5015 14148 5024
rect 14096 4981 14105 5015
rect 14105 4981 14139 5015
rect 14139 4981 14148 5015
rect 14096 4972 14148 4981
rect 14188 5015 14240 5024
rect 14188 4981 14197 5015
rect 14197 4981 14231 5015
rect 14231 4981 14240 5015
rect 14188 4972 14240 4981
rect 15200 4972 15252 5024
rect 18512 4972 18564 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 2228 4768 2280 4820
rect 3332 4811 3384 4820
rect 3332 4777 3341 4811
rect 3341 4777 3375 4811
rect 3375 4777 3384 4811
rect 3332 4768 3384 4777
rect 3700 4768 3752 4820
rect 4988 4768 5040 4820
rect 5172 4768 5224 4820
rect 7104 4811 7156 4820
rect 1860 4700 1912 4752
rect 2228 4632 2280 4684
rect 2872 4632 2924 4684
rect 3608 4607 3660 4616
rect 3608 4573 3617 4607
rect 3617 4573 3651 4607
rect 3651 4573 3660 4607
rect 3608 4564 3660 4573
rect 4252 4632 4304 4684
rect 4712 4632 4764 4684
rect 5448 4632 5500 4684
rect 3148 4496 3200 4548
rect 5172 4564 5224 4616
rect 5908 4700 5960 4752
rect 6276 4700 6328 4752
rect 7104 4777 7113 4811
rect 7113 4777 7147 4811
rect 7147 4777 7156 4811
rect 7104 4768 7156 4777
rect 7380 4811 7432 4820
rect 7380 4777 7389 4811
rect 7389 4777 7423 4811
rect 7423 4777 7432 4811
rect 7380 4768 7432 4777
rect 7748 4811 7800 4820
rect 7748 4777 7757 4811
rect 7757 4777 7791 4811
rect 7791 4777 7800 4811
rect 7748 4768 7800 4777
rect 8852 4768 8904 4820
rect 10140 4811 10192 4820
rect 10140 4777 10149 4811
rect 10149 4777 10183 4811
rect 10183 4777 10192 4811
rect 10140 4768 10192 4777
rect 10876 4811 10928 4820
rect 10416 4700 10468 4752
rect 10876 4777 10885 4811
rect 10885 4777 10919 4811
rect 10919 4777 10928 4811
rect 10876 4768 10928 4777
rect 11152 4768 11204 4820
rect 11428 4768 11480 4820
rect 12072 4768 12124 4820
rect 12440 4768 12492 4820
rect 13912 4811 13964 4820
rect 13912 4777 13921 4811
rect 13921 4777 13955 4811
rect 13955 4777 13964 4811
rect 13912 4768 13964 4777
rect 15200 4768 15252 4820
rect 16028 4768 16080 4820
rect 13084 4700 13136 4752
rect 17224 4768 17276 4820
rect 17776 4811 17828 4820
rect 17776 4777 17785 4811
rect 17785 4777 17819 4811
rect 17819 4777 17828 4811
rect 17776 4768 17828 4777
rect 5724 4675 5776 4684
rect 5724 4641 5733 4675
rect 5733 4641 5767 4675
rect 5767 4641 5776 4675
rect 5724 4632 5776 4641
rect 9680 4632 9732 4684
rect 10876 4632 10928 4684
rect 8392 4564 8444 4616
rect 11060 4607 11112 4616
rect 11060 4573 11069 4607
rect 11069 4573 11103 4607
rect 11103 4573 11112 4607
rect 11060 4564 11112 4573
rect 12164 4607 12216 4616
rect 5632 4496 5684 4548
rect 7656 4496 7708 4548
rect 8300 4496 8352 4548
rect 8852 4496 8904 4548
rect 11428 4496 11480 4548
rect 12164 4573 12173 4607
rect 12173 4573 12207 4607
rect 12207 4573 12216 4607
rect 12164 4564 12216 4573
rect 14280 4632 14332 4684
rect 14740 4632 14792 4684
rect 16212 4632 16264 4684
rect 18696 4700 18748 4752
rect 14188 4564 14240 4616
rect 14464 4564 14516 4616
rect 16028 4564 16080 4616
rect 16856 4607 16908 4616
rect 16856 4573 16865 4607
rect 16865 4573 16899 4607
rect 16899 4573 16908 4607
rect 16856 4564 16908 4573
rect 17040 4607 17092 4616
rect 17040 4573 17049 4607
rect 17049 4573 17083 4607
rect 17083 4573 17092 4607
rect 17040 4564 17092 4573
rect 18788 4632 18840 4684
rect 19524 4675 19576 4684
rect 19524 4641 19533 4675
rect 19533 4641 19567 4675
rect 19567 4641 19576 4675
rect 19524 4632 19576 4641
rect 19800 4632 19852 4684
rect 19616 4607 19668 4616
rect 19616 4573 19625 4607
rect 19625 4573 19659 4607
rect 19659 4573 19668 4607
rect 19616 4564 19668 4573
rect 19708 4607 19760 4616
rect 19708 4573 19717 4607
rect 19717 4573 19751 4607
rect 19751 4573 19760 4607
rect 19708 4564 19760 4573
rect 19892 4564 19944 4616
rect 20168 4496 20220 4548
rect 3976 4428 4028 4480
rect 10968 4428 11020 4480
rect 11704 4428 11756 4480
rect 12900 4428 12952 4480
rect 13084 4428 13136 4480
rect 14832 4471 14884 4480
rect 14832 4437 14841 4471
rect 14841 4437 14875 4471
rect 14875 4437 14884 4471
rect 14832 4428 14884 4437
rect 15108 4428 15160 4480
rect 15660 4428 15712 4480
rect 17316 4428 17368 4480
rect 17408 4428 17460 4480
rect 20076 4428 20128 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 3608 4224 3660 4276
rect 13728 4224 13780 4276
rect 14832 4224 14884 4276
rect 17776 4224 17828 4276
rect 6000 4156 6052 4208
rect 6368 4156 6420 4208
rect 6736 4156 6788 4208
rect 2228 4131 2280 4140
rect 2228 4097 2237 4131
rect 2237 4097 2271 4131
rect 2271 4097 2280 4131
rect 2228 4088 2280 4097
rect 3148 4131 3200 4140
rect 3148 4097 3157 4131
rect 3157 4097 3191 4131
rect 3191 4097 3200 4131
rect 3148 4088 3200 4097
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 5172 4088 5224 4140
rect 4344 4020 4396 4072
rect 5724 4020 5776 4072
rect 6552 4020 6604 4072
rect 2412 3884 2464 3936
rect 4896 3952 4948 4004
rect 5264 3952 5316 4004
rect 6000 3952 6052 4004
rect 7012 4088 7064 4140
rect 8208 4156 8260 4208
rect 8300 4199 8352 4208
rect 8300 4165 8309 4199
rect 8309 4165 8343 4199
rect 8343 4165 8352 4199
rect 8300 4156 8352 4165
rect 9864 4156 9916 4208
rect 10324 4156 10376 4208
rect 7196 4063 7248 4072
rect 7196 4029 7205 4063
rect 7205 4029 7239 4063
rect 7239 4029 7248 4063
rect 7196 4020 7248 4029
rect 7564 4020 7616 4072
rect 8208 4020 8260 4072
rect 11704 4131 11756 4140
rect 11704 4097 11713 4131
rect 11713 4097 11747 4131
rect 11747 4097 11756 4131
rect 11704 4088 11756 4097
rect 11888 4156 11940 4208
rect 12072 4088 12124 4140
rect 13084 4156 13136 4208
rect 14188 4156 14240 4208
rect 14556 4156 14608 4208
rect 15200 4088 15252 4140
rect 17684 4156 17736 4208
rect 10692 4020 10744 4072
rect 11888 4020 11940 4072
rect 10600 3995 10652 4004
rect 10600 3961 10609 3995
rect 10609 3961 10643 3995
rect 10643 3961 10652 3995
rect 12808 4020 12860 4072
rect 13176 4020 13228 4072
rect 10600 3952 10652 3961
rect 3700 3927 3752 3936
rect 3700 3893 3709 3927
rect 3709 3893 3743 3927
rect 3743 3893 3752 3927
rect 3700 3884 3752 3893
rect 3884 3884 3936 3936
rect 4160 3927 4212 3936
rect 4160 3893 4169 3927
rect 4169 3893 4203 3927
rect 4203 3893 4212 3927
rect 4160 3884 4212 3893
rect 4804 3884 4856 3936
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 9864 3884 9916 3936
rect 10232 3884 10284 3936
rect 10324 3884 10376 3936
rect 12624 3952 12676 4004
rect 16028 4088 16080 4140
rect 17960 4088 18012 4140
rect 18052 4131 18104 4140
rect 18052 4097 18061 4131
rect 18061 4097 18095 4131
rect 18095 4097 18104 4131
rect 20536 4224 20588 4276
rect 20260 4156 20312 4208
rect 20904 4199 20956 4208
rect 18052 4088 18104 4097
rect 19984 4088 20036 4140
rect 20904 4165 20913 4199
rect 20913 4165 20947 4199
rect 20947 4165 20956 4199
rect 20904 4156 20956 4165
rect 13360 3995 13412 4004
rect 13360 3961 13394 3995
rect 13394 3961 13412 3995
rect 13360 3952 13412 3961
rect 14096 3952 14148 4004
rect 19800 4020 19852 4072
rect 20536 4020 20588 4072
rect 11520 3884 11572 3936
rect 12440 3884 12492 3936
rect 12808 3884 12860 3936
rect 14004 3884 14056 3936
rect 15108 3927 15160 3936
rect 15108 3893 15117 3927
rect 15117 3893 15151 3927
rect 15151 3893 15160 3927
rect 15108 3884 15160 3893
rect 15200 3927 15252 3936
rect 15200 3893 15209 3927
rect 15209 3893 15243 3927
rect 15243 3893 15252 3927
rect 15200 3884 15252 3893
rect 16304 3927 16356 3936
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 16672 3927 16724 3936
rect 16304 3884 16356 3893
rect 16672 3893 16681 3927
rect 16681 3893 16715 3927
rect 16715 3893 16724 3927
rect 16672 3884 16724 3893
rect 16948 3884 17000 3936
rect 17040 3884 17092 3936
rect 20352 3952 20404 4004
rect 19340 3884 19392 3936
rect 19708 3884 19760 3936
rect 19984 3884 20036 3936
rect 20076 3927 20128 3936
rect 20076 3893 20085 3927
rect 20085 3893 20119 3927
rect 20119 3893 20128 3927
rect 20076 3884 20128 3893
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 2044 3723 2096 3732
rect 2044 3689 2053 3723
rect 2053 3689 2087 3723
rect 2087 3689 2096 3723
rect 2044 3680 2096 3689
rect 2228 3680 2280 3732
rect 3608 3680 3660 3732
rect 3884 3680 3936 3732
rect 4252 3680 4304 3732
rect 4988 3680 5040 3732
rect 7012 3723 7064 3732
rect 7012 3689 7021 3723
rect 7021 3689 7055 3723
rect 7055 3689 7064 3723
rect 7012 3680 7064 3689
rect 9680 3723 9732 3732
rect 1676 3655 1728 3664
rect 1676 3621 1685 3655
rect 1685 3621 1719 3655
rect 1719 3621 1728 3655
rect 1676 3612 1728 3621
rect 7104 3655 7156 3664
rect 1860 3544 1912 3596
rect 3332 3544 3384 3596
rect 4160 3544 4212 3596
rect 6368 3544 6420 3596
rect 5172 3476 5224 3528
rect 4160 3408 4212 3460
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 7104 3621 7113 3655
rect 7113 3621 7147 3655
rect 7147 3621 7156 3655
rect 7104 3612 7156 3621
rect 7288 3612 7340 3664
rect 7380 3612 7432 3664
rect 8024 3655 8076 3664
rect 8024 3621 8033 3655
rect 8033 3621 8067 3655
rect 8067 3621 8076 3655
rect 8024 3612 8076 3621
rect 8944 3612 8996 3664
rect 8484 3544 8536 3596
rect 9680 3689 9689 3723
rect 9689 3689 9723 3723
rect 9723 3689 9732 3723
rect 9680 3680 9732 3689
rect 9772 3680 9824 3732
rect 9956 3612 10008 3664
rect 10692 3680 10744 3732
rect 12440 3723 12492 3732
rect 12440 3689 12449 3723
rect 12449 3689 12483 3723
rect 12483 3689 12492 3723
rect 12440 3680 12492 3689
rect 11060 3655 11112 3664
rect 11060 3621 11094 3655
rect 11094 3621 11112 3655
rect 11060 3612 11112 3621
rect 11244 3612 11296 3664
rect 12900 3655 12952 3664
rect 12900 3621 12909 3655
rect 12909 3621 12943 3655
rect 12943 3621 12952 3655
rect 12900 3612 12952 3621
rect 8392 3476 8444 3528
rect 8576 3476 8628 3528
rect 9772 3476 9824 3528
rect 9956 3476 10008 3528
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 10692 3476 10744 3528
rect 10600 3408 10652 3460
rect 13176 3544 13228 3596
rect 12808 3476 12860 3528
rect 15108 3612 15160 3664
rect 18052 3680 18104 3732
rect 16856 3612 16908 3664
rect 17592 3612 17644 3664
rect 17960 3612 18012 3664
rect 18696 3612 18748 3664
rect 19248 3612 19300 3664
rect 20352 3612 20404 3664
rect 14096 3544 14148 3596
rect 14832 3587 14884 3596
rect 14832 3553 14841 3587
rect 14841 3553 14875 3587
rect 14875 3553 14884 3587
rect 14832 3544 14884 3553
rect 15292 3544 15344 3596
rect 16580 3544 16632 3596
rect 13912 3519 13964 3528
rect 13912 3485 13921 3519
rect 13921 3485 13955 3519
rect 13955 3485 13964 3519
rect 13912 3476 13964 3485
rect 14188 3476 14240 3528
rect 16028 3476 16080 3528
rect 16488 3476 16540 3528
rect 18236 3544 18288 3596
rect 18972 3544 19024 3596
rect 18788 3476 18840 3528
rect 18880 3476 18932 3528
rect 19248 3519 19300 3528
rect 19248 3485 19257 3519
rect 19257 3485 19291 3519
rect 19291 3485 19300 3519
rect 19248 3476 19300 3485
rect 19340 3519 19392 3528
rect 19340 3485 19349 3519
rect 19349 3485 19383 3519
rect 19383 3485 19392 3519
rect 19340 3476 19392 3485
rect 20076 3476 20128 3528
rect 5264 3383 5316 3392
rect 5264 3349 5273 3383
rect 5273 3349 5307 3383
rect 5307 3349 5316 3383
rect 5264 3340 5316 3349
rect 5448 3383 5500 3392
rect 5448 3349 5457 3383
rect 5457 3349 5491 3383
rect 5491 3349 5500 3383
rect 5448 3340 5500 3349
rect 6092 3340 6144 3392
rect 6920 3340 6972 3392
rect 7656 3340 7708 3392
rect 8300 3340 8352 3392
rect 12164 3383 12216 3392
rect 12164 3349 12173 3383
rect 12173 3349 12207 3383
rect 12207 3349 12216 3383
rect 12164 3340 12216 3349
rect 14556 3340 14608 3392
rect 19616 3408 19668 3460
rect 17868 3340 17920 3392
rect 19708 3340 19760 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 1860 3136 1912 3188
rect 2320 3068 2372 3120
rect 2228 3043 2280 3052
rect 2228 3009 2237 3043
rect 2237 3009 2271 3043
rect 2271 3009 2280 3043
rect 2228 3000 2280 3009
rect 3700 3068 3752 3120
rect 3332 3043 3384 3052
rect 3332 3009 3341 3043
rect 3341 3009 3375 3043
rect 3375 3009 3384 3043
rect 3332 3000 3384 3009
rect 6184 3136 6236 3188
rect 6276 3136 6328 3188
rect 8208 3179 8260 3188
rect 8208 3145 8217 3179
rect 8217 3145 8251 3179
rect 8251 3145 8260 3179
rect 8208 3136 8260 3145
rect 8852 3136 8904 3188
rect 5264 3111 5316 3120
rect 5264 3077 5273 3111
rect 5273 3077 5307 3111
rect 5307 3077 5316 3111
rect 5264 3068 5316 3077
rect 6000 3068 6052 3120
rect 9956 3068 10008 3120
rect 10508 3068 10560 3120
rect 12072 3111 12124 3120
rect 12072 3077 12081 3111
rect 12081 3077 12115 3111
rect 12115 3077 12124 3111
rect 12072 3068 12124 3077
rect 12440 3111 12492 3120
rect 12440 3077 12449 3111
rect 12449 3077 12483 3111
rect 12483 3077 12492 3111
rect 12440 3068 12492 3077
rect 3792 2932 3844 2984
rect 6276 3043 6328 3052
rect 6276 3009 6285 3043
rect 6285 3009 6319 3043
rect 6319 3009 6328 3043
rect 6276 3000 6328 3009
rect 7840 3000 7892 3052
rect 8116 3000 8168 3052
rect 4436 2932 4488 2984
rect 5356 2975 5408 2984
rect 5356 2941 5365 2975
rect 5365 2941 5399 2975
rect 5399 2941 5408 2975
rect 5356 2932 5408 2941
rect 6092 2975 6144 2984
rect 6092 2941 6101 2975
rect 6101 2941 6135 2975
rect 6135 2941 6144 2975
rect 6092 2932 6144 2941
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 6828 2932 6880 2941
rect 5172 2864 5224 2916
rect 2044 2839 2096 2848
rect 2044 2805 2053 2839
rect 2053 2805 2087 2839
rect 2087 2805 2096 2839
rect 2044 2796 2096 2805
rect 3056 2839 3108 2848
rect 3056 2805 3065 2839
rect 3065 2805 3099 2839
rect 3099 2805 3108 2839
rect 3056 2796 3108 2805
rect 3700 2839 3752 2848
rect 3700 2805 3709 2839
rect 3709 2805 3743 2839
rect 3743 2805 3752 2839
rect 3700 2796 3752 2805
rect 10232 3000 10284 3052
rect 10692 3043 10744 3052
rect 10692 3009 10701 3043
rect 10701 3009 10735 3043
rect 10735 3009 10744 3043
rect 10692 3000 10744 3009
rect 11796 3000 11848 3052
rect 13084 3043 13136 3052
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 14280 3068 14332 3120
rect 14096 3043 14148 3052
rect 14096 3009 14105 3043
rect 14105 3009 14139 3043
rect 14139 3009 14148 3043
rect 14096 3000 14148 3009
rect 14924 3043 14976 3052
rect 14924 3009 14933 3043
rect 14933 3009 14967 3043
rect 14967 3009 14976 3043
rect 14924 3000 14976 3009
rect 10324 2932 10376 2984
rect 12164 2932 12216 2984
rect 12716 2932 12768 2984
rect 12808 2975 12860 2984
rect 12808 2941 12817 2975
rect 12817 2941 12851 2975
rect 12851 2941 12860 2975
rect 13452 2975 13504 2984
rect 12808 2932 12860 2941
rect 13452 2941 13461 2975
rect 13461 2941 13495 2975
rect 13495 2941 13504 2975
rect 13452 2932 13504 2941
rect 17040 3136 17092 3188
rect 19524 3179 19576 3188
rect 16948 3068 17000 3120
rect 17684 3068 17736 3120
rect 17868 3068 17920 3120
rect 19524 3145 19533 3179
rect 19533 3145 19567 3179
rect 19567 3145 19576 3179
rect 19524 3136 19576 3145
rect 17224 3000 17276 3052
rect 16488 2932 16540 2984
rect 18696 3000 18748 3052
rect 19248 3000 19300 3052
rect 20076 3043 20128 3052
rect 20076 3009 20085 3043
rect 20085 3009 20119 3043
rect 20119 3009 20128 3043
rect 20076 3000 20128 3009
rect 19892 2975 19944 2984
rect 19892 2941 19901 2975
rect 19901 2941 19935 2975
rect 19935 2941 19944 2975
rect 19892 2932 19944 2941
rect 6184 2839 6236 2848
rect 6184 2805 6193 2839
rect 6193 2805 6227 2839
rect 6227 2805 6236 2839
rect 6184 2796 6236 2805
rect 6828 2796 6880 2848
rect 7748 2796 7800 2848
rect 11152 2864 11204 2916
rect 8392 2796 8444 2848
rect 8576 2796 8628 2848
rect 14740 2907 14792 2916
rect 14740 2873 14749 2907
rect 14749 2873 14783 2907
rect 14783 2873 14792 2907
rect 14740 2864 14792 2873
rect 15016 2864 15068 2916
rect 16028 2864 16080 2916
rect 16212 2864 16264 2916
rect 22192 2864 22244 2916
rect 14464 2796 14516 2848
rect 16488 2796 16540 2848
rect 17960 2796 18012 2848
rect 19156 2796 19208 2848
rect 20628 2796 20680 2848
rect 22560 2796 22612 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 2044 2592 2096 2644
rect 2688 2592 2740 2644
rect 2596 2524 2648 2576
rect 3332 2592 3384 2644
rect 5264 2592 5316 2644
rect 5816 2592 5868 2644
rect 6184 2592 6236 2644
rect 7748 2592 7800 2644
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 8668 2592 8720 2644
rect 3148 2524 3200 2576
rect 5448 2524 5500 2576
rect 6092 2524 6144 2576
rect 6644 2524 6696 2576
rect 7656 2524 7708 2576
rect 10324 2592 10376 2644
rect 10508 2592 10560 2644
rect 12808 2592 12860 2644
rect 12992 2635 13044 2644
rect 12992 2601 13001 2635
rect 13001 2601 13035 2635
rect 13035 2601 13044 2635
rect 12992 2592 13044 2601
rect 15936 2592 15988 2644
rect 17132 2592 17184 2644
rect 17500 2592 17552 2644
rect 1952 2456 2004 2508
rect 3424 2456 3476 2508
rect 4436 2499 4488 2508
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 3700 2388 3752 2440
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 4436 2465 4445 2499
rect 4445 2465 4479 2499
rect 4479 2465 4488 2499
rect 4436 2456 4488 2465
rect 4988 2456 5040 2508
rect 7196 2456 7248 2508
rect 9128 2499 9180 2508
rect 3792 2388 3844 2397
rect 5540 2388 5592 2440
rect 7380 2431 7432 2440
rect 7380 2397 7389 2431
rect 7389 2397 7423 2431
rect 7423 2397 7432 2431
rect 7380 2388 7432 2397
rect 9128 2465 9137 2499
rect 9137 2465 9171 2499
rect 9171 2465 9180 2499
rect 9128 2456 9180 2465
rect 9956 2456 10008 2508
rect 10140 2499 10192 2508
rect 10140 2465 10149 2499
rect 10149 2465 10183 2499
rect 10183 2465 10192 2499
rect 10140 2456 10192 2465
rect 10324 2456 10376 2508
rect 8300 2388 8352 2440
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 11612 2456 11664 2508
rect 16396 2524 16448 2576
rect 16856 2524 16908 2576
rect 17592 2567 17644 2576
rect 17592 2533 17601 2567
rect 17601 2533 17635 2567
rect 17635 2533 17644 2567
rect 17592 2524 17644 2533
rect 12256 2456 12308 2508
rect 4160 2320 4212 2372
rect 4344 2363 4396 2372
rect 4344 2329 4353 2363
rect 4353 2329 4387 2363
rect 4387 2329 4396 2363
rect 4344 2320 4396 2329
rect 5908 2320 5960 2372
rect 3792 2252 3844 2304
rect 7840 2252 7892 2304
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 9772 2295 9824 2304
rect 9772 2261 9781 2295
rect 9781 2261 9815 2295
rect 9815 2261 9824 2295
rect 9772 2252 9824 2261
rect 10876 2252 10928 2304
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 12348 2388 12400 2440
rect 13084 2431 13136 2440
rect 13084 2397 13093 2431
rect 13093 2397 13127 2431
rect 13127 2397 13136 2431
rect 13084 2388 13136 2397
rect 13176 2431 13228 2440
rect 13176 2397 13185 2431
rect 13185 2397 13219 2431
rect 13219 2397 13228 2431
rect 13176 2388 13228 2397
rect 12440 2320 12492 2372
rect 15200 2456 15252 2508
rect 15568 2456 15620 2508
rect 17040 2456 17092 2508
rect 17684 2499 17736 2508
rect 17684 2465 17693 2499
rect 17693 2465 17727 2499
rect 17727 2465 17736 2499
rect 17684 2456 17736 2465
rect 17960 2456 18012 2508
rect 19708 2635 19760 2644
rect 18788 2567 18840 2576
rect 18788 2533 18797 2567
rect 18797 2533 18831 2567
rect 18831 2533 18840 2567
rect 18788 2524 18840 2533
rect 19708 2601 19717 2635
rect 19717 2601 19751 2635
rect 19751 2601 19760 2635
rect 19708 2592 19760 2601
rect 20536 2592 20588 2644
rect 20628 2567 20680 2576
rect 20628 2533 20637 2567
rect 20637 2533 20671 2567
rect 20671 2533 20680 2567
rect 20628 2524 20680 2533
rect 19892 2456 19944 2508
rect 18604 2388 18656 2440
rect 18696 2388 18748 2440
rect 19984 2431 20036 2440
rect 14464 2320 14516 2372
rect 17960 2320 18012 2372
rect 18972 2320 19024 2372
rect 16304 2252 16356 2304
rect 17316 2252 17368 2304
rect 19984 2397 19993 2431
rect 19993 2397 20027 2431
rect 20027 2397 20036 2431
rect 19984 2388 20036 2397
rect 19984 2252 20036 2304
rect 20444 2252 20496 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 4160 2048 4212 2100
rect 4988 2048 5040 2100
rect 9956 2048 10008 2100
rect 16212 2048 16264 2100
rect 16580 2048 16632 2100
rect 18604 2048 18656 2100
rect 18788 2048 18840 2100
rect 19432 2048 19484 2100
rect 2780 1980 2832 2032
rect 7012 1980 7064 2032
rect 8208 1980 8260 2032
rect 10876 1980 10928 2032
rect 204 1912 256 1964
rect 8300 1912 8352 1964
rect 9036 1912 9088 1964
rect 9312 1912 9364 1964
rect 21456 1912 21508 1964
rect 6552 1844 6604 1896
rect 10324 1844 10376 1896
rect 11060 1844 11112 1896
rect 19892 1844 19944 1896
rect 4896 1776 4948 1828
rect 9772 1776 9824 1828
rect 10140 1776 10192 1828
rect 10968 1776 11020 1828
rect 11980 1776 12032 1828
rect 18880 1776 18932 1828
rect 20720 1776 20772 1828
rect 572 1708 624 1760
rect 7748 1708 7800 1760
rect 7840 1708 7892 1760
rect 13544 1708 13596 1760
rect 5724 1640 5776 1692
rect 1308 1572 1360 1624
rect 7564 1572 7616 1624
rect 8760 1615 8812 1624
rect 8760 1581 8769 1615
rect 8769 1581 8803 1615
rect 8803 1581 8812 1615
rect 17868 1640 17920 1692
rect 8760 1572 8812 1581
rect 13820 1572 13872 1624
rect 16212 1572 16264 1624
rect 17224 1572 17276 1624
rect 19616 1572 19668 1624
rect 3976 1504 4028 1556
rect 17592 1504 17644 1556
rect 7196 1436 7248 1488
rect 11704 1436 11756 1488
rect 5356 1368 5408 1420
rect 9680 1368 9732 1420
rect 14372 1368 14424 1420
rect 10784 1232 10836 1284
rect 15108 1232 15160 1284
rect 2044 1164 2096 1216
rect 7196 1164 7248 1216
rect 1676 1096 1728 1148
rect 7380 1096 7432 1148
<< metal2 >>
rect 202 22320 258 22800
rect 570 22320 626 22800
rect 938 22320 994 22800
rect 1306 22320 1362 22800
rect 1674 22320 1730 22800
rect 2042 22320 2098 22800
rect 2410 22320 2466 22800
rect 2778 22320 2834 22800
rect 3238 22320 3294 22800
rect 3514 22672 3570 22681
rect 3514 22607 3570 22616
rect 216 17814 244 22320
rect 584 18902 612 22320
rect 952 19242 980 22320
rect 940 19236 992 19242
rect 940 19178 992 19184
rect 1320 19174 1348 22320
rect 1688 20534 1716 22320
rect 1950 20632 2006 20641
rect 1950 20567 2006 20576
rect 1676 20528 1728 20534
rect 1676 20470 1728 20476
rect 1860 19848 1912 19854
rect 1860 19790 1912 19796
rect 1872 19417 1900 19790
rect 1858 19408 1914 19417
rect 1858 19343 1914 19352
rect 1964 19310 1992 20567
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1584 19236 1636 19242
rect 1584 19178 1636 19184
rect 1308 19168 1360 19174
rect 1308 19110 1360 19116
rect 1596 19009 1624 19178
rect 1582 19000 1638 19009
rect 1638 18958 1716 18986
rect 1582 18935 1638 18944
rect 572 18896 624 18902
rect 572 18838 624 18844
rect 1584 18624 1636 18630
rect 1584 18566 1636 18572
rect 1490 17912 1546 17921
rect 1490 17847 1546 17856
rect 204 17808 256 17814
rect 204 17750 256 17756
rect 1216 17128 1268 17134
rect 1216 17070 1268 17076
rect 1122 16280 1178 16289
rect 1122 16215 1178 16224
rect 1136 12442 1164 16215
rect 1228 12481 1256 17070
rect 1504 16250 1532 17847
rect 1596 17513 1624 18566
rect 1688 17882 1716 18958
rect 2056 18766 2084 22320
rect 2424 20074 2452 22320
rect 2792 21162 2820 22320
rect 2792 21134 3004 21162
rect 2870 21040 2926 21049
rect 2870 20975 2926 20984
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 2332 20046 2544 20074
rect 2332 18970 2360 20046
rect 2516 19990 2544 20046
rect 2504 19984 2556 19990
rect 2504 19926 2556 19932
rect 2608 19922 2636 20402
rect 2596 19916 2648 19922
rect 2596 19858 2648 19864
rect 2780 19848 2832 19854
rect 2778 19816 2780 19825
rect 2832 19816 2834 19825
rect 2778 19751 2834 19760
rect 2884 19310 2912 20975
rect 2412 19304 2464 19310
rect 2412 19246 2464 19252
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2320 18964 2372 18970
rect 2320 18906 2372 18912
rect 2424 18850 2452 19246
rect 2504 19236 2556 19242
rect 2504 19178 2556 19184
rect 2136 18828 2188 18834
rect 2136 18770 2188 18776
rect 2332 18822 2452 18850
rect 2044 18760 2096 18766
rect 1950 18728 2006 18737
rect 2044 18702 2096 18708
rect 1950 18663 2006 18672
rect 1964 18426 1992 18663
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1952 18216 2004 18222
rect 1952 18158 2004 18164
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 1858 17912 1914 17921
rect 1676 17876 1728 17882
rect 1858 17847 1914 17856
rect 1676 17818 1728 17824
rect 1872 17814 1900 17847
rect 1860 17808 1912 17814
rect 1860 17750 1912 17756
rect 1582 17504 1638 17513
rect 1582 17439 1638 17448
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 1492 16244 1544 16250
rect 1492 16186 1544 16192
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 1492 15496 1544 15502
rect 1492 15438 1544 15444
rect 1400 13728 1452 13734
rect 1400 13670 1452 13676
rect 1306 13288 1362 13297
rect 1306 13223 1362 13232
rect 1214 12472 1270 12481
rect 1124 12436 1176 12442
rect 1214 12407 1270 12416
rect 1124 12378 1176 12384
rect 1320 10033 1348 13223
rect 1306 10024 1362 10033
rect 1306 9959 1362 9968
rect 1412 8430 1440 13670
rect 1504 12306 1532 15438
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1596 14385 1624 15302
rect 1582 14376 1638 14385
rect 1582 14311 1638 14320
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1596 12986 1624 13330
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1504 8673 1532 12242
rect 1688 11801 1716 15982
rect 1780 14958 1808 17070
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1860 13728 1912 13734
rect 1860 13670 1912 13676
rect 1766 13560 1822 13569
rect 1766 13495 1822 13504
rect 1674 11792 1730 11801
rect 1674 11727 1730 11736
rect 1676 11620 1728 11626
rect 1676 11562 1728 11568
rect 1582 11248 1638 11257
rect 1582 11183 1638 11192
rect 1490 8664 1546 8673
rect 1490 8599 1546 8608
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1400 8288 1452 8294
rect 1400 8230 1452 8236
rect 1412 7002 1440 8230
rect 1400 6996 1452 7002
rect 1400 6938 1452 6944
rect 1596 6458 1624 11183
rect 1688 9042 1716 11562
rect 1780 10266 1808 13495
rect 1872 11778 1900 13670
rect 1964 13190 1992 18158
rect 2056 17134 2084 18158
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 2148 16046 2176 18770
rect 2332 18465 2360 18822
rect 2412 18760 2464 18766
rect 2516 18737 2544 19178
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2700 18902 2728 19110
rect 2688 18896 2740 18902
rect 2688 18838 2740 18844
rect 2688 18760 2740 18766
rect 2412 18702 2464 18708
rect 2502 18728 2558 18737
rect 2318 18456 2374 18465
rect 2424 18426 2452 18702
rect 2688 18702 2740 18708
rect 2502 18663 2558 18672
rect 2318 18391 2374 18400
rect 2412 18420 2464 18426
rect 2412 18362 2464 18368
rect 2410 17776 2466 17785
rect 2410 17711 2466 17720
rect 2596 17740 2648 17746
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2044 16040 2096 16046
rect 2044 15982 2096 15988
rect 2136 16040 2188 16046
rect 2136 15982 2188 15988
rect 2056 14226 2084 15982
rect 2240 15570 2268 17614
rect 2318 17232 2374 17241
rect 2318 17167 2374 17176
rect 2332 16726 2360 17167
rect 2424 16726 2452 17711
rect 2596 17682 2648 17688
rect 2504 17060 2556 17066
rect 2504 17002 2556 17008
rect 2516 16794 2544 17002
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2320 16720 2372 16726
rect 2320 16662 2372 16668
rect 2412 16720 2464 16726
rect 2412 16662 2464 16668
rect 2608 16250 2636 17682
rect 2700 17134 2728 18702
rect 2872 18624 2924 18630
rect 2872 18566 2924 18572
rect 2780 18080 2832 18086
rect 2780 18022 2832 18028
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2700 16590 2728 17070
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 2596 16244 2648 16250
rect 2596 16186 2648 16192
rect 2700 16114 2728 16526
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 2792 16046 2820 18022
rect 2884 17882 2912 18566
rect 2976 18306 3004 21134
rect 3252 20074 3280 22320
rect 3160 20046 3280 20074
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 3068 19145 3096 19246
rect 3054 19136 3110 19145
rect 3054 19071 3110 19080
rect 2976 18278 3096 18306
rect 3068 18222 3096 18278
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 2964 18148 3016 18154
rect 2964 18090 3016 18096
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 2976 17678 3004 18090
rect 3056 17740 3108 17746
rect 3056 17682 3108 17688
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 3068 17105 3096 17682
rect 3160 17354 3188 20046
rect 3240 19916 3292 19922
rect 3240 19858 3292 19864
rect 3252 18970 3280 19858
rect 3332 19440 3384 19446
rect 3332 19382 3384 19388
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 3344 17746 3372 19382
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3436 17882 3464 18702
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3332 17740 3384 17746
rect 3332 17682 3384 17688
rect 3240 17672 3292 17678
rect 3292 17620 3464 17626
rect 3240 17614 3464 17620
rect 3252 17598 3464 17614
rect 3160 17326 3280 17354
rect 3436 17338 3464 17598
rect 3148 17128 3200 17134
rect 3054 17096 3110 17105
rect 3148 17070 3200 17076
rect 3054 17031 3110 17040
rect 2780 16040 2832 16046
rect 2318 16008 2374 16017
rect 2780 15982 2832 15988
rect 2318 15943 2374 15952
rect 2332 15706 2360 15943
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 2228 15564 2280 15570
rect 2228 15506 2280 15512
rect 2424 15450 2452 15846
rect 2594 15736 2650 15745
rect 2594 15671 2650 15680
rect 2608 15570 2636 15671
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2332 15422 2452 15450
rect 2056 14198 2176 14226
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1964 12442 1992 12582
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1872 11750 2084 11778
rect 1860 11620 1912 11626
rect 1860 11562 1912 11568
rect 1872 11218 1900 11562
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1768 9512 1820 9518
rect 1872 9500 1900 10202
rect 1820 9472 1900 9500
rect 1768 9454 1820 9460
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1780 8922 1808 9454
rect 1964 9178 1992 11494
rect 2056 10266 2084 11750
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2042 10160 2098 10169
rect 2042 10095 2098 10104
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1688 8894 1808 8922
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1582 6352 1638 6361
rect 1582 6287 1638 6296
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1412 5846 1440 6190
rect 1400 5840 1452 5846
rect 1400 5782 1452 5788
rect 1596 5370 1624 6287
rect 1688 5545 1716 8894
rect 2056 8616 2084 10095
rect 1964 8588 2084 8616
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1780 7410 1808 7686
rect 1768 7404 1820 7410
rect 1820 7364 1900 7392
rect 1768 7346 1820 7352
rect 1766 7168 1822 7177
rect 1766 7103 1822 7112
rect 1780 6866 1808 7103
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1766 6760 1822 6769
rect 1766 6695 1768 6704
rect 1820 6695 1822 6704
rect 1768 6666 1820 6672
rect 1768 6384 1820 6390
rect 1768 6326 1820 6332
rect 1674 5536 1730 5545
rect 1674 5471 1730 5480
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1674 4992 1730 5001
rect 1674 4927 1730 4936
rect 1122 3904 1178 3913
rect 1122 3839 1178 3848
rect 938 3632 994 3641
rect 938 3567 994 3576
rect 204 1964 256 1970
rect 204 1906 256 1912
rect 216 480 244 1906
rect 572 1760 624 1766
rect 572 1702 624 1708
rect 584 480 612 1702
rect 952 480 980 3567
rect 1136 2961 1164 3839
rect 1688 3670 1716 4927
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1122 2952 1178 2961
rect 1122 2887 1178 2896
rect 1780 2825 1808 6326
rect 1872 5710 1900 7364
rect 1964 6202 1992 8588
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2056 7274 2084 8434
rect 2044 7268 2096 7274
rect 2044 7210 2096 7216
rect 2148 6458 2176 14198
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2240 6474 2268 10406
rect 2332 10130 2360 15422
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2424 15162 2452 15302
rect 2412 15156 2464 15162
rect 2412 15098 2464 15104
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2424 13530 2452 14894
rect 2608 13938 2636 15506
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2792 14890 2820 15438
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2792 14414 2820 14826
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2594 13832 2650 13841
rect 2792 13802 2820 14214
rect 2884 14006 2912 14418
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 2976 13870 3004 15302
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2594 13767 2650 13776
rect 2780 13796 2832 13802
rect 2608 13734 2636 13767
rect 2780 13738 2832 13744
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2424 13394 2452 13466
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2424 12782 2452 13330
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2424 11626 2452 12718
rect 2608 12238 2636 13330
rect 2870 13152 2926 13161
rect 2870 13087 2926 13096
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2412 11620 2464 11626
rect 2412 11562 2464 11568
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2596 10532 2648 10538
rect 2596 10474 2648 10480
rect 2320 10124 2372 10130
rect 2320 10066 2372 10072
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2332 9110 2360 9862
rect 2516 9722 2544 10066
rect 2608 10062 2636 10474
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2608 9586 2636 9998
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2412 9444 2464 9450
rect 2412 9386 2464 9392
rect 2424 9178 2452 9386
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2320 9104 2372 9110
rect 2320 9046 2372 9052
rect 2516 8634 2544 9318
rect 2700 8974 2728 11154
rect 2884 10266 2912 13087
rect 3160 12424 3188 17070
rect 2976 12396 3188 12424
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2780 10192 2832 10198
rect 2976 10146 3004 12396
rect 3146 12336 3202 12345
rect 3146 12271 3202 12280
rect 3054 11928 3110 11937
rect 3054 11863 3110 11872
rect 2780 10134 2832 10140
rect 2792 9178 2820 10134
rect 2884 10118 3004 10146
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2778 8528 2834 8537
rect 2778 8463 2834 8472
rect 2596 7948 2648 7954
rect 2596 7890 2648 7896
rect 2608 7834 2636 7890
rect 2608 7806 2728 7834
rect 2700 7546 2728 7806
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2700 6798 2728 7482
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 2136 6452 2188 6458
rect 2240 6446 2360 6474
rect 2136 6394 2188 6400
rect 2332 6390 2360 6446
rect 2320 6384 2372 6390
rect 2320 6326 2372 6332
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 1964 6174 2084 6202
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1964 5778 1992 6054
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 1872 5234 1900 5646
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1872 4758 1900 5170
rect 1860 4752 1912 4758
rect 1860 4694 1912 4700
rect 1872 3602 1900 4694
rect 2056 3738 2084 6174
rect 2240 5098 2268 6258
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2228 5092 2280 5098
rect 2228 5034 2280 5040
rect 2240 4826 2268 5034
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2228 4684 2280 4690
rect 2228 4626 2280 4632
rect 2240 4146 2268 4626
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2240 3738 2268 4082
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1872 3194 1900 3538
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 2240 3058 2268 3674
rect 2332 3126 2360 6054
rect 2424 3942 2452 6054
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2792 3777 2820 8463
rect 2884 4690 2912 10118
rect 3068 8906 3096 11863
rect 3160 9586 3188 12271
rect 3252 11898 3280 17326
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 3422 16688 3478 16697
rect 3332 16652 3384 16658
rect 3422 16623 3424 16632
rect 3332 16594 3384 16600
rect 3476 16623 3478 16632
rect 3424 16594 3476 16600
rect 3344 16561 3372 16594
rect 3330 16552 3386 16561
rect 3330 16487 3386 16496
rect 3528 15722 3556 22607
rect 3606 22320 3662 22800
rect 3974 22320 4030 22800
rect 4342 22320 4398 22800
rect 4710 22320 4766 22800
rect 5078 22320 5134 22800
rect 5446 22320 5502 22800
rect 5906 22320 5962 22800
rect 6274 22320 6330 22800
rect 6642 22320 6698 22800
rect 7010 22320 7066 22800
rect 7378 22320 7434 22800
rect 7746 22320 7802 22800
rect 8114 22320 8170 22800
rect 8482 22320 8538 22800
rect 8942 22320 8998 22800
rect 9310 22320 9366 22800
rect 9678 22320 9734 22800
rect 10046 22320 10102 22800
rect 10414 22320 10470 22800
rect 10782 22320 10838 22800
rect 11150 22320 11206 22800
rect 11610 22320 11666 22800
rect 11978 22320 12034 22800
rect 12346 22320 12402 22800
rect 12714 22320 12770 22800
rect 13082 22320 13138 22800
rect 13450 22320 13506 22800
rect 13818 22320 13874 22800
rect 14186 22320 14242 22800
rect 14646 22320 14702 22800
rect 15014 22320 15070 22800
rect 15382 22320 15438 22800
rect 15750 22320 15806 22800
rect 16118 22320 16174 22800
rect 16486 22320 16542 22800
rect 16854 22320 16910 22800
rect 17314 22320 17370 22800
rect 17682 22320 17738 22800
rect 18050 22320 18106 22800
rect 18418 22320 18474 22800
rect 18786 22320 18842 22800
rect 19154 22320 19210 22800
rect 19522 22320 19578 22800
rect 19890 22320 19946 22800
rect 20350 22320 20406 22800
rect 20626 22672 20682 22681
rect 20626 22607 20682 22616
rect 3620 18408 3648 22320
rect 3882 22264 3938 22273
rect 3882 22199 3938 22208
rect 3698 21856 3754 21865
rect 3698 21791 3754 21800
rect 3712 21146 3740 21791
rect 3700 21140 3752 21146
rect 3700 21082 3752 21088
rect 3792 20324 3844 20330
rect 3792 20266 3844 20272
rect 3804 20058 3832 20266
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 3792 19440 3844 19446
rect 3792 19382 3844 19388
rect 3620 18380 3740 18408
rect 3606 18320 3662 18329
rect 3606 18255 3662 18264
rect 3620 17610 3648 18255
rect 3712 18057 3740 18380
rect 3804 18222 3832 19382
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 3698 18048 3754 18057
rect 3698 17983 3754 17992
rect 3790 17640 3846 17649
rect 3608 17604 3660 17610
rect 3790 17575 3846 17584
rect 3608 17546 3660 17552
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 3620 17105 3648 17274
rect 3804 17202 3832 17575
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3606 17096 3662 17105
rect 3606 17031 3662 17040
rect 3698 16824 3754 16833
rect 3698 16759 3754 16768
rect 3712 16726 3740 16759
rect 3700 16720 3752 16726
rect 3700 16662 3752 16668
rect 3528 15694 3648 15722
rect 3516 14884 3568 14890
rect 3516 14826 3568 14832
rect 3422 14784 3478 14793
rect 3422 14719 3478 14728
rect 3332 14340 3384 14346
rect 3332 14282 3384 14288
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3344 11778 3372 14282
rect 3436 12646 3464 14719
rect 3528 14328 3556 14826
rect 3620 14550 3648 15694
rect 3896 15586 3924 22199
rect 3988 17134 4016 22320
rect 4356 22250 4384 22320
rect 4172 22222 4384 22250
rect 4066 21448 4122 21457
rect 4066 21383 4068 21392
rect 4120 21383 4122 21392
rect 4068 21354 4120 21360
rect 4068 20256 4120 20262
rect 4066 20224 4068 20233
rect 4120 20224 4122 20233
rect 4066 20159 4122 20168
rect 4172 20074 4200 22222
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 4080 20046 4200 20074
rect 4080 19378 4108 20046
rect 4264 19854 4292 20470
rect 4724 20398 4752 22320
rect 4712 20392 4764 20398
rect 4712 20334 4764 20340
rect 4988 19916 5040 19922
rect 4988 19858 5040 19864
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4160 19780 4212 19786
rect 4160 19722 4212 19728
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 4172 19174 4200 19722
rect 4264 19310 4292 19790
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4344 19372 4396 19378
rect 4396 19332 4476 19360
rect 4344 19314 4396 19320
rect 4252 19304 4304 19310
rect 4252 19246 4304 19252
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 4448 18873 4476 19332
rect 4724 18952 4752 19790
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4632 18924 4752 18952
rect 4434 18864 4490 18873
rect 4434 18799 4490 18808
rect 4632 18714 4660 18924
rect 4816 18902 4844 19246
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4908 18902 4936 19110
rect 4804 18896 4856 18902
rect 4804 18838 4856 18844
rect 4896 18896 4948 18902
rect 4896 18838 4948 18844
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4264 18686 4660 18714
rect 4264 17270 4292 18686
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4724 18154 4752 18770
rect 4816 18714 4844 18838
rect 4816 18686 4936 18714
rect 4802 18592 4858 18601
rect 4802 18527 4858 18536
rect 4816 18426 4844 18527
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4356 17882 4384 18022
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4724 17678 4752 18090
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4252 17264 4304 17270
rect 4252 17206 4304 17212
rect 4712 17196 4764 17202
rect 4816 17184 4844 18226
rect 4908 18086 4936 18686
rect 5000 18193 5028 19858
rect 5092 19417 5120 22320
rect 5172 20392 5224 20398
rect 5172 20334 5224 20340
rect 5078 19408 5134 19417
rect 5078 19343 5134 19352
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 4986 18184 5042 18193
rect 4986 18119 5042 18128
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4764 17156 4844 17184
rect 4712 17138 4764 17144
rect 3976 17128 4028 17134
rect 4724 17105 4752 17138
rect 3976 17070 4028 17076
rect 4710 17096 4766 17105
rect 4710 17031 4766 17040
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 3976 16448 4028 16454
rect 3976 16390 4028 16396
rect 3988 16114 4016 16390
rect 4264 16114 4292 16730
rect 4540 16522 4568 16730
rect 4528 16516 4580 16522
rect 4528 16458 4580 16464
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4620 16176 4672 16182
rect 4724 16164 4752 17031
rect 4908 16658 4936 18022
rect 5092 17882 5120 18906
rect 5080 17876 5132 17882
rect 5080 17818 5132 17824
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 5000 17134 5028 17478
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 5092 16794 5120 16934
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 4988 16720 5040 16726
rect 4988 16662 5040 16668
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4672 16136 4752 16164
rect 4620 16118 4672 16124
rect 4816 16114 4844 16594
rect 4896 16448 4948 16454
rect 4896 16390 4948 16396
rect 3976 16108 4028 16114
rect 3976 16050 4028 16056
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 4620 15972 4672 15978
rect 4620 15914 4672 15920
rect 4066 15872 4122 15881
rect 4066 15807 4122 15816
rect 4080 15706 4108 15807
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4632 15638 4660 15914
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4620 15632 4672 15638
rect 3896 15558 4108 15586
rect 4620 15574 4672 15580
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3882 15464 3938 15473
rect 3608 14544 3660 14550
rect 3608 14486 3660 14492
rect 3608 14340 3660 14346
rect 3528 14300 3608 14328
rect 3528 13938 3556 14300
rect 3608 14282 3660 14288
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3516 13796 3568 13802
rect 3516 13738 3568 13744
rect 3700 13796 3752 13802
rect 3700 13738 3752 13744
rect 3528 13530 3556 13738
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3712 13190 3740 13738
rect 3700 13184 3752 13190
rect 3700 13126 3752 13132
rect 3712 12782 3740 13126
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3252 11750 3372 11778
rect 3252 11234 3280 11750
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3344 11354 3372 11630
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3252 11206 3372 11234
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3252 10810 3280 11018
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3238 10024 3294 10033
rect 3238 9959 3294 9968
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 3252 9466 3280 9959
rect 3344 9586 3372 11206
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3436 9466 3464 12174
rect 3528 11354 3556 12242
rect 3620 12238 3648 12650
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3514 11248 3570 11257
rect 3514 11183 3570 11192
rect 3528 10606 3556 11183
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3528 9518 3556 9862
rect 3620 9738 3648 11834
rect 3712 10810 3740 12582
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3620 9710 3740 9738
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3160 9438 3280 9466
rect 3344 9438 3464 9466
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 2964 6928 3016 6934
rect 2964 6870 3016 6876
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2778 3768 2834 3777
rect 2778 3703 2834 3712
rect 2320 3120 2372 3126
rect 2320 3062 2372 3068
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2044 2848 2096 2854
rect 1766 2816 1822 2825
rect 2044 2790 2096 2796
rect 2686 2816 2742 2825
rect 1766 2751 1822 2760
rect 2056 2650 2084 2790
rect 2686 2751 2742 2760
rect 2410 2680 2466 2689
rect 2044 2644 2096 2650
rect 2700 2650 2728 2751
rect 2410 2615 2466 2624
rect 2688 2644 2740 2650
rect 2044 2586 2096 2592
rect 1950 2544 2006 2553
rect 1950 2479 1952 2488
rect 2004 2479 2006 2488
rect 1952 2450 2004 2456
rect 1308 1624 1360 1630
rect 1308 1566 1360 1572
rect 1320 480 1348 1566
rect 2044 1216 2096 1222
rect 2044 1158 2096 1164
rect 1676 1148 1728 1154
rect 1676 1090 1728 1096
rect 1688 480 1716 1090
rect 2056 480 2084 1158
rect 2424 480 2452 2615
rect 2688 2586 2740 2592
rect 2596 2576 2648 2582
rect 2596 2518 2648 2524
rect 2608 2446 2636 2518
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2976 2145 3004 6870
rect 3068 2854 3096 8366
rect 3160 5250 3188 9438
rect 3240 8900 3292 8906
rect 3240 8842 3292 8848
rect 3252 8498 3280 8842
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3344 8430 3372 9438
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 9178 3464 9318
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3436 8566 3464 8910
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3528 6848 3556 9454
rect 3620 9382 3648 9522
rect 3608 9376 3660 9382
rect 3712 9353 3740 9710
rect 3608 9318 3660 9324
rect 3698 9344 3754 9353
rect 3620 6934 3648 9318
rect 3698 9279 3754 9288
rect 3804 9110 3832 15438
rect 3882 15399 3938 15408
rect 3896 12442 3924 15399
rect 3974 15192 4030 15201
rect 3974 15127 4030 15136
rect 3988 13734 4016 15127
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 4080 13546 4108 15558
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4528 14544 4580 14550
rect 4528 14486 4580 14492
rect 4540 14260 4568 14486
rect 4632 14414 4660 14758
rect 4724 14482 4752 15846
rect 4908 15609 4936 16390
rect 4894 15600 4950 15609
rect 4804 15564 4856 15570
rect 4894 15535 4950 15544
rect 4804 15506 4856 15512
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4540 14232 4752 14260
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4250 13968 4306 13977
rect 4250 13903 4306 13912
rect 3988 13518 4108 13546
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3882 11656 3938 11665
rect 3882 11591 3938 11600
rect 3896 11286 3924 11591
rect 3884 11280 3936 11286
rect 3884 11222 3936 11228
rect 3884 9988 3936 9994
rect 3884 9930 3936 9936
rect 3896 9722 3924 9930
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3792 9104 3844 9110
rect 3698 9072 3754 9081
rect 3792 9046 3844 9052
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3698 9007 3754 9016
rect 3712 8430 3740 9007
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3608 6928 3660 6934
rect 3608 6870 3660 6876
rect 3344 6820 3556 6848
rect 3700 6860 3752 6866
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3252 5370 3280 6054
rect 3344 5692 3372 6820
rect 3700 6802 3752 6808
rect 3422 6760 3478 6769
rect 3422 6695 3478 6704
rect 3606 6760 3662 6769
rect 3606 6695 3662 6704
rect 3436 5817 3464 6695
rect 3620 6662 3648 6695
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3422 5808 3478 5817
rect 3422 5743 3478 5752
rect 3344 5664 3464 5692
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3332 5296 3384 5302
rect 3160 5222 3280 5250
rect 3332 5238 3384 5244
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 3160 4146 3188 4490
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3252 3233 3280 5222
rect 3344 4826 3372 5238
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3344 3602 3372 4082
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 3238 3224 3294 3233
rect 3238 3159 3294 3168
rect 3344 3058 3372 3538
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 2962 2136 3018 2145
rect 2962 2071 3018 2080
rect 2780 2032 2832 2038
rect 2780 1974 2832 1980
rect 2792 480 2820 1974
rect 3068 1737 3096 2790
rect 3344 2650 3372 2994
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 3054 1728 3110 1737
rect 3054 1663 3110 1672
rect 3160 480 3188 2518
rect 3436 2514 3464 5664
rect 3528 5574 3556 6258
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3528 480 3556 5510
rect 3620 5030 3648 6326
rect 3712 5914 3740 6802
rect 3804 6322 3832 8502
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3620 4706 3648 4966
rect 3712 4826 3740 5102
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3620 4678 3740 4706
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3620 4282 3648 4558
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3712 4049 3740 4678
rect 3698 4040 3754 4049
rect 3698 3975 3754 3984
rect 3700 3936 3752 3942
rect 3804 3913 3832 6258
rect 3896 6236 3924 9046
rect 3988 8634 4016 13518
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 4080 12918 4108 13262
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4172 12986 4200 13126
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4068 12912 4120 12918
rect 4264 12866 4292 13903
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4068 12854 4120 12860
rect 4172 12838 4292 12866
rect 4066 12744 4122 12753
rect 4066 12679 4122 12688
rect 4080 11642 4108 12679
rect 4172 11898 4200 12838
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4264 12238 4292 12582
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4356 12084 4384 12174
rect 4724 12102 4752 14232
rect 4816 12628 4844 15506
rect 4896 15428 4948 15434
rect 4896 15370 4948 15376
rect 4908 14006 4936 15370
rect 5000 14414 5028 16662
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 5092 16522 5120 16594
rect 5080 16516 5132 16522
rect 5080 16458 5132 16464
rect 5092 14958 5120 16458
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5078 14784 5134 14793
rect 5078 14719 5134 14728
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 4896 14000 4948 14006
rect 4896 13942 4948 13948
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 5000 13190 5028 13806
rect 5092 13546 5120 14719
rect 5184 13682 5212 20334
rect 5460 20074 5488 22320
rect 5460 20046 5672 20074
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5276 17921 5304 19790
rect 5356 19780 5408 19786
rect 5356 19722 5408 19728
rect 5368 19310 5396 19722
rect 5460 19394 5488 19858
rect 5460 19366 5580 19394
rect 5356 19304 5408 19310
rect 5356 19246 5408 19252
rect 5552 19242 5580 19366
rect 5644 19310 5672 20046
rect 5816 19508 5868 19514
rect 5816 19450 5868 19456
rect 5632 19304 5684 19310
rect 5632 19246 5684 19252
rect 5448 19236 5500 19242
rect 5448 19178 5500 19184
rect 5540 19236 5592 19242
rect 5540 19178 5592 19184
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5368 18154 5396 18566
rect 5347 18148 5399 18154
rect 5347 18090 5399 18096
rect 5460 18086 5488 19178
rect 5828 19174 5856 19450
rect 5816 19168 5868 19174
rect 5630 19136 5686 19145
rect 5816 19110 5868 19116
rect 5630 19071 5686 19080
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5262 17912 5318 17921
rect 5262 17847 5318 17856
rect 5264 17808 5316 17814
rect 5264 17750 5316 17756
rect 5276 15366 5304 17750
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5264 15360 5316 15366
rect 5368 15337 5396 16730
rect 5460 16250 5488 17682
rect 5540 17672 5592 17678
rect 5538 17640 5540 17649
rect 5592 17640 5594 17649
rect 5538 17575 5594 17584
rect 5644 16998 5672 19071
rect 5828 18766 5856 19110
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5736 18426 5764 18566
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5828 18306 5856 18702
rect 5920 18630 5948 22320
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 5908 18624 5960 18630
rect 5908 18566 5960 18572
rect 5736 18278 5856 18306
rect 5736 17202 5764 18278
rect 5816 18080 5868 18086
rect 5816 18022 5868 18028
rect 5828 17746 5856 18022
rect 6104 17882 6132 19858
rect 6184 19712 6236 19718
rect 6184 19654 6236 19660
rect 6196 18970 6224 19654
rect 6184 18964 6236 18970
rect 6184 18906 6236 18912
rect 6288 18290 6316 22320
rect 6656 20210 6684 22320
rect 6656 20182 6868 20210
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 6552 19304 6604 19310
rect 6552 19246 6604 19252
rect 6368 19168 6420 19174
rect 6368 19110 6420 19116
rect 6380 19009 6408 19110
rect 6366 19000 6422 19009
rect 6366 18935 6422 18944
rect 6380 18834 6408 18935
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6276 18284 6328 18290
rect 6276 18226 6328 18232
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6366 18048 6422 18057
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 6092 17876 6144 17882
rect 6092 17818 6144 17824
rect 5816 17740 5868 17746
rect 5816 17682 5868 17688
rect 6012 17610 6040 17818
rect 6288 17678 6316 18022
rect 6366 17983 6422 17992
rect 6276 17672 6328 17678
rect 6380 17649 6408 17983
rect 6276 17614 6328 17620
rect 6366 17640 6422 17649
rect 6000 17604 6052 17610
rect 6366 17575 6422 17584
rect 6000 17546 6052 17552
rect 5816 17332 5868 17338
rect 5816 17274 5868 17280
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 5552 15978 5580 16390
rect 5644 16232 5672 16934
rect 5736 16726 5764 17138
rect 5828 16998 5856 17274
rect 5908 17264 5960 17270
rect 5908 17206 5960 17212
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 5724 16720 5776 16726
rect 5724 16662 5776 16668
rect 5644 16204 5764 16232
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5264 15302 5316 15308
rect 5354 15328 5410 15337
rect 5354 15263 5410 15272
rect 5262 15192 5318 15201
rect 5262 15127 5264 15136
rect 5316 15127 5318 15136
rect 5264 15098 5316 15104
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 5276 13870 5304 14826
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 5368 14385 5396 14418
rect 5354 14376 5410 14385
rect 5354 14311 5410 14320
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5368 13870 5396 14214
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5184 13654 5396 13682
rect 5092 13518 5212 13546
rect 5080 13456 5132 13462
rect 5080 13398 5132 13404
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4816 12600 5028 12628
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4264 12056 4384 12084
rect 4712 12096 4764 12102
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4080 11614 4200 11642
rect 4264 11626 4292 12056
rect 4712 12038 4764 12044
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4816 11830 4844 12242
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4896 11688 4948 11694
rect 4894 11656 4896 11665
rect 4948 11656 4950 11665
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4080 11354 4108 11494
rect 4172 11354 4200 11614
rect 4252 11620 4304 11626
rect 4894 11591 4950 11600
rect 4252 11562 4304 11568
rect 4802 11520 4858 11529
rect 4802 11455 4858 11464
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4712 11280 4764 11286
rect 4712 11222 4764 11228
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4172 10810 4200 11154
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 4080 10130 4108 10678
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4080 8430 4108 10066
rect 4172 9586 4200 10066
rect 4264 9654 4292 11086
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4724 10810 4752 11222
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4540 10266 4568 10610
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4724 10130 4752 10406
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4252 9648 4304 9654
rect 4816 9602 4844 11455
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4908 10305 4936 10542
rect 4894 10296 4950 10305
rect 4894 10231 4950 10240
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 4252 9590 4304 9596
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4693 9574 4844 9602
rect 4172 8974 4200 9522
rect 4693 9466 4721 9574
rect 4802 9480 4858 9489
rect 4693 9438 4752 9466
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4540 9178 4568 9318
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4632 8974 4660 9318
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4620 8968 4672 8974
rect 4724 8945 4752 9438
rect 4802 9415 4858 9424
rect 4620 8910 4672 8916
rect 4710 8936 4766 8945
rect 4710 8871 4766 8880
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4250 8664 4306 8673
rect 4388 8656 4684 8676
rect 4306 8608 4476 8616
rect 4250 8599 4476 8608
rect 4264 8588 4476 8599
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3988 8090 4016 8230
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3988 7721 4016 7822
rect 4080 7750 4108 8366
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4068 7744 4120 7750
rect 3974 7712 4030 7721
rect 4068 7686 4120 7692
rect 3974 7647 4030 7656
rect 4080 7546 4108 7686
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 3976 6656 4028 6662
rect 3974 6624 3976 6633
rect 4028 6624 4030 6633
rect 3974 6559 4030 6568
rect 4080 6390 4108 7210
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 3896 6208 4016 6236
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 3896 5574 3924 5714
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3896 5234 3924 5510
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3988 5114 4016 6208
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4080 5166 4108 6054
rect 3896 5086 4016 5114
rect 4068 5160 4120 5166
rect 4172 5148 4200 8298
rect 4252 7948 4304 7954
rect 4252 7890 4304 7896
rect 4264 6798 4292 7890
rect 4356 7818 4384 8298
rect 4448 7857 4476 8588
rect 4434 7848 4490 7857
rect 4344 7812 4396 7818
rect 4434 7783 4490 7792
rect 4344 7754 4396 7760
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4724 7449 4752 8871
rect 4816 7936 4844 9415
rect 4908 9382 4936 10066
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4908 8430 4936 8978
rect 5000 8838 5028 12600
rect 5092 11218 5120 13398
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 5092 9625 5120 11018
rect 5078 9616 5134 9625
rect 5078 9551 5134 9560
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 4986 8664 5042 8673
rect 4986 8599 5042 8608
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4816 7908 4936 7936
rect 4804 7812 4856 7818
rect 4804 7754 4856 7760
rect 4710 7440 4766 7449
rect 4710 7375 4766 7384
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4250 6488 4306 6497
rect 4388 6480 4684 6500
rect 4250 6423 4252 6432
rect 4304 6423 4306 6432
rect 4252 6394 4304 6400
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4724 5953 4752 6258
rect 4710 5944 4766 5953
rect 4710 5879 4766 5888
rect 4724 5846 4752 5879
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4724 5234 4752 5782
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4252 5160 4304 5166
rect 4172 5120 4252 5148
rect 4068 5102 4120 5108
rect 4252 5102 4304 5108
rect 4344 5092 4396 5098
rect 3896 3942 3924 5086
rect 4344 5034 4396 5040
rect 4252 4684 4304 4690
rect 4356 4672 4384 5034
rect 4816 5001 4844 7754
rect 4908 5545 4936 7908
rect 5000 5681 5028 8599
rect 5092 8430 5120 9386
rect 5184 9353 5212 13518
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5276 9382 5304 12582
rect 5368 11937 5396 13654
rect 5460 13530 5488 15506
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5552 14618 5580 15302
rect 5644 15162 5672 15846
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 14074 5580 14214
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5736 13818 5764 16204
rect 5552 13790 5764 13818
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5460 12986 5488 13330
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5354 11928 5410 11937
rect 5354 11863 5410 11872
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5368 11082 5396 11698
rect 5552 11150 5580 13790
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5644 11898 5672 13262
rect 5736 12850 5764 13262
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5736 12442 5764 12786
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5736 11218 5764 11562
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5356 11076 5408 11082
rect 5356 11018 5408 11024
rect 5538 10976 5594 10985
rect 5538 10911 5594 10920
rect 5354 10704 5410 10713
rect 5354 10639 5410 10648
rect 5448 10668 5500 10674
rect 5368 9382 5396 10639
rect 5448 10610 5500 10616
rect 5460 9586 5488 10610
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5264 9376 5316 9382
rect 5170 9344 5226 9353
rect 5264 9318 5316 9324
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5170 9279 5226 9288
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 5184 8634 5212 9114
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5170 7712 5226 7721
rect 5170 7647 5226 7656
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5092 7206 5120 7346
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 5092 6798 5120 7142
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 5078 6216 5134 6225
rect 5078 6151 5134 6160
rect 4986 5672 5042 5681
rect 4986 5607 5042 5616
rect 5092 5574 5120 6151
rect 5080 5568 5132 5574
rect 4894 5536 4950 5545
rect 5080 5510 5132 5516
rect 4894 5471 4950 5480
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4802 4992 4858 5001
rect 4802 4927 4858 4936
rect 4908 4740 4936 5306
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4986 4992 5042 5001
rect 4986 4927 5042 4936
rect 5000 4826 5028 4927
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4816 4712 4936 4740
rect 4304 4644 4384 4672
rect 4712 4684 4764 4690
rect 4252 4626 4304 4632
rect 4712 4626 4764 4632
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3884 3936 3936 3942
rect 3700 3878 3752 3884
rect 3790 3904 3846 3913
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3620 921 3648 3674
rect 3712 3126 3740 3878
rect 3884 3878 3936 3884
rect 3790 3839 3846 3848
rect 3896 3738 3924 3878
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3882 3224 3938 3233
rect 3882 3159 3938 3168
rect 3700 3120 3752 3126
rect 3700 3062 3752 3068
rect 3790 3088 3846 3097
rect 3790 3023 3846 3032
rect 3804 2990 3832 3023
rect 3792 2984 3844 2990
rect 3698 2952 3754 2961
rect 3792 2926 3844 2932
rect 3698 2887 3754 2896
rect 3712 2854 3740 2887
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3700 2440 3752 2446
rect 3700 2382 3752 2388
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3712 1873 3740 2382
rect 3804 2310 3832 2382
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 3698 1864 3754 1873
rect 3698 1799 3754 1808
rect 3606 912 3662 921
rect 3606 847 3662 856
rect 3896 480 3924 3159
rect 3988 1562 4016 4422
rect 4160 3936 4212 3942
rect 4080 3896 4160 3924
rect 3976 1556 4028 1562
rect 3976 1498 4028 1504
rect 4080 1442 4108 3896
rect 4160 3878 4212 3884
rect 4264 3738 4292 4626
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4342 4176 4398 4185
rect 4342 4111 4398 4120
rect 4356 4078 4384 4111
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4724 3754 4752 4626
rect 4816 3942 4844 4712
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4252 3732 4304 3738
rect 4724 3726 4844 3754
rect 4252 3674 4304 3680
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4172 3505 4200 3538
rect 4158 3496 4214 3505
rect 4342 3496 4398 3505
rect 4158 3431 4160 3440
rect 4212 3431 4214 3440
rect 4264 3454 4342 3482
rect 4160 3402 4212 3408
rect 4264 3369 4292 3454
rect 4342 3431 4398 3440
rect 4250 3360 4306 3369
rect 4250 3295 4306 3304
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4436 2984 4488 2990
rect 4436 2926 4488 2932
rect 4250 2816 4306 2825
rect 4250 2751 4306 2760
rect 4158 2544 4214 2553
rect 4158 2479 4214 2488
rect 4172 2378 4200 2479
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 4160 2100 4212 2106
rect 4160 2042 4212 2048
rect 3988 1414 4108 1442
rect 202 0 258 480
rect 570 0 626 480
rect 938 0 994 480
rect 1306 0 1362 480
rect 1674 0 1730 480
rect 2042 0 2098 480
rect 2410 0 2466 480
rect 2778 0 2834 480
rect 3146 0 3202 480
rect 3514 0 3570 480
rect 3882 0 3938 480
rect 3988 241 4016 1414
rect 4172 1329 4200 2042
rect 4158 1320 4214 1329
rect 4158 1255 4214 1264
rect 4264 480 4292 2751
rect 4448 2514 4476 2926
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 4342 2408 4398 2417
rect 4342 2343 4344 2352
rect 4396 2343 4398 2352
rect 4344 2314 4396 2320
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4816 2088 4844 3726
rect 4632 2060 4844 2088
rect 4632 480 4660 2060
rect 4908 1834 4936 3946
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 5000 3738 5028 3878
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 5092 3618 5120 5102
rect 5184 4826 5212 7647
rect 5276 5370 5304 9318
rect 5368 8945 5396 9318
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5354 8936 5410 8945
rect 5354 8871 5410 8880
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5262 5264 5318 5273
rect 5262 5199 5318 5208
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5184 4146 5212 4558
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5000 3590 5120 3618
rect 5000 2514 5028 3590
rect 5184 3534 5212 4082
rect 5276 4010 5304 5199
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5262 3768 5318 3777
rect 5262 3703 5318 3712
rect 5172 3528 5224 3534
rect 5078 3496 5134 3505
rect 5172 3470 5224 3476
rect 5078 3431 5134 3440
rect 4988 2508 5040 2514
rect 4988 2450 5040 2456
rect 5000 2106 5028 2450
rect 4988 2100 5040 2106
rect 4988 2042 5040 2048
rect 4896 1828 4948 1834
rect 4896 1770 4948 1776
rect 5092 1442 5120 3431
rect 5184 2922 5212 3470
rect 5276 3398 5304 3703
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5368 3210 5396 8774
rect 5460 8566 5488 9046
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5460 7546 5488 7890
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5552 6882 5580 10911
rect 5630 10704 5686 10713
rect 5630 10639 5686 10648
rect 5644 10606 5672 10639
rect 5632 10600 5684 10606
rect 5684 10560 5764 10588
rect 5632 10542 5684 10548
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5644 8294 5672 10202
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5736 7562 5764 10560
rect 5460 6854 5580 6882
rect 5644 7534 5764 7562
rect 5460 6633 5488 6854
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5446 6624 5502 6633
rect 5446 6559 5502 6568
rect 5460 5658 5488 6559
rect 5552 5846 5580 6734
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5460 5642 5580 5658
rect 5460 5636 5592 5642
rect 5460 5630 5540 5636
rect 5540 5578 5592 5584
rect 5446 5536 5502 5545
rect 5446 5471 5502 5480
rect 5460 4690 5488 5471
rect 5538 5400 5594 5409
rect 5538 5335 5594 5344
rect 5552 5098 5580 5335
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5644 4554 5672 7534
rect 5828 6984 5856 16934
rect 5920 16658 5948 17206
rect 6012 16658 6040 17546
rect 6380 16794 6408 17575
rect 6564 17338 6592 19246
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6368 16788 6420 16794
rect 6368 16730 6420 16736
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 5920 15745 5948 16594
rect 6184 16176 6236 16182
rect 6184 16118 6236 16124
rect 5906 15736 5962 15745
rect 5906 15671 5962 15680
rect 6092 15700 6144 15706
rect 5920 12753 5948 15671
rect 6092 15642 6144 15648
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 6012 14074 6040 15438
rect 6104 15094 6132 15642
rect 6196 15502 6224 16118
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6288 15706 6316 15846
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6380 15586 6408 15846
rect 6458 15736 6514 15745
rect 6458 15671 6514 15680
rect 6288 15558 6408 15586
rect 6472 15570 6500 15671
rect 6460 15564 6512 15570
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 6092 15088 6144 15094
rect 6092 15030 6144 15036
rect 6196 14822 6224 15438
rect 6288 15434 6316 15558
rect 6460 15506 6512 15512
rect 6276 15428 6328 15434
rect 6276 15370 6328 15376
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6380 14958 6408 15302
rect 6460 15020 6512 15026
rect 6460 14962 6512 14968
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6276 14884 6328 14890
rect 6276 14826 6328 14832
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6288 14770 6316 14826
rect 6288 14742 6408 14770
rect 6090 14104 6146 14113
rect 6000 14068 6052 14074
rect 6090 14039 6146 14048
rect 6000 14010 6052 14016
rect 6104 13938 6132 14039
rect 6182 13968 6238 13977
rect 6092 13932 6144 13938
rect 6182 13903 6238 13912
rect 6092 13874 6144 13880
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 5906 12744 5962 12753
rect 5906 12679 5962 12688
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5920 12170 5948 12582
rect 5908 12164 5960 12170
rect 5908 12106 5960 12112
rect 5906 11792 5962 11801
rect 5906 11727 5962 11736
rect 5920 11558 5948 11727
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5908 10464 5960 10470
rect 5906 10432 5908 10441
rect 5960 10432 5962 10441
rect 5906 10367 5962 10376
rect 6012 10010 6040 13670
rect 6092 13252 6144 13258
rect 6092 13194 6144 13200
rect 6104 12918 6132 13194
rect 6092 12912 6144 12918
rect 6092 12854 6144 12860
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 6104 12306 6132 12582
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6196 11558 6224 13903
rect 6276 13728 6328 13734
rect 6276 13670 6328 13676
rect 6288 13462 6316 13670
rect 6276 13456 6328 13462
rect 6380 13433 6408 14742
rect 6276 13398 6328 13404
rect 6366 13424 6422 13433
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6090 10704 6146 10713
rect 6090 10639 6146 10648
rect 6104 10538 6132 10639
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 6090 10296 6146 10305
rect 6196 10266 6224 10542
rect 6090 10231 6146 10240
rect 6184 10260 6236 10266
rect 6104 10146 6132 10231
rect 6184 10202 6236 10208
rect 6104 10118 6224 10146
rect 5920 9982 6040 10010
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 5920 7002 5948 9982
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 6012 8090 6040 9862
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6012 7206 6040 7686
rect 6104 7410 6132 9998
rect 6196 9178 6224 10118
rect 6288 9489 6316 13398
rect 6366 13359 6422 13368
rect 6380 12866 6408 13359
rect 6472 12986 6500 14962
rect 6564 13920 6592 17274
rect 6656 17066 6684 19994
rect 6736 19916 6788 19922
rect 6736 19858 6788 19864
rect 6748 18834 6776 19858
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6840 18329 6868 20182
rect 6920 19984 6972 19990
rect 6920 19926 6972 19932
rect 6826 18320 6882 18329
rect 6826 18255 6882 18264
rect 6932 18222 6960 19926
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6734 17912 6790 17921
rect 6734 17847 6790 17856
rect 6748 17746 6776 17847
rect 6736 17740 6788 17746
rect 6736 17682 6788 17688
rect 6840 17082 6868 18022
rect 6644 17060 6696 17066
rect 6644 17002 6696 17008
rect 6748 17054 6868 17082
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6656 15473 6684 16730
rect 6642 15464 6698 15473
rect 6642 15399 6698 15408
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6656 15026 6684 15302
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6748 14074 6776 17054
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6840 16794 6868 16934
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6736 13932 6788 13938
rect 6564 13892 6684 13920
rect 6552 13796 6604 13802
rect 6552 13738 6604 13744
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6380 12838 6500 12866
rect 6368 12708 6420 12714
rect 6368 12650 6420 12656
rect 6380 11898 6408 12650
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6472 11257 6500 12838
rect 6564 12782 6592 13738
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6656 12646 6684 13892
rect 6840 13920 6868 16594
rect 6932 16522 6960 16662
rect 6920 16516 6972 16522
rect 6920 16458 6972 16464
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6932 14618 6960 15914
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6788 13892 6868 13920
rect 6736 13874 6788 13880
rect 6734 13696 6790 13705
rect 6734 13631 6790 13640
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6458 11248 6514 11257
rect 6368 11212 6420 11218
rect 6458 11183 6514 11192
rect 6368 11154 6420 11160
rect 6274 9480 6330 9489
rect 6380 9450 6408 11154
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6274 9415 6330 9424
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6196 8634 6224 8978
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6196 8090 6224 8570
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 6182 7984 6238 7993
rect 6288 7954 6316 9318
rect 6380 9110 6408 9386
rect 6472 9178 6500 9454
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6564 9024 6592 12310
rect 6642 11928 6698 11937
rect 6642 11863 6698 11872
rect 6656 10266 6684 11863
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6656 9625 6684 9998
rect 6642 9616 6698 9625
rect 6642 9551 6698 9560
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6472 8996 6592 9024
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 6380 8294 6408 8842
rect 6472 8514 6500 8996
rect 6656 8922 6684 9454
rect 6564 8894 6684 8922
rect 6564 8634 6592 8894
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6656 8634 6684 8774
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6472 8486 6684 8514
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6368 8288 6420 8294
rect 6472 8265 6500 8366
rect 6552 8288 6604 8294
rect 6368 8230 6420 8236
rect 6458 8256 6514 8265
rect 6552 8230 6604 8236
rect 6458 8191 6514 8200
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6472 7993 6500 8026
rect 6458 7984 6514 7993
rect 6182 7919 6238 7928
rect 6276 7948 6328 7954
rect 6196 7585 6224 7919
rect 6458 7919 6514 7928
rect 6276 7890 6328 7896
rect 6182 7576 6238 7585
rect 6182 7511 6238 7520
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 5736 6956 5856 6984
rect 5908 6996 5960 7002
rect 5736 6497 5764 6956
rect 5908 6938 5960 6944
rect 6288 6934 6316 7890
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6366 7304 6422 7313
rect 6366 7239 6422 7248
rect 6380 7206 6408 7239
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6472 7002 6500 7482
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6184 6928 6236 6934
rect 6184 6870 6236 6876
rect 6276 6928 6328 6934
rect 6276 6870 6328 6876
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5722 6488 5778 6497
rect 5722 6423 5778 6432
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5736 6225 5764 6258
rect 5722 6216 5778 6225
rect 5722 6151 5778 6160
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5736 4690 5764 5646
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5632 4548 5684 4554
rect 5632 4490 5684 4496
rect 5446 4312 5502 4321
rect 5446 4247 5502 4256
rect 5460 3398 5488 4247
rect 5538 4040 5594 4049
rect 5538 3975 5594 3984
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5368 3182 5488 3210
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 5354 3088 5410 3097
rect 5172 2916 5224 2922
rect 5172 2858 5224 2864
rect 5276 2650 5304 3062
rect 5354 3023 5410 3032
rect 5368 2990 5396 3023
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 5460 2582 5488 3182
rect 5448 2576 5500 2582
rect 5448 2518 5500 2524
rect 5552 2446 5580 3975
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5000 1414 5120 1442
rect 5644 1442 5672 4490
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5736 1698 5764 4014
rect 5828 2650 5856 6802
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5920 4758 5948 6734
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 6012 5166 6040 6598
rect 6092 6180 6144 6186
rect 6092 6122 6144 6128
rect 6104 5914 6132 6122
rect 6196 5914 6224 6870
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6288 6390 6316 6598
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 6104 4604 6132 5578
rect 6276 5296 6328 5302
rect 6380 5250 6408 6938
rect 6564 6322 6592 8230
rect 6656 7041 6684 8486
rect 6642 7032 6698 7041
rect 6642 6967 6698 6976
rect 6656 6390 6684 6967
rect 6748 6866 6776 13631
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6840 12714 6868 12922
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 6932 12322 6960 14418
rect 7024 12617 7052 22320
rect 7392 22273 7420 22320
rect 7378 22264 7434 22273
rect 7378 22199 7434 22208
rect 7104 19984 7156 19990
rect 7104 19926 7156 19932
rect 7472 19984 7524 19990
rect 7472 19926 7524 19932
rect 7116 19530 7144 19926
rect 7116 19514 7236 19530
rect 7116 19508 7248 19514
rect 7116 19502 7196 19508
rect 7116 19310 7144 19502
rect 7196 19450 7248 19456
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7116 18834 7144 19246
rect 7104 18828 7156 18834
rect 7104 18770 7156 18776
rect 7116 18154 7144 18770
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7288 18352 7340 18358
rect 7288 18294 7340 18300
rect 7104 18148 7156 18154
rect 7104 18090 7156 18096
rect 7194 18048 7250 18057
rect 7194 17983 7250 17992
rect 7208 17320 7236 17983
rect 7300 17513 7328 18294
rect 7286 17504 7342 17513
rect 7286 17439 7342 17448
rect 7116 17292 7236 17320
rect 7010 12608 7066 12617
rect 7010 12543 7066 12552
rect 7116 12442 7144 17292
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7208 16454 7236 17138
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7208 15978 7236 16390
rect 7196 15972 7248 15978
rect 7196 15914 7248 15920
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7196 15564 7248 15570
rect 7300 15552 7328 15846
rect 7248 15524 7328 15552
rect 7196 15506 7248 15512
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7208 12986 7236 15098
rect 7286 15056 7342 15065
rect 7286 14991 7342 15000
rect 7300 14550 7328 14991
rect 7288 14544 7340 14550
rect 7288 14486 7340 14492
rect 7300 13870 7328 14486
rect 7392 14414 7420 18566
rect 7484 18426 7512 19926
rect 7760 19394 7788 22320
rect 8128 20346 8156 22320
rect 8128 20318 8248 20346
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7668 19366 7788 19394
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7484 16726 7512 17614
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7484 15910 7512 16526
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7470 15736 7526 15745
rect 7470 15671 7526 15680
rect 7484 15570 7512 15671
rect 7472 15564 7524 15570
rect 7472 15506 7524 15512
rect 7576 14521 7604 18226
rect 7562 14512 7618 14521
rect 7668 14482 7696 19366
rect 7748 19236 7800 19242
rect 7748 19178 7800 19184
rect 7760 18680 7788 19178
rect 8220 19122 8248 20318
rect 8298 19952 8354 19961
rect 8298 19887 8354 19896
rect 8392 19916 8444 19922
rect 8312 19242 8340 19887
rect 8392 19858 8444 19864
rect 8404 19786 8432 19858
rect 8392 19780 8444 19786
rect 8392 19722 8444 19728
rect 8404 19514 8432 19722
rect 8392 19508 8444 19514
rect 8392 19450 8444 19456
rect 8300 19236 8352 19242
rect 8300 19178 8352 19184
rect 8392 19168 8444 19174
rect 8220 19094 8340 19122
rect 8392 19110 8444 19116
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 8206 19000 8262 19009
rect 8128 18944 8206 18952
rect 8128 18935 8262 18944
rect 8128 18924 8248 18935
rect 7760 18652 7880 18680
rect 7852 18612 7880 18652
rect 8024 18624 8076 18630
rect 7746 18592 7802 18601
rect 7746 18527 7802 18536
rect 7852 18584 8024 18612
rect 7760 18358 7788 18527
rect 7748 18352 7800 18358
rect 7748 18294 7800 18300
rect 7852 18272 7880 18584
rect 8024 18566 8076 18572
rect 8022 18456 8078 18465
rect 8128 18442 8156 18924
rect 8078 18414 8156 18442
rect 8022 18391 8078 18400
rect 8116 18284 8168 18290
rect 7852 18244 8116 18272
rect 8116 18226 8168 18232
rect 8312 18170 8340 19094
rect 8404 18902 8432 19110
rect 8392 18896 8444 18902
rect 8392 18838 8444 18844
rect 8496 18737 8524 22320
rect 8760 21140 8812 21146
rect 8760 21082 8812 21088
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 8482 18728 8538 18737
rect 8482 18663 8538 18672
rect 8588 18612 8616 20402
rect 8666 19544 8722 19553
rect 8666 19479 8722 19488
rect 8680 19310 8708 19479
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 7748 18148 7800 18154
rect 7748 18090 7800 18096
rect 8220 18142 8340 18170
rect 8496 18584 8616 18612
rect 7760 16590 7788 18090
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 7932 17808 7984 17814
rect 7932 17750 7984 17756
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 7852 17270 7880 17682
rect 7944 17338 7972 17750
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 7840 17264 7892 17270
rect 7840 17206 7892 17212
rect 8024 17264 8076 17270
rect 8024 17206 8076 17212
rect 8036 17105 8064 17206
rect 8022 17096 8078 17105
rect 8022 17031 8078 17040
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7760 16250 7788 16526
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7760 15348 7788 16186
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 7840 15360 7892 15366
rect 7760 15320 7840 15348
rect 7760 15065 7788 15320
rect 8116 15360 8168 15366
rect 7840 15302 7892 15308
rect 7930 15328 7986 15337
rect 8116 15302 8168 15308
rect 7930 15263 7986 15272
rect 7746 15056 7802 15065
rect 7746 14991 7802 15000
rect 7944 14958 7972 15263
rect 8128 15094 8156 15302
rect 8116 15088 8168 15094
rect 8116 15030 8168 15036
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 7760 14550 7788 14894
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 7930 14512 7986 14521
rect 7562 14447 7618 14456
rect 7656 14476 7708 14482
rect 7930 14447 7932 14456
rect 7656 14418 7708 14424
rect 7984 14447 7986 14456
rect 7932 14418 7984 14424
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7300 13462 7328 13806
rect 7392 13530 7420 14350
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7288 13456 7340 13462
rect 7288 13398 7340 13404
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7196 12776 7248 12782
rect 7300 12753 7328 13262
rect 7484 12986 7512 14214
rect 8128 14113 8156 14350
rect 8114 14104 8170 14113
rect 8114 14039 8170 14048
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7840 13456 7892 13462
rect 7840 13398 7892 13404
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7196 12718 7248 12724
rect 7286 12744 7342 12753
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7116 12345 7144 12378
rect 6840 12294 6960 12322
rect 7102 12336 7158 12345
rect 6840 11642 6868 12294
rect 7102 12271 7158 12280
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6932 11762 6960 12174
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6840 11614 7052 11642
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 10305 6868 11494
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6826 10296 6882 10305
rect 6826 10231 6882 10240
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6840 7342 6868 9862
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6932 7274 6960 10542
rect 7024 10305 7052 11614
rect 7116 11082 7144 12106
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7010 10296 7066 10305
rect 7010 10231 7066 10240
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6644 6384 6696 6390
rect 6644 6326 6696 6332
rect 6840 6322 6868 6734
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6564 5953 6592 6258
rect 6644 6112 6696 6118
rect 6642 6080 6644 6089
rect 6696 6080 6698 6089
rect 6642 6015 6698 6024
rect 6550 5944 6606 5953
rect 6550 5879 6606 5888
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6328 5244 6408 5250
rect 6276 5238 6408 5244
rect 6288 5222 6408 5238
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 5920 4576 6132 4604
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 5920 2378 5948 4576
rect 5998 4312 6054 4321
rect 5998 4247 6054 4256
rect 6012 4214 6040 4247
rect 6000 4208 6052 4214
rect 6000 4150 6052 4156
rect 5998 4040 6054 4049
rect 5998 3975 6000 3984
rect 6052 3975 6054 3984
rect 6000 3946 6052 3952
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6012 3126 6040 3470
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 6104 2990 6132 3334
rect 6196 3194 6224 5102
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6288 3194 6316 4694
rect 6380 4214 6408 5222
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6288 3058 6316 3130
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 6196 2650 6224 2790
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 6092 2576 6144 2582
rect 6092 2518 6144 2524
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 5724 1692 5776 1698
rect 5724 1634 5776 1640
rect 5356 1420 5408 1426
rect 5000 480 5028 1414
rect 5644 1414 5764 1442
rect 5356 1362 5408 1368
rect 5368 480 5396 1362
rect 5736 480 5764 1414
rect 6104 513 6132 2518
rect 6380 2009 6408 3538
rect 6472 3505 6500 5714
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6458 3496 6514 3505
rect 6458 3431 6514 3440
rect 6366 2000 6422 2009
rect 6366 1935 6422 1944
rect 6564 1902 6592 4014
rect 6656 2582 6684 6015
rect 6826 5944 6882 5953
rect 6826 5879 6882 5888
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6748 5098 6776 5646
rect 6840 5166 6868 5879
rect 7024 5710 7052 10066
rect 7116 8362 7144 11018
rect 7208 10266 7236 12718
rect 7484 12714 7512 12922
rect 7286 12679 7342 12688
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7300 11218 7328 12582
rect 7378 12472 7434 12481
rect 7668 12442 7696 13126
rect 7378 12407 7380 12416
rect 7432 12407 7434 12416
rect 7656 12436 7708 12442
rect 7380 12378 7432 12384
rect 7656 12378 7708 12384
rect 7654 12336 7710 12345
rect 7564 12300 7616 12306
rect 7654 12271 7710 12280
rect 7564 12242 7616 12248
rect 7470 12064 7526 12073
rect 7470 11999 7526 12008
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7392 11082 7420 11834
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7484 10962 7512 11999
rect 7392 10934 7512 10962
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7208 9450 7236 10202
rect 7300 9994 7328 10610
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7300 9450 7328 9930
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7194 9072 7250 9081
rect 7194 9007 7250 9016
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 7208 7426 7236 9007
rect 7300 7750 7328 9386
rect 7392 7834 7420 10934
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7484 10033 7512 10746
rect 7470 10024 7526 10033
rect 7470 9959 7472 9968
rect 7524 9959 7526 9968
rect 7472 9930 7524 9936
rect 7484 9899 7512 9930
rect 7470 9616 7526 9625
rect 7470 9551 7526 9560
rect 7484 9178 7512 9551
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7470 8664 7526 8673
rect 7470 8599 7526 8608
rect 7484 7954 7512 8599
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7392 7806 7512 7834
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7116 7398 7236 7426
rect 7286 7440 7342 7449
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7116 5522 7144 7398
rect 7286 7375 7342 7384
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7208 7002 7236 7278
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7208 5953 7236 6938
rect 7194 5944 7250 5953
rect 7300 5914 7328 7375
rect 7392 7002 7420 7686
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7484 6644 7512 7806
rect 7576 6798 7604 12242
rect 7668 7954 7696 12271
rect 7760 11121 7788 13330
rect 7852 12714 7880 13398
rect 7840 12708 7892 12714
rect 7840 12650 7892 12656
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 8116 12368 8168 12374
rect 7930 12336 7986 12345
rect 8116 12310 8168 12316
rect 7930 12271 7986 12280
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7852 11898 7880 12174
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7944 11830 7972 12271
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 8128 11762 8156 12310
rect 8220 12186 8248 18142
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8312 17921 8340 18022
rect 8298 17912 8354 17921
rect 8298 17847 8354 17856
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 8312 16726 8340 17614
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8312 15434 8340 16662
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 8312 13326 8340 14214
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8312 12374 8340 12582
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8220 12158 8340 12186
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8116 11756 8168 11762
rect 8116 11698 8168 11704
rect 8220 11694 8248 12038
rect 8312 11801 8340 12158
rect 8404 11898 8432 17138
rect 8496 16153 8524 18584
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 8588 17882 8616 18090
rect 8680 18057 8708 18770
rect 8666 18048 8722 18057
rect 8666 17983 8722 17992
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 8668 16720 8720 16726
rect 8668 16662 8720 16668
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8482 16144 8538 16153
rect 8482 16079 8538 16088
rect 8482 15192 8538 15201
rect 8482 15127 8538 15136
rect 8496 14550 8524 15127
rect 8588 14618 8616 16594
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8484 14544 8536 14550
rect 8484 14486 8536 14492
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8496 12918 8524 13262
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8588 12186 8616 14350
rect 8680 12424 8708 16662
rect 8772 16114 8800 21082
rect 8850 19136 8906 19145
rect 8850 19071 8906 19080
rect 8864 18465 8892 19071
rect 8850 18456 8906 18465
rect 8850 18391 8906 18400
rect 8852 18080 8904 18086
rect 8852 18022 8904 18028
rect 8864 17338 8892 18022
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8956 17218 8984 22320
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 9048 18426 9076 19790
rect 9220 19780 9272 19786
rect 9220 19722 9272 19728
rect 9232 19666 9260 19722
rect 9140 19638 9260 19666
rect 9140 18766 9168 19638
rect 9218 19408 9274 19417
rect 9218 19343 9274 19352
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9036 18080 9088 18086
rect 9036 18022 9088 18028
rect 9048 17921 9076 18022
rect 9034 17912 9090 17921
rect 9034 17847 9090 17856
rect 9140 17678 9168 18702
rect 9232 17882 9260 19343
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 9220 17740 9272 17746
rect 9220 17682 9272 17688
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 8864 17202 8984 17218
rect 9140 17202 9168 17614
rect 8852 17196 8984 17202
rect 8904 17190 8984 17196
rect 9128 17196 9180 17202
rect 8852 17138 8904 17144
rect 9128 17138 9180 17144
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8864 16250 8892 16934
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8944 16040 8996 16046
rect 8850 16008 8906 16017
rect 8944 15982 8996 15988
rect 8850 15943 8906 15952
rect 8864 15910 8892 15943
rect 8852 15904 8904 15910
rect 8758 15872 8814 15881
rect 8852 15846 8904 15852
rect 8758 15807 8814 15816
rect 8772 15722 8800 15807
rect 8772 15694 8892 15722
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 8772 14414 8800 15302
rect 8864 14618 8892 15694
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8864 13734 8892 13806
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8772 12986 8800 13330
rect 8956 13297 8984 15982
rect 8942 13288 8998 13297
rect 8942 13223 8998 13232
rect 9048 13002 9076 16594
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 9140 15502 9168 15914
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9140 14414 9168 15438
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 8760 12980 8812 12986
rect 9048 12974 9168 13002
rect 8760 12922 8812 12928
rect 9036 12912 9088 12918
rect 9036 12854 9088 12860
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8956 12442 8984 12582
rect 8944 12436 8996 12442
rect 8680 12396 8800 12424
rect 8668 12300 8720 12306
rect 8668 12242 8720 12248
rect 8496 12158 8616 12186
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8298 11792 8354 11801
rect 8298 11727 8354 11736
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 7840 11688 7892 11694
rect 7838 11656 7840 11665
rect 8208 11688 8260 11694
rect 7892 11656 7894 11665
rect 8208 11630 8260 11636
rect 7838 11591 7894 11600
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8312 11132 8340 11290
rect 8404 11286 8432 11698
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 8496 11218 8524 12158
rect 8576 12096 8628 12102
rect 8574 12064 8576 12073
rect 8628 12064 8630 12073
rect 8574 11999 8630 12008
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8392 11144 8444 11150
rect 7746 11112 7802 11121
rect 7746 11047 7802 11056
rect 8206 11112 8262 11121
rect 8312 11104 8392 11132
rect 8392 11086 8444 11092
rect 8206 11047 8262 11056
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7760 10130 7788 10950
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 8220 10266 8248 11047
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8390 10432 8446 10441
rect 8312 10266 8340 10406
rect 8390 10367 8446 10376
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 7838 10160 7894 10169
rect 7748 10124 7800 10130
rect 7838 10095 7894 10104
rect 8024 10124 8076 10130
rect 7748 10066 7800 10072
rect 7852 9994 7880 10095
rect 8024 10066 8076 10072
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 7840 9988 7892 9994
rect 7840 9930 7892 9936
rect 8036 9489 8064 10066
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8022 9480 8078 9489
rect 8022 9415 8078 9424
rect 8128 9364 8156 9930
rect 8128 9336 8248 9364
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 7748 9172 7800 9178
rect 7800 9132 7880 9160
rect 7748 9114 7800 9120
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7760 8634 7788 8978
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7760 7886 7788 8570
rect 7852 8566 7880 9132
rect 8220 8634 8248 9336
rect 8312 8673 8340 10066
rect 8404 9994 8432 10367
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8404 9217 8432 9318
rect 8390 9208 8446 9217
rect 8390 9143 8446 9152
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8298 8664 8354 8673
rect 8208 8628 8260 8634
rect 8298 8599 8354 8608
rect 8208 8570 8260 8576
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 8404 8498 8432 8978
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8220 8072 8248 8434
rect 8496 8378 8524 11154
rect 8588 10305 8616 11834
rect 8680 10810 8708 12242
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8666 10432 8722 10441
rect 8666 10367 8722 10376
rect 8574 10296 8630 10305
rect 8574 10231 8630 10240
rect 8588 8838 8616 10231
rect 8680 10130 8708 10367
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8772 10062 8800 12396
rect 8944 12378 8996 12384
rect 9048 12345 9076 12854
rect 9034 12336 9090 12345
rect 9034 12271 9090 12280
rect 9048 12238 9076 12271
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 8864 11393 8892 12174
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 8850 11384 8906 11393
rect 8850 11319 8906 11328
rect 8942 11248 8998 11257
rect 8942 11183 8998 11192
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 8864 10713 8892 10950
rect 8850 10704 8906 10713
rect 8850 10639 8906 10648
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8864 10062 8892 10542
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8574 8664 8630 8673
rect 8574 8599 8630 8608
rect 8588 8498 8616 8599
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8404 8350 8524 8378
rect 8128 8044 8248 8072
rect 8300 8084 8352 8090
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7748 7880 7800 7886
rect 7654 7848 7710 7857
rect 7748 7822 7800 7828
rect 7654 7783 7710 7792
rect 7668 7002 7696 7783
rect 7760 7342 7788 7822
rect 7852 7546 7880 7890
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 8128 7342 8156 8044
rect 8300 8026 8352 8032
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8220 7546 8248 7890
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8312 7410 8340 8026
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 7852 7188 7880 7278
rect 7760 7160 7880 7188
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7760 6934 7788 7160
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7748 6928 7800 6934
rect 7748 6870 7800 6876
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8036 6662 8064 6734
rect 8024 6656 8076 6662
rect 7484 6616 7604 6644
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7194 5879 7250 5888
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7392 5778 7420 6054
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7300 5658 7328 5714
rect 7300 5630 7420 5658
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6736 5092 6788 5098
rect 6736 5034 6788 5040
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6644 2576 6696 2582
rect 6644 2518 6696 2524
rect 6552 1896 6604 1902
rect 6552 1838 6604 1844
rect 6182 1592 6238 1601
rect 6182 1527 6238 1536
rect 6090 504 6146 513
rect 3974 232 4030 241
rect 3974 167 4030 176
rect 4250 0 4306 480
rect 4618 0 4674 480
rect 4986 0 5042 480
rect 5354 0 5410 480
rect 5722 0 5778 480
rect 6196 480 6224 1527
rect 6748 1170 6776 4150
rect 6840 2990 6868 5102
rect 7024 4146 7052 5510
rect 7116 5494 7328 5522
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 7116 4826 7144 5034
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7208 4078 7236 5306
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 6920 3392 6972 3398
rect 7024 3369 7052 3674
rect 7300 3670 7328 5494
rect 7392 4826 7420 5630
rect 7472 5092 7524 5098
rect 7472 5034 7524 5040
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7104 3664 7156 3670
rect 7104 3606 7156 3612
rect 7288 3664 7340 3670
rect 7380 3664 7432 3670
rect 7288 3606 7340 3612
rect 7378 3632 7380 3641
rect 7432 3632 7434 3641
rect 6920 3334 6972 3340
rect 7010 3360 7066 3369
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6840 2854 6868 2926
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6564 1142 6776 1170
rect 6564 480 6592 1142
rect 6932 480 6960 3334
rect 7010 3295 7066 3304
rect 7024 2038 7052 3295
rect 7116 2689 7144 3606
rect 7378 3567 7434 3576
rect 7484 3233 7512 5034
rect 7576 4078 7604 6616
rect 8024 6598 8076 6604
rect 7654 6488 7710 6497
rect 7654 6423 7710 6432
rect 7668 6390 7696 6423
rect 8128 6390 8156 6870
rect 7656 6384 7708 6390
rect 8024 6384 8076 6390
rect 7656 6326 7708 6332
rect 7930 6352 7986 6361
rect 8024 6326 8076 6332
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 7930 6287 7986 6296
rect 7944 6254 7972 6287
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 8036 6186 8064 6326
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7760 4826 7788 6054
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7852 5137 7880 5510
rect 8128 5234 8156 5578
rect 8220 5370 8248 7346
rect 8404 6338 8432 8350
rect 8680 8294 8708 9658
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8312 6310 8432 6338
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 7838 5128 7894 5137
rect 7838 5063 7894 5072
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7668 3398 7696 4490
rect 8220 4214 8248 5306
rect 8312 4554 8340 6310
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8404 5710 8432 6190
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8404 4622 8432 5646
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8220 3720 8248 4014
rect 8128 3692 8248 3720
rect 8024 3664 8076 3670
rect 8024 3606 8076 3612
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7470 3224 7526 3233
rect 8036 3176 8064 3606
rect 7470 3159 7526 3168
rect 7576 3148 8064 3176
rect 7102 2680 7158 2689
rect 7102 2615 7158 2624
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 7012 2032 7064 2038
rect 7012 1974 7064 1980
rect 7208 1494 7236 2450
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7392 2145 7420 2382
rect 7378 2136 7434 2145
rect 7378 2071 7434 2080
rect 7286 1728 7342 1737
rect 7286 1663 7342 1672
rect 7196 1488 7248 1494
rect 7196 1430 7248 1436
rect 7208 1222 7236 1430
rect 7196 1216 7248 1222
rect 7196 1158 7248 1164
rect 7300 480 7328 1663
rect 7392 1154 7420 2071
rect 7576 1630 7604 3148
rect 8128 3058 8156 3692
rect 8312 3398 8340 4150
rect 8404 3534 8432 4558
rect 8496 3602 8524 8230
rect 8772 7936 8800 9998
rect 8956 9489 8984 11183
rect 9048 10674 9076 11834
rect 9140 11558 9168 12974
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9034 10432 9090 10441
rect 9034 10367 9090 10376
rect 9048 10266 9076 10367
rect 9036 10260 9088 10266
rect 9140 10248 9168 11494
rect 9232 10849 9260 17682
rect 9324 16658 9352 22320
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9416 18850 9444 20334
rect 9692 19990 9720 22320
rect 9680 19984 9732 19990
rect 9680 19926 9732 19932
rect 10060 19718 10088 22320
rect 10232 20052 10284 20058
rect 10232 19994 10284 20000
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9508 18970 9536 19450
rect 9692 19310 9720 19654
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9588 19236 9640 19242
rect 9588 19178 9640 19184
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 9600 18902 9628 19178
rect 9784 19122 9812 19654
rect 9956 19236 10008 19242
rect 9956 19178 10008 19184
rect 9692 19094 9812 19122
rect 9588 18896 9640 18902
rect 9416 18822 9536 18850
rect 9692 18873 9720 19094
rect 9588 18838 9640 18844
rect 9678 18864 9734 18873
rect 9402 18456 9458 18465
rect 9402 18391 9458 18400
rect 9416 18222 9444 18391
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9508 17513 9536 18822
rect 9600 18290 9628 18838
rect 9968 18834 9996 19178
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 10060 18970 10088 19110
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 9864 18828 9916 18834
rect 9678 18799 9734 18808
rect 9784 18788 9864 18816
rect 9784 18578 9812 18788
rect 9864 18770 9916 18776
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9784 18550 9996 18578
rect 9770 18456 9826 18465
rect 9770 18391 9826 18400
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9494 17504 9550 17513
rect 9494 17439 9550 17448
rect 9600 17202 9628 18226
rect 9784 17814 9812 18391
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9876 17921 9904 18022
rect 9862 17912 9918 17921
rect 9862 17847 9918 17856
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9508 16726 9536 16934
rect 9600 16794 9628 17138
rect 9680 17060 9732 17066
rect 9680 17002 9732 17008
rect 9692 16969 9720 17002
rect 9678 16960 9734 16969
rect 9678 16895 9734 16904
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9600 16114 9628 16730
rect 9312 16108 9364 16114
rect 9588 16108 9640 16114
rect 9312 16050 9364 16056
rect 9508 16068 9588 16096
rect 9324 13512 9352 16050
rect 9508 15434 9536 16068
rect 9588 16050 9640 16056
rect 9680 15904 9732 15910
rect 9784 15892 9812 17274
rect 9732 15864 9812 15892
rect 9680 15846 9732 15852
rect 9678 15736 9734 15745
rect 9678 15671 9680 15680
rect 9732 15671 9734 15680
rect 9680 15642 9732 15648
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9416 13705 9444 14758
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9508 13870 9536 14554
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9402 13696 9458 13705
rect 9402 13631 9458 13640
rect 9324 13484 9444 13512
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 9324 12481 9352 13330
rect 9416 13190 9444 13484
rect 9508 13326 9536 13806
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9310 12472 9366 12481
rect 9310 12407 9366 12416
rect 9310 12200 9366 12209
rect 9310 12135 9366 12144
rect 9324 11830 9352 12135
rect 9312 11824 9364 11830
rect 9312 11766 9364 11772
rect 9416 11393 9444 12718
rect 9600 12481 9628 15506
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9692 14074 9720 14826
rect 9784 14482 9812 15864
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9692 13938 9720 14010
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9586 12472 9642 12481
rect 9586 12407 9642 12416
rect 9496 12368 9548 12374
rect 9784 12356 9812 14418
rect 9876 14414 9904 17478
rect 9968 16658 9996 18550
rect 10152 18426 10180 19858
rect 10244 18902 10272 19994
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 10336 19446 10364 19858
rect 10324 19440 10376 19446
rect 10324 19382 10376 19388
rect 10324 19168 10376 19174
rect 10324 19110 10376 19116
rect 10232 18896 10284 18902
rect 10232 18838 10284 18844
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10138 18320 10194 18329
rect 10336 18306 10364 19110
rect 10138 18255 10194 18264
rect 10244 18278 10364 18306
rect 10428 18290 10456 22320
rect 10508 21412 10560 21418
rect 10508 21354 10560 21360
rect 10520 19174 10548 21354
rect 10796 20398 10824 22320
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10876 20324 10928 20330
rect 10876 20266 10928 20272
rect 10888 19922 10916 20266
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 10876 19916 10928 19922
rect 10876 19858 10928 19864
rect 10600 19712 10652 19718
rect 10600 19654 10652 19660
rect 10508 19168 10560 19174
rect 10508 19110 10560 19116
rect 10508 18692 10560 18698
rect 10508 18634 10560 18640
rect 10416 18284 10468 18290
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 10060 16833 10088 17682
rect 10046 16824 10102 16833
rect 10046 16759 10102 16768
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9496 12310 9548 12316
rect 9600 12328 9812 12356
rect 9402 11384 9458 11393
rect 9508 11354 9536 12310
rect 9402 11319 9458 11328
rect 9496 11348 9548 11354
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 9416 11234 9444 11319
rect 9496 11290 9548 11296
rect 9218 10840 9274 10849
rect 9324 10810 9352 11222
rect 9416 11206 9536 11234
rect 9218 10775 9274 10784
rect 9312 10804 9364 10810
rect 9232 10577 9260 10775
rect 9312 10746 9364 10752
rect 9218 10568 9274 10577
rect 9218 10503 9274 10512
rect 9402 10432 9458 10441
rect 9402 10367 9458 10376
rect 9140 10220 9260 10248
rect 9036 10202 9088 10208
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 8942 9480 8998 9489
rect 8852 9444 8904 9450
rect 8942 9415 8998 9424
rect 8852 9386 8904 9392
rect 8864 9110 8892 9386
rect 8852 9104 8904 9110
rect 8852 9046 8904 9052
rect 8864 8974 8892 9046
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8864 8430 8892 8774
rect 8947 8650 8975 8842
rect 9048 8809 9076 9998
rect 9140 9722 9168 9998
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9232 9568 9260 10220
rect 9140 9540 9260 9568
rect 9034 8800 9090 8809
rect 9034 8735 9090 8744
rect 8947 8622 9076 8650
rect 9048 8498 9076 8622
rect 9140 8548 9168 9540
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9220 9444 9272 9450
rect 9220 9386 9272 9392
rect 9232 9178 9260 9386
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9232 8906 9260 9114
rect 9324 9110 9352 9454
rect 9312 9104 9364 9110
rect 9312 9046 9364 9052
rect 9220 8900 9272 8906
rect 9220 8842 9272 8848
rect 9140 8520 9352 8548
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 8852 8288 8904 8294
rect 8904 8248 8984 8276
rect 8852 8230 8904 8236
rect 8772 7908 8892 7936
rect 8864 7834 8892 7908
rect 8772 7806 8892 7834
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8588 7002 8616 7278
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8680 6934 8708 7482
rect 8668 6928 8720 6934
rect 8668 6870 8720 6876
rect 8574 6352 8630 6361
rect 8574 6287 8576 6296
rect 8628 6287 8630 6296
rect 8576 6258 8628 6264
rect 8574 6216 8630 6225
rect 8574 6151 8576 6160
rect 8628 6151 8630 6160
rect 8576 6122 8628 6128
rect 8574 5944 8630 5953
rect 8574 5879 8576 5888
rect 8628 5879 8630 5888
rect 8576 5850 8628 5856
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8574 4448 8630 4457
rect 8574 4383 8630 4392
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8588 3534 8616 4383
rect 8392 3528 8444 3534
rect 8576 3528 8628 3534
rect 8392 3470 8444 3476
rect 8482 3496 8538 3505
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8298 3224 8354 3233
rect 8208 3188 8260 3194
rect 8298 3159 8354 3168
rect 8208 3130 8260 3136
rect 7840 3052 7892 3058
rect 7760 3012 7840 3040
rect 7760 2854 7788 3012
rect 7840 2994 7892 3000
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 7564 1624 7616 1630
rect 7564 1566 7616 1572
rect 7380 1148 7432 1154
rect 7380 1090 7432 1096
rect 7668 480 7696 2518
rect 7760 1766 7788 2586
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 7852 1766 7880 2246
rect 8220 2038 8248 3130
rect 8312 2650 8340 3159
rect 8404 2854 8432 3470
rect 8576 3470 8628 3476
rect 8482 3431 8538 3440
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8496 2666 8524 3431
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8404 2638 8524 2666
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8208 2032 8260 2038
rect 8208 1974 8260 1980
rect 8312 1970 8340 2382
rect 8300 1964 8352 1970
rect 8300 1906 8352 1912
rect 7748 1760 7800 1766
rect 7748 1702 7800 1708
rect 7840 1760 7892 1766
rect 7840 1702 7892 1708
rect 8022 1592 8078 1601
rect 8022 1527 8078 1536
rect 8036 480 8064 1527
rect 8404 480 8432 2638
rect 8588 2446 8616 2790
rect 8680 2650 8708 5170
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8772 1630 8800 7806
rect 8850 7576 8906 7585
rect 8850 7511 8906 7520
rect 8864 7313 8892 7511
rect 8850 7304 8906 7313
rect 8850 7239 8906 7248
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8864 5098 8892 7142
rect 8852 5092 8904 5098
rect 8852 5034 8904 5040
rect 8850 4992 8906 5001
rect 8956 4978 8984 8248
rect 9140 8090 9168 8366
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9140 7750 9168 8026
rect 9324 7857 9352 8520
rect 9310 7848 9366 7857
rect 9220 7812 9272 7818
rect 9310 7783 9366 7792
rect 9220 7754 9272 7760
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9232 7546 9260 7754
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9220 7404 9272 7410
rect 9324 7392 9352 7686
rect 9416 7585 9444 10367
rect 9508 8129 9536 11206
rect 9494 8120 9550 8129
rect 9494 8055 9550 8064
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9600 7834 9628 12328
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 9784 11354 9812 12106
rect 9876 11898 9904 13398
rect 9968 12481 9996 15438
rect 9954 12472 10010 12481
rect 9954 12407 10010 12416
rect 10060 12288 10088 15914
rect 10152 12481 10180 18255
rect 10244 14618 10272 18278
rect 10416 18226 10468 18232
rect 10520 18222 10548 18634
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10336 17746 10364 18158
rect 10416 18148 10468 18154
rect 10416 18090 10468 18096
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10428 16998 10456 18090
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10322 16688 10378 16697
rect 10322 16623 10378 16632
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10244 13326 10272 13874
rect 10336 13734 10364 16623
rect 10520 16590 10548 18158
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10520 16046 10548 16526
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10520 15638 10548 15982
rect 10508 15632 10560 15638
rect 10508 15574 10560 15580
rect 10324 13728 10376 13734
rect 10376 13688 10456 13716
rect 10324 13670 10376 13676
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10322 13288 10378 13297
rect 10322 13223 10324 13232
rect 10376 13223 10378 13232
rect 10324 13194 10376 13200
rect 10336 12782 10364 13194
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10428 12628 10456 13688
rect 10612 13444 10640 19654
rect 10782 19544 10838 19553
rect 10782 19479 10838 19488
rect 10796 18766 10824 19479
rect 10888 19417 10916 19858
rect 10874 19408 10930 19417
rect 10874 19343 10930 19352
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 10690 18592 10746 18601
rect 10690 18527 10746 18536
rect 10704 16969 10732 18527
rect 10796 18465 10824 18702
rect 10782 18456 10838 18465
rect 10782 18391 10838 18400
rect 10782 18320 10838 18329
rect 10782 18255 10838 18264
rect 10796 17134 10824 18255
rect 10888 17338 10916 19343
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10690 16960 10746 16969
rect 10746 16918 10824 16946
rect 10690 16895 10746 16904
rect 10692 16448 10744 16454
rect 10690 16416 10692 16425
rect 10744 16416 10746 16425
rect 10690 16351 10746 16360
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10520 13416 10640 13444
rect 10520 13025 10548 13416
rect 10600 13320 10652 13326
rect 10704 13308 10732 15506
rect 10652 13280 10732 13308
rect 10600 13262 10652 13268
rect 10506 13016 10562 13025
rect 10506 12951 10508 12960
rect 10560 12951 10562 12960
rect 10508 12922 10560 12928
rect 10520 12891 10548 12922
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10244 12600 10456 12628
rect 10138 12472 10194 12481
rect 10138 12407 10194 12416
rect 10060 12260 10180 12288
rect 10046 12200 10102 12209
rect 10046 12135 10102 12144
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 10060 11665 10088 12135
rect 10046 11656 10102 11665
rect 10046 11591 10102 11600
rect 10060 11558 10088 11591
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9692 8022 9720 9862
rect 9784 9586 9812 10542
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9876 9926 9904 10066
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9862 9752 9918 9761
rect 9862 9687 9918 9696
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9876 9518 9904 9687
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 9402 7576 9458 7585
rect 9508 7546 9536 7822
rect 9600 7806 9720 7834
rect 9402 7511 9458 7520
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9272 7364 9352 7392
rect 9404 7404 9456 7410
rect 9220 7346 9272 7352
rect 9456 7364 9536 7392
rect 9404 7346 9456 7352
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 9404 7268 9456 7274
rect 9404 7210 9456 7216
rect 9048 7002 9076 7210
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 9416 6780 9444 7210
rect 9508 6866 9536 7364
rect 9600 7002 9628 7482
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9140 6752 9444 6780
rect 9036 6384 9088 6390
rect 9036 6326 9088 6332
rect 9048 5778 9076 6326
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 9048 5370 9076 5714
rect 9140 5370 9168 6752
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9232 6254 9260 6598
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9324 6118 9352 6598
rect 9402 6352 9458 6361
rect 9402 6287 9458 6296
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 8906 4950 8984 4978
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 8850 4927 8906 4936
rect 8864 4826 8892 4927
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8852 4548 8904 4554
rect 8904 4508 8984 4536
rect 8852 4490 8904 4496
rect 8850 4176 8906 4185
rect 8850 4111 8906 4120
rect 8864 3516 8892 4111
rect 8956 3670 8984 4508
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8864 3488 8984 3516
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8864 3097 8892 3130
rect 8850 3088 8906 3097
rect 8850 3023 8906 3032
rect 8760 1624 8812 1630
rect 8760 1566 8812 1572
rect 8956 1306 8984 3488
rect 9048 1970 9076 4966
rect 9140 3369 9168 5306
rect 9126 3360 9182 3369
rect 9126 3295 9182 3304
rect 9324 3233 9352 5850
rect 9416 5409 9444 6287
rect 9508 6186 9536 6802
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9600 6089 9628 6734
rect 9586 6080 9642 6089
rect 9586 6015 9642 6024
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9402 5400 9458 5409
rect 9402 5335 9458 5344
rect 9600 5166 9628 5510
rect 9588 5160 9640 5166
rect 9692 5137 9720 7806
rect 9784 6662 9812 9386
rect 9968 9110 9996 9998
rect 9956 9104 10008 9110
rect 9956 9046 10008 9052
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9876 8922 9904 8978
rect 9876 8894 9996 8922
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9876 8566 9904 8774
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9968 8412 9996 8894
rect 9876 8384 9996 8412
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9876 6474 9904 8384
rect 10060 8378 10088 11494
rect 10152 10849 10180 12260
rect 10138 10840 10194 10849
rect 10138 10775 10194 10784
rect 10140 10532 10192 10538
rect 10140 10474 10192 10480
rect 10152 9722 10180 10474
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10152 8498 10180 8910
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10060 8350 10180 8378
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9968 8090 9996 8230
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9784 6446 9904 6474
rect 9588 5102 9640 5108
rect 9678 5128 9734 5137
rect 9404 5092 9456 5098
rect 9678 5063 9734 5072
rect 9404 5034 9456 5040
rect 9416 3380 9444 5034
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9692 3738 9720 4626
rect 9784 3738 9812 6446
rect 9862 5128 9918 5137
rect 9862 5063 9918 5072
rect 9876 4214 9904 5063
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9876 3618 9904 3878
rect 9968 3670 9996 7890
rect 10060 5030 10088 8026
rect 10152 5166 10180 8350
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10152 4729 10180 4762
rect 10138 4720 10194 4729
rect 10138 4655 10194 4664
rect 10244 4536 10272 12600
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10336 10690 10364 12378
rect 10414 12336 10470 12345
rect 10414 12271 10470 12280
rect 10428 10810 10456 12271
rect 10520 11762 10548 12786
rect 10612 12442 10640 13262
rect 10796 12968 10824 16918
rect 10980 15994 11008 19926
rect 11058 19816 11114 19825
rect 11058 19751 11114 19760
rect 11072 19009 11100 19751
rect 11058 19000 11114 19009
rect 11058 18935 11114 18944
rect 11164 18850 11192 22320
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11624 19514 11652 22320
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11992 19394 12020 22320
rect 12254 19952 12310 19961
rect 12254 19887 12310 19896
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 11072 18822 11192 18850
rect 11624 19366 12020 19394
rect 12084 19378 12112 19790
rect 12072 19372 12124 19378
rect 11072 16794 11100 18822
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 11164 17746 11192 18702
rect 11624 18630 11652 19366
rect 12072 19314 12124 19320
rect 11888 19236 11940 19242
rect 11888 19178 11940 19184
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11716 18630 11744 19110
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11808 17921 11836 19110
rect 11900 18358 11928 19178
rect 12084 18834 12112 19314
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 12176 18970 12204 19110
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12084 18426 12112 18770
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 11888 18352 11940 18358
rect 11888 18294 11940 18300
rect 12268 18290 12296 19887
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 11978 18184 12034 18193
rect 11888 18148 11940 18154
rect 11978 18119 11980 18128
rect 11888 18090 11940 18096
rect 12032 18119 12034 18128
rect 12162 18184 12218 18193
rect 12162 18119 12218 18128
rect 11980 18090 12032 18096
rect 11794 17912 11850 17921
rect 11794 17847 11850 17856
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 11796 17604 11848 17610
rect 11796 17546 11848 17552
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11164 17202 11192 17478
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11152 17196 11204 17202
rect 11152 17138 11204 17144
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 10888 15966 11008 15994
rect 10888 14822 10916 15966
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10888 13938 10916 14350
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10876 13456 10928 13462
rect 10876 13398 10928 13404
rect 10704 12940 10824 12968
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10598 11792 10654 11801
rect 10508 11756 10560 11762
rect 10598 11727 10654 11736
rect 10508 11698 10560 11704
rect 10612 11529 10640 11727
rect 10704 11694 10732 12940
rect 10782 12880 10838 12889
rect 10782 12815 10838 12824
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10796 11626 10824 12815
rect 10888 12714 10916 13398
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10888 12617 10916 12650
rect 10874 12608 10930 12617
rect 10874 12543 10930 12552
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10888 11642 10916 12378
rect 10980 12209 11008 15846
rect 11164 15745 11192 17002
rect 11808 16658 11836 17546
rect 11900 17134 11928 18090
rect 11980 17808 12032 17814
rect 12176 17785 12204 18119
rect 12360 17882 12388 22320
rect 12728 20074 12756 22320
rect 12544 20046 12756 20074
rect 12438 19544 12494 19553
rect 12438 19479 12440 19488
rect 12492 19479 12494 19488
rect 12440 19450 12492 19456
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12256 17808 12308 17814
rect 11980 17750 12032 17756
rect 12162 17776 12218 17785
rect 11888 17128 11940 17134
rect 11992 17105 12020 17750
rect 12256 17750 12308 17756
rect 12162 17711 12218 17720
rect 12164 17672 12216 17678
rect 12070 17640 12126 17649
rect 12164 17614 12216 17620
rect 12070 17575 12126 17584
rect 11888 17070 11940 17076
rect 11978 17096 12034 17105
rect 11900 16794 11928 17070
rect 11978 17031 12034 17040
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11992 16658 12020 16934
rect 12084 16697 12112 17575
rect 12070 16688 12126 16697
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11980 16652 12032 16658
rect 12070 16623 12126 16632
rect 11980 16594 12032 16600
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11612 15972 11664 15978
rect 11612 15914 11664 15920
rect 11150 15736 11206 15745
rect 11150 15671 11206 15680
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11624 15162 11652 15914
rect 11808 15910 11836 16594
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 12084 15638 12112 16526
rect 12072 15632 12124 15638
rect 12072 15574 12124 15580
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11518 15056 11574 15065
rect 11518 14991 11574 15000
rect 11428 14884 11480 14890
rect 11428 14826 11480 14832
rect 11440 14521 11468 14826
rect 11426 14512 11482 14521
rect 11060 14476 11112 14482
rect 11426 14447 11482 14456
rect 11060 14418 11112 14424
rect 11072 13530 11100 14418
rect 11532 14414 11560 14991
rect 11624 14482 11652 15098
rect 12084 14804 12112 15574
rect 12176 15026 12204 17614
rect 12268 15366 12296 17750
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12256 15360 12308 15366
rect 12254 15328 12256 15337
rect 12308 15328 12310 15337
rect 12254 15263 12310 15272
rect 12268 15237 12296 15263
rect 12360 15178 12388 17614
rect 12452 17338 12480 19246
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12544 17270 12572 20046
rect 12992 19984 13044 19990
rect 12992 19926 13044 19932
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 12636 18426 12664 19858
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12716 18896 12768 18902
rect 12716 18838 12768 18844
rect 12728 18426 12756 18838
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12532 17264 12584 17270
rect 12532 17206 12584 17212
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12636 17105 12664 17206
rect 12622 17096 12678 17105
rect 12532 17060 12584 17066
rect 12622 17031 12678 17040
rect 12532 17002 12584 17008
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12452 16153 12480 16594
rect 12544 16454 12572 17002
rect 12728 16980 12756 18158
rect 12820 18086 12848 19654
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12636 16952 12756 16980
rect 12808 16992 12860 16998
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12438 16144 12494 16153
rect 12438 16079 12494 16088
rect 12452 15745 12480 16079
rect 12438 15736 12494 15745
rect 12438 15671 12494 15680
rect 12268 15150 12388 15178
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12164 14816 12216 14822
rect 12084 14776 12164 14804
rect 12164 14758 12216 14764
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11978 14512 12034 14521
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11520 14408 11572 14414
rect 11518 14376 11520 14385
rect 11572 14376 11574 14385
rect 11518 14311 11574 14320
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11072 12850 11100 13126
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 11164 12782 11192 14214
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11426 13968 11482 13977
rect 11426 13903 11482 13912
rect 11440 13734 11468 13903
rect 11428 13728 11480 13734
rect 11428 13670 11480 13676
rect 11440 13394 11468 13670
rect 11518 13560 11574 13569
rect 11518 13495 11520 13504
rect 11572 13495 11574 13504
rect 11520 13466 11572 13472
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11624 12986 11652 14214
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11716 13462 11744 13670
rect 11704 13456 11756 13462
rect 11704 13398 11756 13404
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11150 12472 11206 12481
rect 11150 12407 11206 12416
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10966 12200 11022 12209
rect 10966 12135 11022 12144
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10980 11762 11008 12038
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10784 11620 10836 11626
rect 10888 11614 11008 11642
rect 10784 11562 10836 11568
rect 10598 11520 10654 11529
rect 10598 11455 10654 11464
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10336 10662 10456 10690
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10336 8022 10364 9998
rect 10428 9489 10456 10662
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10520 10130 10548 10202
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10612 10062 10640 11455
rect 10690 10976 10746 10985
rect 10690 10911 10746 10920
rect 10704 10810 10732 10911
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10704 10266 10732 10406
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10600 10056 10652 10062
rect 10652 10016 10732 10044
rect 10600 9998 10652 10004
rect 10508 9988 10560 9994
rect 10508 9930 10560 9936
rect 10520 9761 10548 9930
rect 10598 9888 10654 9897
rect 10598 9823 10654 9832
rect 10506 9752 10562 9761
rect 10506 9687 10562 9696
rect 10414 9480 10470 9489
rect 10414 9415 10470 9424
rect 10416 9376 10468 9382
rect 10520 9353 10548 9687
rect 10612 9518 10640 9823
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10600 9376 10652 9382
rect 10416 9318 10468 9324
rect 10506 9344 10562 9353
rect 10428 9178 10456 9318
rect 10600 9318 10652 9324
rect 10506 9279 10562 9288
rect 10612 9217 10640 9318
rect 10598 9208 10654 9217
rect 10416 9172 10468 9178
rect 10704 9178 10732 10016
rect 10598 9143 10654 9152
rect 10692 9172 10744 9178
rect 10416 9114 10468 9120
rect 10692 9114 10744 9120
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10324 8016 10376 8022
rect 10324 7958 10376 7964
rect 10612 7954 10640 8978
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10704 8265 10732 8298
rect 10690 8256 10746 8265
rect 10690 8191 10746 8200
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10416 7812 10468 7818
rect 10416 7754 10468 7760
rect 10322 7576 10378 7585
rect 10322 7511 10378 7520
rect 10060 4508 10272 4536
rect 9692 3590 9904 3618
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9416 3352 9536 3380
rect 9310 3224 9366 3233
rect 9310 3159 9366 3168
rect 9126 2816 9182 2825
rect 9126 2751 9182 2760
rect 9140 2514 9168 2751
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 9312 2304 9364 2310
rect 9126 2272 9182 2281
rect 9312 2246 9364 2252
rect 9126 2207 9182 2216
rect 9036 1964 9088 1970
rect 9036 1906 9088 1912
rect 8772 1278 8984 1306
rect 8772 480 8800 1278
rect 9140 480 9168 2207
rect 9324 1970 9352 2246
rect 9312 1964 9364 1970
rect 9312 1906 9364 1912
rect 9508 480 9536 3352
rect 9692 1426 9720 3590
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9784 2825 9812 3470
rect 9968 3126 9996 3470
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 10060 2972 10088 4508
rect 10336 4434 10364 7511
rect 10428 7410 10456 7754
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10520 7274 10548 7822
rect 10796 7392 10824 11562
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10612 7364 10824 7392
rect 10508 7268 10560 7274
rect 10508 7210 10560 7216
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10428 6916 10456 7142
rect 10428 6888 10548 6916
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10428 5574 10456 6734
rect 10520 6089 10548 6888
rect 10506 6080 10562 6089
rect 10506 6015 10562 6024
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10428 4758 10456 4966
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 9876 2944 10088 2972
rect 10152 4406 10364 4434
rect 9770 2816 9826 2825
rect 9770 2751 9826 2760
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9784 1834 9812 2246
rect 9772 1828 9824 1834
rect 9772 1770 9824 1776
rect 9680 1420 9732 1426
rect 9680 1362 9732 1368
rect 9876 480 9904 2944
rect 10152 2514 10180 4406
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10336 3942 10364 4150
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10244 3534 10272 3878
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10244 3058 10272 3470
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10336 2990 10364 3878
rect 10324 2984 10376 2990
rect 10230 2952 10286 2961
rect 10324 2926 10376 2932
rect 10230 2887 10286 2896
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 9968 2106 9996 2450
rect 9956 2100 10008 2106
rect 9956 2042 10008 2048
rect 10152 1834 10180 2450
rect 10140 1828 10192 1834
rect 10140 1770 10192 1776
rect 10244 480 10272 2887
rect 10322 2680 10378 2689
rect 10322 2615 10324 2624
rect 10376 2615 10378 2624
rect 10324 2586 10376 2592
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 10336 1902 10364 2450
rect 10428 2446 10456 4694
rect 10612 4196 10640 7364
rect 10888 7290 10916 11494
rect 10980 7585 11008 11614
rect 11072 10810 11100 12242
rect 11164 11694 11192 12407
rect 11716 12073 11744 13262
rect 11702 12064 11758 12073
rect 11252 11996 11548 12016
rect 11702 11999 11758 12008
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11808 11914 11836 13330
rect 11900 12850 11928 14486
rect 11978 14447 12034 14456
rect 11992 12918 12020 14447
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12084 13530 12112 13806
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11886 12608 11942 12617
rect 11886 12543 11942 12552
rect 11900 12345 11928 12543
rect 12084 12481 12112 12922
rect 12176 12782 12204 14758
rect 12268 14385 12296 15150
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12254 14376 12310 14385
rect 12254 14311 12310 14320
rect 12268 13802 12296 14311
rect 12256 13796 12308 13802
rect 12256 13738 12308 13744
rect 12254 13696 12310 13705
rect 12254 13631 12310 13640
rect 12268 12986 12296 13631
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 12070 12472 12126 12481
rect 11980 12436 12032 12442
rect 12070 12407 12126 12416
rect 11980 12378 12032 12384
rect 11886 12336 11942 12345
rect 11886 12271 11942 12280
rect 11992 12209 12020 12378
rect 12070 12336 12126 12345
rect 12070 12271 12126 12280
rect 12254 12336 12310 12345
rect 12254 12271 12310 12280
rect 11978 12200 12034 12209
rect 11978 12135 12034 12144
rect 11624 11886 11836 11914
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11072 10266 11100 10746
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11164 10146 11192 11086
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11072 10130 11192 10146
rect 11060 10124 11192 10130
rect 11112 10118 11192 10124
rect 11060 10066 11112 10072
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 11072 9450 11100 9930
rect 11348 9908 11376 10474
rect 11624 9994 11652 11886
rect 11980 11824 12032 11830
rect 11794 11792 11850 11801
rect 11704 11756 11756 11762
rect 11980 11766 12032 11772
rect 11794 11727 11850 11736
rect 11888 11756 11940 11762
rect 11704 11698 11756 11704
rect 11716 10062 11744 11698
rect 11808 11558 11836 11727
rect 11888 11698 11940 11704
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11808 10130 11836 11154
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11808 9908 11836 10066
rect 11164 9880 11376 9908
rect 11716 9880 11836 9908
rect 11164 9704 11192 9880
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11164 9676 11376 9704
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 11164 9330 11192 9522
rect 11072 9302 11192 9330
rect 11072 8498 11100 9302
rect 11150 9208 11206 9217
rect 11150 9143 11206 9152
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11164 8401 11192 9143
rect 11348 8945 11376 9676
rect 11518 9616 11574 9625
rect 11518 9551 11574 9560
rect 11532 8945 11560 9551
rect 11610 9344 11666 9353
rect 11610 9279 11666 9288
rect 11334 8936 11390 8945
rect 11334 8871 11390 8880
rect 11518 8936 11574 8945
rect 11518 8871 11574 8880
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11150 8392 11206 8401
rect 11150 8327 11206 8336
rect 11058 8120 11114 8129
rect 11058 8055 11114 8064
rect 10966 7576 11022 7585
rect 10966 7511 11022 7520
rect 11072 7449 11100 8055
rect 11242 7848 11298 7857
rect 11164 7806 11242 7834
rect 11058 7440 11114 7449
rect 10968 7404 11020 7410
rect 11058 7375 11114 7384
rect 10968 7346 11020 7352
rect 10796 7262 10916 7290
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10704 5642 10732 6598
rect 10796 6089 10824 7262
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10888 7002 10916 7142
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10980 6100 11008 7346
rect 11164 7313 11192 7806
rect 11242 7783 11298 7792
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11624 7546 11652 9279
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11150 7304 11206 7313
rect 11060 7268 11112 7274
rect 11518 7304 11574 7313
rect 11150 7239 11206 7248
rect 11428 7268 11480 7274
rect 11060 7210 11112 7216
rect 11518 7239 11574 7248
rect 11428 7210 11480 7216
rect 11072 6730 11100 7210
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11256 6905 11284 6938
rect 11242 6896 11298 6905
rect 11242 6831 11298 6840
rect 11440 6798 11468 7210
rect 11532 6934 11560 7239
rect 11520 6928 11572 6934
rect 11520 6870 11572 6876
rect 11624 6866 11652 7346
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 11612 6656 11664 6662
rect 11058 6624 11114 6633
rect 11612 6598 11664 6604
rect 11058 6559 11114 6568
rect 11072 6390 11100 6559
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11060 6112 11112 6118
rect 10782 6080 10838 6089
rect 10980 6072 11060 6100
rect 11060 6054 11112 6060
rect 10782 6015 10838 6024
rect 11072 5846 11100 6054
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11624 5778 11652 6598
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 10692 5636 10744 5642
rect 10692 5578 10744 5584
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10704 5001 10732 5306
rect 10966 5128 11022 5137
rect 10966 5063 11022 5072
rect 10784 5024 10836 5030
rect 10690 4992 10746 5001
rect 10784 4966 10836 4972
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10690 4927 10746 4936
rect 10520 4168 10640 4196
rect 10520 3346 10548 4168
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10612 3466 10640 3946
rect 10704 3738 10732 4014
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10600 3460 10652 3466
rect 10600 3402 10652 3408
rect 10704 3369 10732 3470
rect 10690 3360 10746 3369
rect 10520 3318 10640 3346
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10520 2650 10548 3062
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10324 1896 10376 1902
rect 10324 1838 10376 1844
rect 10612 480 10640 3318
rect 10690 3295 10746 3304
rect 10704 3058 10732 3295
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10796 1290 10824 4966
rect 10888 4826 10916 4966
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10980 4706 11008 5063
rect 11164 4826 11192 5510
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11716 5137 11744 9880
rect 11900 9722 11928 11698
rect 11992 9738 12020 11766
rect 12084 11218 12112 12271
rect 12162 12064 12218 12073
rect 12162 11999 12218 12008
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12070 10840 12126 10849
rect 12070 10775 12126 10784
rect 12084 10538 12112 10775
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 12176 10470 12204 11999
rect 12268 11898 12296 12271
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12254 11792 12310 11801
rect 12254 11727 12310 11736
rect 12268 11393 12296 11727
rect 12254 11384 12310 11393
rect 12254 11319 12310 11328
rect 12360 11268 12388 14962
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 14113 12480 14894
rect 12530 14240 12586 14249
rect 12530 14175 12586 14184
rect 12438 14104 12494 14113
rect 12438 14039 12494 14048
rect 12544 14006 12572 14175
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12452 12102 12480 12718
rect 12636 12458 12664 16952
rect 12808 16934 12860 16940
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 12728 16153 12756 16662
rect 12714 16144 12770 16153
rect 12714 16079 12770 16088
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12728 15026 12756 15846
rect 12820 15162 12848 16934
rect 12912 16250 12940 19654
rect 13004 16250 13032 19926
rect 13096 19242 13124 22320
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 13084 19236 13136 19242
rect 13084 19178 13136 19184
rect 13084 18896 13136 18902
rect 13084 18838 13136 18844
rect 13096 18290 13124 18838
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 13096 17202 13124 18022
rect 13188 17814 13216 20198
rect 13464 19938 13492 22320
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13372 19910 13492 19938
rect 13268 18420 13320 18426
rect 13268 18362 13320 18368
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13280 17252 13308 18362
rect 13372 17882 13400 19910
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13464 19310 13492 19790
rect 13740 19786 13768 20198
rect 13728 19780 13780 19786
rect 13728 19722 13780 19728
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13452 19304 13504 19310
rect 13452 19246 13504 19252
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 13280 17224 13400 17252
rect 13084 17196 13136 17202
rect 13136 17156 13308 17184
rect 13084 17138 13136 17144
rect 13174 17096 13230 17105
rect 13174 17031 13230 17040
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 13096 16794 13124 16934
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 13084 16652 13136 16658
rect 13188 16640 13216 17031
rect 13136 16612 13216 16640
rect 13084 16594 13136 16600
rect 12900 16244 12952 16250
rect 12900 16186 12952 16192
rect 12992 16244 13044 16250
rect 12992 16186 13044 16192
rect 13280 16114 13308 17156
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13268 15972 13320 15978
rect 13268 15914 13320 15920
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12716 14544 12768 14550
rect 12716 14486 12768 14492
rect 12728 14074 12756 14486
rect 12820 14074 12848 14758
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12714 13016 12770 13025
rect 12714 12951 12770 12960
rect 12728 12918 12756 12951
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12636 12430 12848 12458
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12452 11762 12480 12038
rect 12530 11792 12586 11801
rect 12440 11756 12492 11762
rect 12530 11727 12586 11736
rect 12440 11698 12492 11704
rect 12268 11240 12388 11268
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 12072 9920 12124 9926
rect 12070 9888 12072 9897
rect 12124 9888 12126 9897
rect 12070 9823 12126 9832
rect 11888 9716 11940 9722
rect 11992 9710 12112 9738
rect 11888 9658 11940 9664
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11808 8945 11836 9114
rect 11794 8936 11850 8945
rect 11794 8871 11850 8880
rect 11794 8800 11850 8809
rect 11794 8735 11850 8744
rect 11808 8430 11836 8735
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11702 5128 11758 5137
rect 11612 5092 11664 5098
rect 11702 5063 11758 5072
rect 11612 5034 11664 5040
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11440 4826 11468 4966
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 10888 4690 11008 4706
rect 10876 4684 11008 4690
rect 10928 4678 11008 4684
rect 10876 4626 10928 4632
rect 10888 2666 10916 4626
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10980 3505 11008 4422
rect 11072 3670 11100 4558
rect 11440 4554 11468 4762
rect 11428 4548 11480 4554
rect 11428 4490 11480 4496
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11624 3992 11652 5034
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11716 4146 11744 4422
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11808 4060 11836 8366
rect 11900 6866 11928 9658
rect 11980 9648 12032 9654
rect 11978 9616 11980 9625
rect 12032 9616 12034 9625
rect 11978 9551 12034 9560
rect 11980 9444 12032 9450
rect 11980 9386 12032 9392
rect 11992 8673 12020 9386
rect 11978 8664 12034 8673
rect 11978 8599 12034 8608
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 11992 8401 12020 8502
rect 11978 8392 12034 8401
rect 11978 8327 12034 8336
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11992 7954 12020 8230
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 12084 7834 12112 9710
rect 12176 9450 12204 9930
rect 12268 9761 12296 11240
rect 12452 11218 12480 11698
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12544 11098 12572 11727
rect 12636 11676 12664 12038
rect 12728 11898 12756 12242
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12716 11688 12768 11694
rect 12636 11648 12716 11676
rect 12716 11630 12768 11636
rect 12622 11384 12678 11393
rect 12820 11354 12848 12430
rect 12622 11319 12624 11328
rect 12676 11319 12678 11328
rect 12808 11348 12860 11354
rect 12624 11290 12676 11296
rect 12808 11290 12860 11296
rect 12912 11234 12940 15846
rect 13084 14952 13136 14958
rect 13004 14912 13084 14940
rect 13004 14260 13032 14912
rect 13084 14894 13136 14900
rect 13082 14512 13138 14521
rect 13082 14447 13138 14456
rect 13096 14414 13124 14447
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13004 14232 13124 14260
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 13004 12442 13032 13262
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12990 12336 13046 12345
rect 12990 12271 13046 12280
rect 13004 12102 13032 12271
rect 13096 12170 13124 14232
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13188 13433 13216 14010
rect 13174 13424 13230 13433
rect 13174 13359 13230 13368
rect 13084 12164 13136 12170
rect 13084 12106 13136 12112
rect 12992 12096 13044 12102
rect 13188 12050 13216 13359
rect 13280 12646 13308 15914
rect 13372 14346 13400 17224
rect 13464 14804 13492 17682
rect 13556 15745 13584 18838
rect 13636 18828 13688 18834
rect 13636 18770 13688 18776
rect 13648 17134 13676 18770
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 13648 16454 13676 17070
rect 13740 16794 13768 19314
rect 13832 19174 13860 22320
rect 14200 19938 14228 22320
rect 14464 20732 14516 20738
rect 14464 20674 14516 20680
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14384 20058 14412 20334
rect 14372 20052 14424 20058
rect 14372 19994 14424 20000
rect 13924 19910 14228 19938
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13832 17066 13860 18770
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13542 15736 13598 15745
rect 13542 15671 13598 15680
rect 13544 15632 13596 15638
rect 13544 15574 13596 15580
rect 13556 14906 13584 15574
rect 13636 15564 13688 15570
rect 13740 15552 13768 16730
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13832 15706 13860 15846
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13688 15524 13860 15552
rect 13636 15506 13688 15512
rect 13728 14952 13780 14958
rect 13556 14878 13676 14906
rect 13728 14894 13780 14900
rect 13464 14776 13584 14804
rect 13556 14346 13584 14776
rect 13360 14340 13412 14346
rect 13360 14282 13412 14288
rect 13544 14340 13596 14346
rect 13544 14282 13596 14288
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13358 13424 13414 13433
rect 13358 13359 13414 13368
rect 13372 12889 13400 13359
rect 13358 12880 13414 12889
rect 13358 12815 13414 12824
rect 13464 12782 13492 14214
rect 13544 13796 13596 13802
rect 13544 13738 13596 13744
rect 13556 13326 13584 13738
rect 13648 13394 13676 14878
rect 13740 14074 13768 14894
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13726 13152 13782 13161
rect 13726 13087 13782 13096
rect 13634 12880 13690 12889
rect 13634 12815 13690 12824
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 13544 12708 13596 12714
rect 13544 12650 13596 12656
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 12992 12038 13044 12044
rect 13096 12022 13216 12050
rect 12990 11928 13046 11937
rect 12990 11863 13046 11872
rect 13004 11694 13032 11863
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 12360 11070 12572 11098
rect 12728 11206 12940 11234
rect 12254 9752 12310 9761
rect 12254 9687 12310 9696
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12176 8956 12204 9386
rect 12268 9092 12296 9522
rect 12360 9518 12388 11070
rect 12438 10840 12494 10849
rect 12438 10775 12494 10784
rect 12452 10742 12480 10775
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12452 9178 12480 9862
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12348 9104 12400 9110
rect 12268 9064 12348 9092
rect 12400 9052 12480 9058
rect 12348 9046 12480 9052
rect 12360 9030 12480 9046
rect 12176 8928 12388 8956
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12176 8022 12204 8774
rect 12254 8664 12310 8673
rect 12254 8599 12310 8608
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 12268 7936 12296 8599
rect 12360 8090 12388 8928
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12452 7954 12480 9030
rect 12544 8634 12572 10134
rect 12636 8945 12664 10202
rect 12622 8936 12678 8945
rect 12622 8871 12678 8880
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12636 8514 12664 8774
rect 12544 8486 12664 8514
rect 12440 7948 12492 7954
rect 12268 7908 12388 7936
rect 12084 7806 12296 7834
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11992 6798 12020 7686
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12084 7313 12112 7346
rect 12070 7304 12126 7313
rect 12070 7239 12126 7248
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12176 7002 12204 7142
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12072 6928 12124 6934
rect 12072 6870 12124 6876
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11886 6488 11942 6497
rect 11886 6423 11942 6432
rect 11900 6390 11928 6423
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11888 6180 11940 6186
rect 11888 6122 11940 6128
rect 11900 4214 11928 6122
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 11888 4072 11940 4078
rect 11808 4032 11888 4060
rect 11992 4049 12020 6258
rect 12084 4826 12112 6870
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12176 5574 12204 5646
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12176 5234 12204 5510
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 11888 4014 11940 4020
rect 11978 4040 12034 4049
rect 11624 3964 11744 3992
rect 11978 3975 12034 3984
rect 11520 3936 11572 3942
rect 11572 3896 11652 3924
rect 11520 3878 11572 3884
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 11244 3664 11296 3670
rect 11244 3606 11296 3612
rect 11256 3516 11284 3606
rect 10966 3496 11022 3505
rect 10966 3431 11022 3440
rect 11072 3488 11284 3516
rect 11072 3369 11100 3488
rect 11058 3360 11114 3369
rect 11058 3295 11114 3304
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 10888 2638 11100 2666
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 10888 2038 10916 2246
rect 10876 2032 10928 2038
rect 10876 1974 10928 1980
rect 11072 1902 11100 2638
rect 11060 1896 11112 1902
rect 11060 1838 11112 1844
rect 10968 1828 11020 1834
rect 10968 1770 11020 1776
rect 10784 1284 10836 1290
rect 10784 1226 10836 1232
rect 10980 480 11008 1770
rect 11164 1442 11192 2858
rect 11624 2514 11652 3896
rect 11612 2508 11664 2514
rect 11612 2450 11664 2456
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11716 1494 11744 3964
rect 11978 3632 12034 3641
rect 11978 3567 12034 3576
rect 11794 3224 11850 3233
rect 11794 3159 11850 3168
rect 11808 3058 11836 3159
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11992 2836 12020 3567
rect 12084 3126 12112 4082
rect 12176 3398 12204 4558
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 12176 2990 12204 3334
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 11794 2816 11850 2825
rect 11992 2808 12204 2836
rect 11794 2751 11850 2760
rect 11704 1488 11756 1494
rect 11164 1414 11376 1442
rect 11704 1430 11756 1436
rect 11348 480 11376 1414
rect 11808 480 11836 2751
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 11992 1834 12020 2382
rect 11980 1828 12032 1834
rect 11980 1770 12032 1776
rect 12176 480 12204 2808
rect 12268 2514 12296 7806
rect 12360 5914 12388 7908
rect 12440 7890 12492 7896
rect 12452 7410 12480 7890
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12452 6236 12480 7346
rect 12544 6866 12572 8486
rect 12728 7834 12756 11206
rect 13096 11132 13124 12022
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 12806 11112 12862 11121
rect 12806 11047 12862 11056
rect 12912 11104 13124 11132
rect 12820 11014 12848 11047
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12820 8566 12848 10406
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12806 8392 12862 8401
rect 12806 8327 12862 8336
rect 12636 7806 12756 7834
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12532 6248 12584 6254
rect 12452 6208 12532 6236
rect 12532 6190 12584 6196
rect 12438 6080 12494 6089
rect 12438 6015 12494 6024
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12452 5794 12480 6015
rect 12360 5778 12480 5794
rect 12348 5772 12480 5778
rect 12400 5766 12480 5772
rect 12544 5760 12572 6190
rect 12636 5953 12664 7806
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12622 5944 12678 5953
rect 12622 5879 12678 5888
rect 12624 5772 12676 5778
rect 12544 5732 12624 5760
rect 12348 5714 12400 5720
rect 12624 5714 12676 5720
rect 12438 5672 12494 5681
rect 12438 5607 12494 5616
rect 12624 5636 12676 5642
rect 12452 5370 12480 5607
rect 12624 5578 12676 5584
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12440 5024 12492 5030
rect 12346 4992 12402 5001
rect 12636 5001 12664 5578
rect 12440 4966 12492 4972
rect 12622 4992 12678 5001
rect 12346 4927 12402 4936
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 12360 2446 12388 4927
rect 12452 4826 12480 4966
rect 12622 4927 12678 4936
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12622 4040 12678 4049
rect 12622 3975 12624 3984
rect 12676 3975 12678 3984
rect 12624 3946 12676 3952
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12452 3738 12480 3878
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12530 3496 12586 3505
rect 12530 3431 12586 3440
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12452 2378 12480 3062
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 12544 480 12572 3431
rect 12728 3346 12756 7686
rect 12820 7002 12848 8327
rect 12912 7041 12940 11104
rect 12990 10976 13046 10985
rect 12990 10911 13046 10920
rect 13004 10062 13032 10911
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 13004 9704 13032 9998
rect 13084 9716 13136 9722
rect 13004 9676 13084 9704
rect 13004 9042 13032 9676
rect 13084 9658 13136 9664
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 12990 8800 13046 8809
rect 12990 8735 13046 8744
rect 13004 7313 13032 8735
rect 13096 8498 13124 9318
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 13082 7576 13138 7585
rect 13082 7511 13138 7520
rect 12990 7304 13046 7313
rect 12990 7239 13046 7248
rect 12898 7032 12954 7041
rect 12808 6996 12860 7002
rect 12898 6967 12954 6976
rect 12808 6938 12860 6944
rect 13096 6934 13124 7511
rect 13188 7002 13216 11290
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 12900 6928 12952 6934
rect 12898 6896 12900 6905
rect 13084 6928 13136 6934
rect 12952 6896 12954 6905
rect 13084 6870 13136 6876
rect 12898 6831 12954 6840
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12820 5914 12848 6054
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12912 4570 12940 6831
rect 13188 6798 13216 6938
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13280 6458 13308 12582
rect 13372 11937 13400 12650
rect 13556 12374 13584 12650
rect 13648 12646 13676 12815
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13544 12368 13596 12374
rect 13450 12336 13506 12345
rect 13544 12310 13596 12316
rect 13450 12271 13506 12280
rect 13358 11928 13414 11937
rect 13358 11863 13414 11872
rect 13372 6662 13400 11863
rect 13464 10810 13492 12271
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13556 11354 13584 12174
rect 13636 12164 13688 12170
rect 13636 12106 13688 12112
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13556 11257 13584 11290
rect 13542 11248 13598 11257
rect 13648 11218 13676 12106
rect 13740 11626 13768 13087
rect 13832 12850 13860 15524
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13832 12424 13860 12786
rect 13924 12714 13952 19910
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 14200 19417 14228 19790
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14186 19408 14242 19417
rect 14186 19343 14242 19352
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 14016 18193 14044 19246
rect 14292 18698 14320 19450
rect 14370 19136 14426 19145
rect 14370 19071 14426 19080
rect 14384 18970 14412 19071
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 14108 18426 14136 18566
rect 14096 18420 14148 18426
rect 14096 18362 14148 18368
rect 14200 18306 14228 18566
rect 14108 18290 14228 18306
rect 14108 18284 14240 18290
rect 14108 18278 14188 18284
rect 14002 18184 14058 18193
rect 14002 18119 14058 18128
rect 14108 17320 14136 18278
rect 14188 18226 14240 18232
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14200 18195 14228 18226
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14016 17292 14136 17320
rect 14016 17066 14044 17292
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 14016 16522 14044 17002
rect 14094 16960 14150 16969
rect 14094 16895 14150 16904
rect 14108 16590 14136 16895
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 14200 16538 14228 17614
rect 14292 16726 14320 18226
rect 14476 18170 14504 20674
rect 14660 20346 14688 22320
rect 14568 20318 14688 20346
rect 14568 18465 14596 20318
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 14554 18456 14610 18465
rect 14554 18391 14610 18400
rect 14556 18352 14608 18358
rect 14556 18294 14608 18300
rect 14384 18142 14504 18170
rect 14384 17678 14412 18142
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14280 16720 14332 16726
rect 14280 16662 14332 16668
rect 14004 16516 14056 16522
rect 14200 16510 14320 16538
rect 14004 16458 14056 16464
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 14094 15736 14150 15745
rect 14094 15671 14150 15680
rect 14108 15570 14136 15671
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 14094 15056 14150 15065
rect 14094 14991 14096 15000
rect 14148 14991 14150 15000
rect 14096 14962 14148 14968
rect 14200 13870 14228 16186
rect 14292 15502 14320 16510
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14096 13456 14148 13462
rect 14096 13398 14148 13404
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 14004 12708 14056 12714
rect 14004 12650 14056 12656
rect 13832 12396 13952 12424
rect 13924 12306 13952 12396
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13832 11506 13860 12242
rect 13912 11824 13964 11830
rect 13912 11766 13964 11772
rect 13740 11478 13860 11506
rect 13542 11183 13598 11192
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13648 10674 13676 11018
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13464 10130 13492 10542
rect 13542 10432 13598 10441
rect 13542 10367 13598 10376
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13556 10033 13584 10367
rect 13542 10024 13598 10033
rect 13542 9959 13598 9968
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13464 9217 13492 9862
rect 13450 9208 13506 9217
rect 13450 9143 13506 9152
rect 13452 8832 13504 8838
rect 13556 8820 13584 9862
rect 13648 9518 13676 10610
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13636 8832 13688 8838
rect 13556 8792 13636 8820
rect 13452 8774 13504 8780
rect 13636 8774 13688 8780
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13372 6338 13400 6394
rect 13188 6310 13400 6338
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 13004 5846 13032 6122
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 13082 5808 13138 5817
rect 13188 5778 13216 6310
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 13082 5743 13138 5752
rect 13176 5772 13228 5778
rect 13096 5642 13124 5743
rect 13176 5714 13228 5720
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 13004 5234 13032 5510
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13082 5128 13138 5137
rect 13082 5063 13138 5072
rect 13096 4865 13124 5063
rect 13082 4856 13138 4865
rect 13082 4791 13138 4800
rect 13096 4758 13124 4791
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 12912 4542 13032 4570
rect 12900 4480 12952 4486
rect 12806 4448 12862 4457
rect 12900 4422 12952 4428
rect 12806 4383 12862 4392
rect 12820 4078 12848 4383
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12820 3777 12848 3878
rect 12806 3768 12862 3777
rect 12806 3703 12862 3712
rect 12912 3670 12940 4422
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12636 3318 12756 3346
rect 12636 2530 12664 3318
rect 12820 3210 12848 3470
rect 12728 3182 12848 3210
rect 12728 2990 12756 3182
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 13004 2938 13032 4542
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13096 4214 13124 4422
rect 13084 4208 13136 4214
rect 13084 4150 13136 4156
rect 13188 4078 13216 5714
rect 13372 5545 13400 5782
rect 13358 5536 13414 5545
rect 13358 5471 13414 5480
rect 13266 5400 13322 5409
rect 13266 5335 13322 5344
rect 13280 5030 13308 5335
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13280 4593 13308 4966
rect 13266 4584 13322 4593
rect 13266 4519 13322 4528
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13082 3904 13138 3913
rect 13082 3839 13138 3848
rect 13096 3058 13124 3839
rect 13188 3602 13216 4014
rect 13372 4010 13400 5170
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 13266 3088 13322 3097
rect 13084 3052 13136 3058
rect 13266 3023 13322 3032
rect 13084 2994 13136 3000
rect 12820 2650 12848 2926
rect 13004 2910 13216 2938
rect 12990 2816 13046 2825
rect 12990 2751 13046 2760
rect 13004 2650 13032 2751
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 13082 2544 13138 2553
rect 12636 2502 12940 2530
rect 12912 480 12940 2502
rect 13082 2479 13138 2488
rect 13096 2446 13124 2479
rect 13188 2446 13216 2910
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13280 480 13308 3023
rect 13464 2990 13492 8774
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13556 6798 13584 8434
rect 13648 7154 13676 8570
rect 13740 8537 13768 11478
rect 13924 11150 13952 11766
rect 14016 11257 14044 12650
rect 14108 12442 14136 13398
rect 14200 12918 14228 13806
rect 14292 13394 14320 13874
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14188 12912 14240 12918
rect 14188 12854 14240 12860
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14186 12472 14242 12481
rect 14096 12436 14148 12442
rect 14186 12407 14242 12416
rect 14096 12378 14148 12384
rect 14200 12374 14228 12407
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14188 12164 14240 12170
rect 14188 12106 14240 12112
rect 14200 11762 14228 12106
rect 14292 11830 14320 12718
rect 14384 12238 14412 14010
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14280 11824 14332 11830
rect 14280 11766 14332 11772
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14188 11620 14240 11626
rect 14108 11580 14188 11608
rect 14108 11286 14136 11580
rect 14188 11562 14240 11568
rect 14186 11384 14242 11393
rect 14186 11319 14242 11328
rect 14096 11280 14148 11286
rect 14002 11248 14058 11257
rect 14096 11222 14148 11228
rect 14002 11183 14058 11192
rect 13912 11144 13964 11150
rect 13910 11112 13912 11121
rect 14004 11144 14056 11150
rect 13964 11112 13966 11121
rect 14004 11086 14056 11092
rect 13910 11047 13966 11056
rect 13924 11021 13952 11047
rect 14016 10985 14044 11086
rect 14096 11076 14148 11082
rect 14096 11018 14148 11024
rect 14002 10976 14058 10985
rect 14002 10911 14058 10920
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13820 10600 13872 10606
rect 13872 10560 13952 10588
rect 13820 10542 13872 10548
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13726 8528 13782 8537
rect 13726 8463 13782 8472
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13740 7721 13768 8366
rect 13832 8090 13860 10406
rect 13924 9489 13952 10560
rect 13910 9480 13966 9489
rect 13910 9415 13966 9424
rect 14016 9058 14044 10610
rect 14108 9178 14136 11018
rect 14200 10985 14228 11319
rect 14186 10976 14242 10985
rect 14186 10911 14242 10920
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14200 10062 14228 10746
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14200 9586 14228 9998
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14016 9030 14136 9058
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 13912 8900 13964 8906
rect 13912 8842 13964 8848
rect 13924 8634 13952 8842
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13924 8129 13952 8366
rect 13910 8120 13966 8129
rect 13820 8084 13872 8090
rect 13910 8055 13966 8064
rect 13820 8026 13872 8032
rect 13726 7712 13782 7721
rect 13726 7647 13782 7656
rect 13728 7472 13780 7478
rect 13728 7414 13780 7420
rect 13740 7290 13768 7414
rect 13740 7262 13860 7290
rect 13648 7126 13768 7154
rect 13634 7032 13690 7041
rect 13634 6967 13690 6976
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 13556 1766 13584 6598
rect 13648 4457 13676 6967
rect 13740 5658 13768 7126
rect 13832 6254 13860 7262
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 13924 6390 13952 6802
rect 14016 6458 14044 8910
rect 14108 8498 14136 9030
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14108 7954 14136 8434
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14200 7750 14228 9522
rect 14292 9518 14320 11766
rect 14384 11393 14412 12174
rect 14370 11384 14426 11393
rect 14370 11319 14426 11328
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14384 10470 14412 11154
rect 14372 10464 14424 10470
rect 14476 10441 14504 18022
rect 14568 17882 14596 18294
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14844 17338 14872 17614
rect 15028 17513 15056 22320
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 15120 17785 15148 19790
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 15212 18290 15240 19654
rect 15396 18873 15424 22320
rect 15474 19408 15530 19417
rect 15474 19343 15530 19352
rect 15488 18902 15516 19343
rect 15476 18896 15528 18902
rect 15382 18864 15438 18873
rect 15292 18828 15344 18834
rect 15476 18838 15528 18844
rect 15382 18799 15438 18808
rect 15292 18770 15344 18776
rect 15304 18465 15332 18770
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15290 18456 15346 18465
rect 15290 18391 15346 18400
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 15384 18148 15436 18154
rect 15384 18090 15436 18096
rect 15198 17912 15254 17921
rect 15198 17847 15254 17856
rect 15212 17814 15240 17847
rect 15200 17808 15252 17814
rect 15106 17776 15162 17785
rect 15200 17750 15252 17756
rect 15106 17711 15162 17720
rect 15014 17504 15070 17513
rect 15014 17439 15070 17448
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 14554 16688 14610 16697
rect 14554 16623 14610 16632
rect 14568 13462 14596 16623
rect 15120 16250 15148 17711
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15200 17060 15252 17066
rect 15200 17002 15252 17008
rect 15212 16658 15240 17002
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15198 16416 15254 16425
rect 15198 16351 15254 16360
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15108 16108 15160 16114
rect 15212 16096 15240 16351
rect 15160 16068 15240 16096
rect 15108 16050 15160 16056
rect 15120 15881 15148 16050
rect 15106 15872 15162 15881
rect 14684 15804 14980 15824
rect 15106 15807 15162 15816
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 15106 15736 15162 15745
rect 15106 15671 15162 15680
rect 15014 15600 15070 15609
rect 15014 15535 15070 15544
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14660 14890 14688 15302
rect 15028 15162 15056 15535
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 15014 15056 15070 15065
rect 15014 14991 15070 15000
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14646 14512 14702 14521
rect 14646 14447 14702 14456
rect 14660 13870 14688 14447
rect 14924 14340 14976 14346
rect 14924 14282 14976 14288
rect 14648 13864 14700 13870
rect 14646 13832 14648 13841
rect 14700 13832 14702 13841
rect 14646 13767 14702 13776
rect 14936 13716 14964 14282
rect 15028 13870 15056 14991
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14936 13688 15056 13716
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14556 13456 14608 13462
rect 14556 13398 14608 13404
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14660 13161 14688 13330
rect 14646 13152 14702 13161
rect 14646 13087 14702 13096
rect 14830 13152 14886 13161
rect 14830 13087 14886 13096
rect 14844 12986 14872 13087
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 14554 12744 14610 12753
rect 14936 12714 14964 12922
rect 14554 12679 14610 12688
rect 14924 12708 14976 12714
rect 14568 12646 14596 12679
rect 14924 12650 14976 12656
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14752 12294 14964 12322
rect 14554 12200 14610 12209
rect 14554 12135 14610 12144
rect 14568 11121 14596 12135
rect 14648 11620 14700 11626
rect 14752 11608 14780 12294
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14844 11626 14872 12174
rect 14936 12170 14964 12294
rect 14924 12164 14976 12170
rect 14924 12106 14976 12112
rect 14700 11580 14780 11608
rect 14832 11620 14884 11626
rect 14648 11562 14700 11568
rect 14832 11562 14884 11568
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 14740 11280 14792 11286
rect 14740 11222 14792 11228
rect 14554 11112 14610 11121
rect 14554 11047 14610 11056
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14372 10406 14424 10412
rect 14462 10432 14518 10441
rect 14462 10367 14518 10376
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14476 9926 14504 10202
rect 14568 10130 14596 10950
rect 14752 10520 14780 11222
rect 14832 10532 14884 10538
rect 14752 10492 14832 10520
rect 14832 10474 14884 10480
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14936 9625 14964 9998
rect 14922 9616 14978 9625
rect 14922 9551 14978 9560
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14370 9208 14426 9217
rect 14370 9143 14426 9152
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14292 8498 14320 8910
rect 14384 8498 14412 9143
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14476 8566 14504 8978
rect 14464 8560 14516 8566
rect 14464 8502 14516 8508
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14464 8288 14516 8294
rect 14278 8256 14334 8265
rect 14464 8230 14516 8236
rect 14278 8191 14334 8200
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14094 7576 14150 7585
rect 14094 7511 14150 7520
rect 14108 7478 14136 7511
rect 14096 7472 14148 7478
rect 14096 7414 14148 7420
rect 14200 7274 14228 7686
rect 14188 7268 14240 7274
rect 14188 7210 14240 7216
rect 14188 6928 14240 6934
rect 14188 6870 14240 6876
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13910 6080 13966 6089
rect 13910 6015 13966 6024
rect 13740 5630 13860 5658
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13634 4448 13690 4457
rect 13634 4383 13690 4392
rect 13740 4282 13768 5510
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13832 4049 13860 5630
rect 13924 5409 13952 6015
rect 14016 5545 14044 6394
rect 14108 6361 14136 6734
rect 14094 6352 14150 6361
rect 14094 6287 14150 6296
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 14108 5914 14136 6054
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14200 5778 14228 6870
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14002 5536 14058 5545
rect 14002 5471 14058 5480
rect 13910 5400 13966 5409
rect 13910 5335 13966 5344
rect 14200 5030 14228 5714
rect 13912 5024 13964 5030
rect 14096 5024 14148 5030
rect 13912 4966 13964 4972
rect 14094 4992 14096 5001
rect 14188 5024 14240 5030
rect 14148 4992 14150 5001
rect 13924 4826 13952 4966
rect 14188 4966 14240 4972
rect 14094 4927 14150 4936
rect 14094 4856 14150 4865
rect 13912 4820 13964 4826
rect 14094 4791 14150 4800
rect 13912 4762 13964 4768
rect 13910 4176 13966 4185
rect 13910 4111 13966 4120
rect 13818 4040 13874 4049
rect 13818 3975 13874 3984
rect 13818 3768 13874 3777
rect 13818 3703 13874 3712
rect 13634 2000 13690 2009
rect 13634 1935 13690 1944
rect 13544 1760 13596 1766
rect 13544 1702 13596 1708
rect 13648 480 13676 1935
rect 13832 1630 13860 3703
rect 13924 3534 13952 4111
rect 14108 4010 14136 4791
rect 14292 4690 14320 8191
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14384 7410 14412 8026
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14372 7268 14424 7274
rect 14476 7256 14504 8230
rect 14568 8004 14596 9318
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 15028 9042 15056 13688
rect 15120 13138 15148 15671
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 15212 14521 15240 15506
rect 15198 14512 15254 14521
rect 15198 14447 15254 14456
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15212 13977 15240 14350
rect 15198 13968 15254 13977
rect 15198 13903 15254 13912
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 15212 13326 15240 13738
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15120 13110 15240 13138
rect 15212 12918 15240 13110
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15198 12200 15254 12209
rect 15108 12164 15160 12170
rect 15198 12135 15254 12144
rect 15108 12106 15160 12112
rect 15120 11558 15148 12106
rect 15108 11552 15160 11558
rect 15106 11520 15108 11529
rect 15160 11520 15162 11529
rect 15106 11455 15162 11464
rect 15212 11014 15240 12135
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15120 9722 15148 10406
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 15212 9330 15240 10610
rect 15304 9586 15332 17614
rect 15396 17610 15424 18090
rect 15384 17604 15436 17610
rect 15384 17546 15436 17552
rect 15488 17218 15516 18702
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15396 17202 15516 17218
rect 15384 17196 15516 17202
rect 15436 17190 15516 17196
rect 15384 17138 15436 17144
rect 15396 15065 15424 17138
rect 15580 16794 15608 17682
rect 15672 17338 15700 17818
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15488 16114 15516 16594
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15488 15434 15516 16050
rect 15568 15496 15620 15502
rect 15566 15464 15568 15473
rect 15620 15464 15622 15473
rect 15476 15428 15528 15434
rect 15566 15399 15622 15408
rect 15476 15370 15528 15376
rect 15672 15201 15700 17274
rect 15764 15609 15792 22320
rect 16132 19938 16160 22320
rect 16040 19910 16160 19938
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15856 17513 15884 17614
rect 15948 17542 15976 19790
rect 16040 18057 16068 19910
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 16132 18834 16160 19790
rect 16212 19780 16264 19786
rect 16212 19722 16264 19728
rect 16120 18828 16172 18834
rect 16120 18770 16172 18776
rect 16118 18456 16174 18465
rect 16118 18391 16174 18400
rect 16132 18222 16160 18391
rect 16120 18216 16172 18222
rect 16120 18158 16172 18164
rect 16026 18048 16082 18057
rect 16026 17983 16082 17992
rect 16028 17672 16080 17678
rect 16026 17640 16028 17649
rect 16080 17640 16082 17649
rect 16026 17575 16082 17584
rect 15936 17536 15988 17542
rect 15842 17504 15898 17513
rect 15936 17478 15988 17484
rect 15842 17439 15898 17448
rect 16026 16824 16082 16833
rect 15936 16788 15988 16794
rect 16026 16759 16082 16768
rect 15936 16730 15988 16736
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15856 16250 15884 16390
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15750 15600 15806 15609
rect 15750 15535 15806 15544
rect 15842 15464 15898 15473
rect 15842 15399 15898 15408
rect 15658 15192 15714 15201
rect 15658 15127 15714 15136
rect 15382 15056 15438 15065
rect 15382 14991 15384 15000
rect 15436 14991 15438 15000
rect 15384 14962 15436 14968
rect 15396 14931 15424 14962
rect 15476 14952 15528 14958
rect 15474 14920 15476 14929
rect 15528 14920 15530 14929
rect 15856 14890 15884 15399
rect 15474 14855 15530 14864
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 15476 14816 15528 14822
rect 15396 14776 15476 14804
rect 15396 13190 15424 14776
rect 15476 14758 15528 14764
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15566 14104 15622 14113
rect 15566 14039 15622 14048
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 13530 15516 13670
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15580 13274 15608 14039
rect 15488 13246 15608 13274
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15488 12918 15516 13246
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15488 12617 15516 12854
rect 15474 12608 15530 12617
rect 15474 12543 15530 12552
rect 15474 12472 15530 12481
rect 15474 12407 15530 12416
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15396 11762 15424 12174
rect 15488 11801 15516 12407
rect 15580 12322 15608 13126
rect 15764 12442 15792 14758
rect 15844 14476 15896 14482
rect 15844 14418 15896 14424
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15580 12294 15792 12322
rect 15568 12164 15620 12170
rect 15568 12106 15620 12112
rect 15474 11792 15530 11801
rect 15384 11756 15436 11762
rect 15474 11727 15530 11736
rect 15384 11698 15436 11704
rect 15488 11150 15516 11727
rect 15580 11393 15608 12106
rect 15566 11384 15622 11393
rect 15566 11319 15622 11328
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15476 11144 15528 11150
rect 15672 11121 15700 11290
rect 15476 11086 15528 11092
rect 15658 11112 15714 11121
rect 15658 11047 15714 11056
rect 15384 10600 15436 10606
rect 15436 10560 15516 10588
rect 15384 10542 15436 10548
rect 15382 10432 15438 10441
rect 15382 10367 15438 10376
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15120 9302 15240 9330
rect 15120 9058 15148 9302
rect 15198 9208 15254 9217
rect 15198 9143 15200 9152
rect 15252 9143 15254 9152
rect 15200 9114 15252 9120
rect 15292 9104 15344 9110
rect 15016 9036 15068 9042
rect 15120 9030 15240 9058
rect 15292 9046 15344 9052
rect 15016 8978 15068 8984
rect 14752 8894 14964 8922
rect 14646 8528 14702 8537
rect 14752 8514 14780 8894
rect 14936 8838 14964 8894
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14702 8486 14780 8514
rect 15016 8492 15068 8498
rect 14646 8463 14702 8472
rect 15016 8434 15068 8440
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 15028 8090 15056 8434
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 14648 8016 14700 8022
rect 14568 7976 14648 8004
rect 14648 7958 14700 7964
rect 14660 7342 14688 7958
rect 15028 7886 15056 8026
rect 15120 8022 15148 8366
rect 15212 8294 15240 9030
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 15304 8090 15332 9046
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15108 8016 15160 8022
rect 15108 7958 15160 7964
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14936 7478 14964 7686
rect 15396 7562 15424 10367
rect 15488 7954 15516 10560
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15764 10418 15792 12294
rect 15856 12170 15884 14418
rect 15948 14278 15976 16730
rect 16040 16590 16068 16759
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 16132 16153 16160 18158
rect 16224 16425 16252 19722
rect 16302 19544 16358 19553
rect 16302 19479 16358 19488
rect 16316 18272 16344 19479
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16408 18601 16436 19110
rect 16394 18592 16450 18601
rect 16394 18527 16450 18536
rect 16316 18244 16436 18272
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16316 17338 16344 18090
rect 16408 18086 16436 18244
rect 16500 18193 16528 22320
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16486 18184 16542 18193
rect 16486 18119 16542 18128
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16210 16416 16266 16425
rect 16210 16351 16266 16360
rect 16118 16144 16174 16153
rect 16118 16079 16174 16088
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16316 15994 16344 16730
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16408 16114 16436 16526
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16028 15904 16080 15910
rect 16028 15846 16080 15852
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16040 15366 16068 15846
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 16026 15192 16082 15201
rect 16026 15127 16082 15136
rect 16040 14482 16068 15127
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 15948 13569 15976 14214
rect 15934 13560 15990 13569
rect 15934 13495 15990 13504
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15948 12918 15976 13262
rect 16040 12986 16068 14214
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 16026 12608 16082 12617
rect 16026 12543 16082 12552
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 15844 12164 15896 12170
rect 15844 12106 15896 12112
rect 15842 11928 15898 11937
rect 15948 11898 15976 12378
rect 15842 11863 15844 11872
rect 15896 11863 15898 11872
rect 15936 11892 15988 11898
rect 15844 11834 15896 11840
rect 15936 11834 15988 11840
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 15856 11286 15884 11698
rect 15948 11694 15976 11834
rect 16040 11694 16068 12543
rect 16132 12481 16160 15846
rect 16224 12753 16252 15982
rect 16316 15966 16436 15994
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16316 15706 16344 15846
rect 16304 15700 16356 15706
rect 16304 15642 16356 15648
rect 16302 15056 16358 15065
rect 16302 14991 16358 15000
rect 16316 14074 16344 14991
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16302 13968 16358 13977
rect 16302 13903 16358 13912
rect 16316 12782 16344 13903
rect 16408 13297 16436 15966
rect 16500 14521 16528 17682
rect 16592 16794 16620 19858
rect 16776 19689 16804 19858
rect 16762 19680 16818 19689
rect 16762 19615 16818 19624
rect 16868 19242 16896 22320
rect 16948 19984 17000 19990
rect 16948 19926 17000 19932
rect 16960 19378 16988 19926
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 16856 19236 16908 19242
rect 16856 19178 16908 19184
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16856 18692 16908 18698
rect 16856 18634 16908 18640
rect 16764 18624 16816 18630
rect 16684 18584 16764 18612
rect 16684 17338 16712 18584
rect 16764 18566 16816 18572
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16580 16516 16632 16522
rect 16580 16458 16632 16464
rect 16486 14512 16542 14521
rect 16486 14447 16542 14456
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16394 13288 16450 13297
rect 16394 13223 16450 13232
rect 16304 12776 16356 12782
rect 16210 12744 16266 12753
rect 16304 12718 16356 12724
rect 16210 12679 16266 12688
rect 16118 12472 16174 12481
rect 16118 12407 16174 12416
rect 16224 12186 16252 12679
rect 16408 12617 16436 13223
rect 16500 12986 16528 14350
rect 16592 13394 16620 16458
rect 16684 15434 16712 17138
rect 16776 16182 16804 18158
rect 16868 16522 16896 18634
rect 16960 16998 16988 18770
rect 17052 18766 17080 19246
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 17052 18329 17080 18702
rect 17038 18320 17094 18329
rect 17038 18255 17094 18264
rect 17040 17740 17092 17746
rect 17040 17682 17092 17688
rect 17052 17134 17080 17682
rect 17040 17128 17092 17134
rect 17040 17070 17092 17076
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 16856 16516 16908 16522
rect 16856 16458 16908 16464
rect 16764 16176 16816 16182
rect 16764 16118 16816 16124
rect 16960 16114 16988 16934
rect 17052 16697 17080 16934
rect 17144 16794 17172 19654
rect 17328 18970 17356 22320
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17512 19825 17540 19858
rect 17498 19816 17554 19825
rect 17498 19751 17554 19760
rect 17590 19680 17646 19689
rect 17590 19615 17646 19624
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 17236 18873 17264 18906
rect 17222 18864 17278 18873
rect 17222 18799 17278 18808
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17236 18426 17264 18566
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 17224 18216 17276 18222
rect 17224 18158 17276 18164
rect 17236 18057 17264 18158
rect 17222 18048 17278 18057
rect 17222 17983 17278 17992
rect 17328 17338 17356 18226
rect 17316 17332 17368 17338
rect 17316 17274 17368 17280
rect 17222 16960 17278 16969
rect 17222 16895 17278 16904
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 17038 16688 17094 16697
rect 17038 16623 17094 16632
rect 17144 16572 17172 16730
rect 17052 16544 17172 16572
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 17052 15722 17080 16544
rect 17132 16176 17184 16182
rect 17132 16118 17184 16124
rect 17144 15910 17172 16118
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17052 15694 17172 15722
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 16672 15428 16724 15434
rect 16672 15370 16724 15376
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16684 14414 16712 14826
rect 16776 14618 16804 15506
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16684 13938 16712 14350
rect 16764 14340 16816 14346
rect 16764 14282 16816 14288
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16580 13388 16632 13394
rect 16632 13348 16712 13376
rect 16580 13330 16632 13336
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16580 12640 16632 12646
rect 16394 12608 16450 12617
rect 16580 12582 16632 12588
rect 16394 12543 16450 12552
rect 16302 12472 16358 12481
rect 16302 12407 16358 12416
rect 16132 12158 16252 12186
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 16132 11529 16160 12158
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16224 11898 16252 12038
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16118 11520 16174 11529
rect 16118 11455 16174 11464
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15856 10606 15884 11086
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15672 10169 15700 10406
rect 15764 10390 15884 10418
rect 15658 10160 15714 10169
rect 15658 10095 15714 10104
rect 15856 10010 15884 10390
rect 15580 9982 15884 10010
rect 15580 9353 15608 9982
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15842 9616 15898 9625
rect 15566 9344 15622 9353
rect 15566 9279 15622 9288
rect 15568 9104 15620 9110
rect 15566 9072 15568 9081
rect 15620 9072 15622 9081
rect 15566 9007 15622 9016
rect 15566 8800 15622 8809
rect 15566 8735 15622 8744
rect 15580 8430 15608 8735
rect 15568 8424 15620 8430
rect 15568 8366 15620 8372
rect 15672 8090 15700 9590
rect 15752 9580 15804 9586
rect 15842 9551 15844 9560
rect 15752 9522 15804 9528
rect 15896 9551 15898 9560
rect 15844 9522 15896 9528
rect 15764 9160 15792 9522
rect 15844 9172 15896 9178
rect 15764 9132 15844 9160
rect 15844 9114 15896 9120
rect 15750 9072 15806 9081
rect 15750 9007 15806 9016
rect 15764 8498 15792 9007
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15856 8294 15884 8774
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15476 7948 15528 7954
rect 15476 7890 15528 7896
rect 15750 7576 15806 7585
rect 15396 7534 15608 7562
rect 14924 7472 14976 7478
rect 14924 7414 14976 7420
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14424 7228 14504 7256
rect 14372 7210 14424 7216
rect 14370 7168 14426 7177
rect 14370 7103 14426 7112
rect 14384 6934 14412 7103
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14200 4214 14228 4558
rect 14384 4264 14412 6326
rect 14476 6254 14504 7228
rect 14556 7268 14608 7274
rect 14556 7210 14608 7216
rect 15108 7268 15160 7274
rect 15108 7210 15160 7216
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14476 5216 14504 5578
rect 14568 5370 14596 7210
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 15120 6934 15148 7210
rect 15108 6928 15160 6934
rect 15108 6870 15160 6876
rect 15108 6656 15160 6662
rect 14922 6624 14978 6633
rect 14922 6559 14978 6568
rect 15106 6624 15108 6633
rect 15160 6624 15162 6633
rect 15106 6559 15162 6568
rect 14936 6361 14964 6559
rect 15212 6497 15240 7346
rect 15292 7200 15344 7206
rect 15290 7168 15292 7177
rect 15344 7168 15346 7177
rect 15290 7103 15346 7112
rect 15396 6798 15424 7346
rect 15476 7268 15528 7274
rect 15476 7210 15528 7216
rect 15488 7002 15516 7210
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15198 6488 15254 6497
rect 15198 6423 15254 6432
rect 14922 6352 14978 6361
rect 14922 6287 14978 6296
rect 15396 6186 15424 6734
rect 15384 6180 15436 6186
rect 15384 6122 15436 6128
rect 15200 6112 15252 6118
rect 15252 6072 15332 6100
rect 15200 6054 15252 6060
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 14556 5364 14608 5370
rect 14608 5324 14688 5352
rect 14556 5306 14608 5312
rect 14660 5234 14688 5324
rect 14556 5228 14608 5234
rect 14476 5188 14556 5216
rect 14556 5170 14608 5176
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14292 4236 14412 4264
rect 14188 4208 14240 4214
rect 14188 4150 14240 4156
rect 14096 4004 14148 4010
rect 14096 3946 14148 3952
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 13820 1624 13872 1630
rect 13820 1566 13872 1572
rect 14016 480 14044 3878
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14108 3058 14136 3538
rect 14200 3534 14228 4150
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14292 3126 14320 4236
rect 14476 3913 14504 4558
rect 14568 4214 14596 5170
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14752 4321 14780 4626
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14738 4312 14794 4321
rect 14844 4282 14872 4422
rect 14738 4247 14794 4256
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 14556 4208 14608 4214
rect 14556 4150 14608 4156
rect 14462 3904 14518 3913
rect 14462 3839 14518 3848
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14830 3632 14886 3641
rect 14830 3567 14832 3576
rect 14884 3567 14886 3576
rect 14832 3538 14884 3544
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14462 3224 14518 3233
rect 14462 3159 14518 3168
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14476 2854 14504 3159
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 14462 2408 14518 2417
rect 14462 2343 14464 2352
rect 14516 2343 14518 2352
rect 14464 2314 14516 2320
rect 14568 1442 14596 3334
rect 14922 3088 14978 3097
rect 14922 3023 14924 3032
rect 14976 3023 14978 3032
rect 14924 2994 14976 3000
rect 14738 2952 14794 2961
rect 15028 2922 15056 5850
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15120 4865 15148 5714
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15212 5030 15240 5646
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15106 4856 15162 4865
rect 15106 4791 15162 4800
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 15120 3942 15148 4422
rect 15212 4146 15240 4762
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15198 4040 15254 4049
rect 15198 3975 15254 3984
rect 15304 3992 15332 6072
rect 15396 5234 15424 6122
rect 15474 5264 15530 5273
rect 15384 5228 15436 5234
rect 15474 5199 15530 5208
rect 15384 5170 15436 5176
rect 15488 4185 15516 5199
rect 15474 4176 15530 4185
rect 15474 4111 15530 4120
rect 15212 3942 15240 3975
rect 15304 3964 15516 3992
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15382 3904 15438 3913
rect 15106 3768 15162 3777
rect 15106 3703 15162 3712
rect 15212 3720 15240 3878
rect 15382 3839 15438 3848
rect 15120 3670 15148 3703
rect 15212 3692 15332 3720
rect 15108 3664 15160 3670
rect 15108 3606 15160 3612
rect 15198 3632 15254 3641
rect 15304 3602 15332 3692
rect 15198 3567 15254 3576
rect 15292 3596 15344 3602
rect 14738 2887 14740 2896
rect 14792 2887 14794 2896
rect 15016 2916 15068 2922
rect 14740 2858 14792 2864
rect 15016 2858 15068 2864
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 15212 2514 15240 3567
rect 15292 3538 15344 3544
rect 15396 3233 15424 3839
rect 15382 3224 15438 3233
rect 15382 3159 15438 3168
rect 15382 2952 15438 2961
rect 15382 2887 15438 2896
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15396 2281 15424 2887
rect 15382 2272 15438 2281
rect 15382 2207 15438 2216
rect 14372 1420 14424 1426
rect 14568 1414 14780 1442
rect 14372 1362 14424 1368
rect 14384 480 14412 1362
rect 14752 480 14780 1414
rect 15108 1284 15160 1290
rect 15108 1226 15160 1232
rect 15120 480 15148 1226
rect 15488 480 15516 3964
rect 15580 2514 15608 7534
rect 15750 7511 15806 7520
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15672 7002 15700 7142
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15764 6934 15792 7511
rect 15842 7304 15898 7313
rect 15842 7239 15898 7248
rect 15752 6928 15804 6934
rect 15752 6870 15804 6876
rect 15764 5930 15792 6870
rect 15672 5902 15792 5930
rect 15672 4486 15700 5902
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 15672 4049 15700 4422
rect 15658 4040 15714 4049
rect 15658 3975 15714 3984
rect 15764 3074 15792 5714
rect 15856 5681 15884 7239
rect 15842 5672 15898 5681
rect 15842 5607 15898 5616
rect 15842 5264 15898 5273
rect 15842 5199 15898 5208
rect 15856 5098 15884 5199
rect 15844 5092 15896 5098
rect 15844 5034 15896 5040
rect 15764 3046 15884 3074
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15856 480 15884 3046
rect 15948 2650 15976 10950
rect 16316 10690 16344 12407
rect 16394 11928 16450 11937
rect 16394 11863 16450 11872
rect 16408 11694 16436 11863
rect 16592 11801 16620 12582
rect 16578 11792 16634 11801
rect 16578 11727 16634 11736
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 16578 11656 16634 11665
rect 16578 11591 16634 11600
rect 16486 11520 16542 11529
rect 16486 11455 16542 11464
rect 16394 11384 16450 11393
rect 16394 11319 16450 11328
rect 16132 10662 16344 10690
rect 16132 10266 16160 10662
rect 16302 10568 16358 10577
rect 16302 10503 16304 10512
rect 16356 10503 16358 10512
rect 16304 10474 16356 10480
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16224 10266 16252 10406
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16210 10160 16266 10169
rect 16210 10095 16266 10104
rect 16026 9616 16082 9625
rect 16026 9551 16082 9560
rect 16040 8838 16068 9551
rect 16118 9480 16174 9489
rect 16118 9415 16174 9424
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 16040 8430 16068 8774
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 16040 7886 16068 8366
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 16040 7546 16068 7822
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16040 6390 16068 6734
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 16040 5710 16068 6326
rect 16132 5914 16160 9415
rect 16224 8514 16252 10095
rect 16408 9625 16436 11319
rect 16394 9616 16450 9625
rect 16394 9551 16450 9560
rect 16302 9480 16358 9489
rect 16302 9415 16304 9424
rect 16356 9415 16358 9424
rect 16304 9386 16356 9392
rect 16394 9344 16450 9353
rect 16394 9279 16450 9288
rect 16304 8900 16356 8906
rect 16304 8842 16356 8848
rect 16316 8809 16344 8842
rect 16302 8800 16358 8809
rect 16302 8735 16358 8744
rect 16224 8486 16344 8514
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 16224 7546 16252 8298
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16212 7200 16264 7206
rect 16210 7168 16212 7177
rect 16264 7168 16266 7177
rect 16210 7103 16266 7112
rect 16316 7018 16344 8486
rect 16408 8378 16436 9279
rect 16500 9178 16528 11455
rect 16592 10470 16620 11591
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16592 9217 16620 9658
rect 16578 9208 16634 9217
rect 16488 9172 16540 9178
rect 16578 9143 16634 9152
rect 16488 9114 16540 9120
rect 16486 9072 16542 9081
rect 16486 9007 16542 9016
rect 16580 9036 16632 9042
rect 16500 8537 16528 9007
rect 16580 8978 16632 8984
rect 16486 8528 16542 8537
rect 16486 8463 16542 8472
rect 16408 8350 16528 8378
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16224 6990 16344 7018
rect 16224 6769 16252 6990
rect 16210 6760 16266 6769
rect 16210 6695 16266 6704
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 16040 5098 16068 5646
rect 16028 5092 16080 5098
rect 16028 5034 16080 5040
rect 16040 4826 16068 5034
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 16040 4146 16068 4558
rect 16224 4298 16252 4626
rect 16224 4270 16344 4298
rect 16028 4140 16080 4146
rect 16028 4082 16080 4088
rect 16040 3534 16068 4082
rect 16316 3942 16344 4270
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 16040 2922 16068 3470
rect 16028 2916 16080 2922
rect 16028 2858 16080 2864
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16224 2106 16252 2858
rect 16408 2582 16436 8230
rect 16500 7410 16528 8350
rect 16592 7993 16620 8978
rect 16578 7984 16634 7993
rect 16578 7919 16634 7928
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16500 6769 16528 7346
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16486 6760 16542 6769
rect 16486 6695 16542 6704
rect 16592 5642 16620 7142
rect 16580 5636 16632 5642
rect 16580 5578 16632 5584
rect 16578 5400 16634 5409
rect 16578 5335 16634 5344
rect 16592 3602 16620 5335
rect 16684 3942 16712 13348
rect 16776 12782 16804 14282
rect 16868 14074 16896 15438
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 16948 14884 17000 14890
rect 16948 14826 17000 14832
rect 16960 14385 16988 14826
rect 17052 14482 17080 14894
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 16946 14376 17002 14385
rect 16946 14311 17002 14320
rect 17052 14074 17080 14418
rect 16856 14068 16908 14074
rect 17040 14068 17092 14074
rect 16856 14010 16908 14016
rect 16960 14028 17040 14056
rect 16856 13796 16908 13802
rect 16856 13738 16908 13744
rect 16868 13462 16896 13738
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16960 13410 16988 14028
rect 17040 14010 17092 14016
rect 17144 13954 17172 15694
rect 17052 13926 17172 13954
rect 17052 13569 17080 13926
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17038 13560 17094 13569
rect 17144 13530 17172 13670
rect 17038 13495 17094 13504
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 16960 13382 17080 13410
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16868 13161 16896 13262
rect 16854 13152 16910 13161
rect 16854 13087 16910 13096
rect 16960 12850 16988 13262
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 17052 12442 17080 13382
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 17236 12220 17264 16895
rect 17316 16720 17368 16726
rect 17314 16688 17316 16697
rect 17368 16688 17370 16697
rect 17314 16623 17370 16632
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17328 15638 17356 15846
rect 17316 15632 17368 15638
rect 17316 15574 17368 15580
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17420 15450 17448 19314
rect 17500 19304 17552 19310
rect 17498 19272 17500 19281
rect 17552 19272 17554 19281
rect 17498 19207 17554 19216
rect 17604 19145 17632 19615
rect 17590 19136 17646 19145
rect 17590 19071 17646 19080
rect 17696 18986 17724 22320
rect 17958 21040 18014 21049
rect 17958 20975 18014 20984
rect 17972 19990 18000 20975
rect 18064 20058 18092 22320
rect 18142 21448 18198 21457
rect 18142 21383 18198 21392
rect 18156 20738 18184 21383
rect 18144 20732 18196 20738
rect 18144 20674 18196 20680
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 17960 19984 18012 19990
rect 17960 19926 18012 19932
rect 18432 19802 18460 22320
rect 18800 20754 18828 22320
rect 18800 20726 19012 20754
rect 18786 20632 18842 20641
rect 18786 20567 18842 20576
rect 18432 19774 18552 19802
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17776 19236 17828 19242
rect 17776 19178 17828 19184
rect 17604 18958 17724 18986
rect 17604 18902 17632 18958
rect 17592 18896 17644 18902
rect 17592 18838 17644 18844
rect 17682 18864 17738 18873
rect 17500 18828 17552 18834
rect 17682 18799 17738 18808
rect 17500 18770 17552 18776
rect 17512 17678 17540 18770
rect 17696 18193 17724 18799
rect 17682 18184 17738 18193
rect 17682 18119 17738 18128
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 17590 17776 17646 17785
rect 17590 17711 17646 17720
rect 17604 17678 17632 17711
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17512 15570 17540 17274
rect 17604 17134 17632 17478
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17604 16697 17632 16730
rect 17590 16688 17646 16697
rect 17590 16623 17646 16632
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 17328 14822 17356 15438
rect 17420 15422 17540 15450
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17328 14482 17356 14758
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17328 13326 17356 14418
rect 17420 13530 17448 15302
rect 17512 15094 17540 15422
rect 17500 15088 17552 15094
rect 17500 15030 17552 15036
rect 17604 14793 17632 16390
rect 17696 16114 17724 18022
rect 17788 16590 17816 19178
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17880 17882 17908 19110
rect 17972 18873 18000 19450
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 17958 18864 18014 18873
rect 17958 18799 18014 18808
rect 18156 18737 18184 19178
rect 18142 18728 18198 18737
rect 18142 18663 18198 18672
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 17960 18352 18012 18358
rect 17958 18320 17960 18329
rect 18012 18320 18014 18329
rect 18524 18290 18552 19774
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18616 18737 18644 19654
rect 18696 19304 18748 19310
rect 18696 19246 18748 19252
rect 18602 18728 18658 18737
rect 18602 18663 18658 18672
rect 18604 18352 18656 18358
rect 18604 18294 18656 18300
rect 17958 18255 18014 18264
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17880 17377 17908 17478
rect 17866 17368 17922 17377
rect 17866 17303 17922 17312
rect 17972 17241 18000 18090
rect 18236 18080 18288 18086
rect 18420 18080 18472 18086
rect 18236 18022 18288 18028
rect 18418 18048 18420 18057
rect 18472 18048 18474 18057
rect 18248 17921 18276 18022
rect 18418 17983 18474 17992
rect 18050 17912 18106 17921
rect 18050 17847 18106 17856
rect 18234 17912 18290 17921
rect 18234 17847 18290 17856
rect 18064 17814 18092 17847
rect 18052 17808 18104 17814
rect 18052 17750 18104 17756
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 17958 17232 18014 17241
rect 17958 17167 18014 17176
rect 18616 17105 18644 18294
rect 18602 17096 18658 17105
rect 18328 17060 18380 17066
rect 18602 17031 18658 17040
rect 18328 17002 18380 17008
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17868 16516 17920 16522
rect 17868 16458 17920 16464
rect 17774 16144 17830 16153
rect 17684 16108 17736 16114
rect 17774 16079 17830 16088
rect 17684 16050 17736 16056
rect 17590 14784 17646 14793
rect 17590 14719 17646 14728
rect 17788 14618 17816 16079
rect 17880 15609 17908 16458
rect 17972 16250 18000 16934
rect 18340 16658 18368 17002
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 18432 16522 18460 16934
rect 18420 16516 18472 16522
rect 18420 16458 18472 16464
rect 18604 16516 18656 16522
rect 18604 16458 18656 16464
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 17866 15600 17922 15609
rect 17866 15535 17922 15544
rect 17960 15496 18012 15502
rect 17880 15456 17960 15484
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17316 12912 17368 12918
rect 17316 12854 17368 12860
rect 16868 12192 17264 12220
rect 16762 11928 16818 11937
rect 16762 11863 16818 11872
rect 16776 11558 16804 11863
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16762 10976 16818 10985
rect 16762 10911 16818 10920
rect 16776 9722 16804 10911
rect 16764 9716 16816 9722
rect 16764 9658 16816 9664
rect 16868 9654 16896 12192
rect 17328 11830 17356 12854
rect 17512 12306 17540 14010
rect 17604 13734 17632 14418
rect 17880 14396 17908 15456
rect 17960 15438 18012 15444
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17972 14550 18000 15302
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18524 15144 18552 16186
rect 18616 16017 18644 16458
rect 18602 16008 18658 16017
rect 18602 15943 18658 15952
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18616 15745 18644 15846
rect 18602 15736 18658 15745
rect 18602 15671 18658 15680
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18340 15116 18552 15144
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 18142 14784 18198 14793
rect 18142 14719 18198 14728
rect 17960 14544 18012 14550
rect 17960 14486 18012 14492
rect 18052 14544 18104 14550
rect 18052 14486 18104 14492
rect 18064 14396 18092 14486
rect 17682 14376 17738 14385
rect 17682 14311 17738 14320
rect 17880 14368 18092 14396
rect 17696 14278 17724 14311
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17682 13968 17738 13977
rect 17682 13903 17738 13912
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17590 12880 17646 12889
rect 17590 12815 17646 12824
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17316 11824 17368 11830
rect 16946 11792 17002 11801
rect 17316 11766 17368 11772
rect 16946 11727 17002 11736
rect 16856 9648 16908 9654
rect 16856 9590 16908 9596
rect 16762 8664 16818 8673
rect 16762 8599 16818 8608
rect 16776 8401 16804 8599
rect 16868 8430 16896 9590
rect 16960 9353 16988 11727
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17144 11286 17172 11494
rect 17132 11280 17184 11286
rect 17132 11222 17184 11228
rect 17236 11150 17264 11630
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 17224 11144 17276 11150
rect 17224 11086 17276 11092
rect 17052 10266 17080 11086
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17144 10674 17172 10950
rect 17328 10810 17356 11494
rect 17420 11218 17448 11494
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17512 10674 17540 12242
rect 17604 11218 17632 12815
rect 17696 11898 17724 13903
rect 17788 13394 17816 14214
rect 17880 13802 17908 14368
rect 18156 14346 18184 14719
rect 18248 14521 18276 14962
rect 18234 14512 18290 14521
rect 18234 14447 18236 14456
rect 18288 14447 18290 14456
rect 18236 14418 18288 14424
rect 18340 14396 18368 15116
rect 18418 14920 18474 14929
rect 18418 14855 18420 14864
rect 18472 14855 18474 14864
rect 18420 14826 18472 14832
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18524 14521 18552 14758
rect 18510 14512 18566 14521
rect 18510 14447 18566 14456
rect 18340 14368 18552 14396
rect 18144 14340 18196 14346
rect 17972 14300 18144 14328
rect 17972 13938 18000 14300
rect 18144 14282 18196 14288
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 18050 13832 18106 13841
rect 17868 13796 17920 13802
rect 18050 13767 18106 13776
rect 17868 13738 17920 13744
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17776 13388 17828 13394
rect 17776 13330 17828 13336
rect 17776 12300 17828 12306
rect 17880 12288 17908 13466
rect 17972 12646 18000 13670
rect 18064 13394 18092 13767
rect 18418 13560 18474 13569
rect 18418 13495 18474 13504
rect 18234 13424 18290 13433
rect 18052 13388 18104 13394
rect 18234 13359 18290 13368
rect 18052 13330 18104 13336
rect 18248 13326 18276 13359
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18432 13172 18460 13495
rect 18524 13444 18552 14368
rect 18616 13546 18644 15506
rect 18708 13705 18736 19246
rect 18800 18902 18828 20567
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 18892 19825 18920 19858
rect 18878 19816 18934 19825
rect 18878 19751 18934 19760
rect 18892 19514 18920 19751
rect 18880 19508 18932 19514
rect 18880 19450 18932 19456
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 18788 18896 18840 18902
rect 18788 18838 18840 18844
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18800 16522 18828 18702
rect 18892 17513 18920 19110
rect 18984 18834 19012 20726
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 18972 18828 19024 18834
rect 18972 18770 19024 18776
rect 18972 18624 19024 18630
rect 18972 18566 19024 18572
rect 18878 17504 18934 17513
rect 18878 17439 18934 17448
rect 18880 17196 18932 17202
rect 18880 17138 18932 17144
rect 18892 17105 18920 17138
rect 18878 17096 18934 17105
rect 18878 17031 18934 17040
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18788 16516 18840 16522
rect 18788 16458 18840 16464
rect 18800 16250 18828 16458
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 18892 15688 18920 16934
rect 18984 16182 19012 18566
rect 19076 17762 19104 20198
rect 19168 19009 19196 22320
rect 19246 22264 19302 22273
rect 19246 22199 19302 22208
rect 19154 19000 19210 19009
rect 19154 18935 19210 18944
rect 19156 18828 19208 18834
rect 19156 18770 19208 18776
rect 19168 18426 19196 18770
rect 19156 18420 19208 18426
rect 19156 18362 19208 18368
rect 19260 18290 19288 22199
rect 19340 18896 19392 18902
rect 19340 18838 19392 18844
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19156 18216 19208 18222
rect 19154 18184 19156 18193
rect 19208 18184 19210 18193
rect 19154 18119 19210 18128
rect 19156 18080 19208 18086
rect 19154 18048 19156 18057
rect 19208 18048 19210 18057
rect 19154 17983 19210 17992
rect 19076 17734 19288 17762
rect 19064 17672 19116 17678
rect 19064 17614 19116 17620
rect 18972 16176 19024 16182
rect 18972 16118 19024 16124
rect 18800 15660 18920 15688
rect 18694 13696 18750 13705
rect 18694 13631 18750 13640
rect 18616 13518 18736 13546
rect 18708 13462 18736 13518
rect 18696 13456 18748 13462
rect 18524 13416 18644 13444
rect 18616 13308 18644 13416
rect 18696 13398 18748 13404
rect 18800 13376 18828 15660
rect 18972 15632 19024 15638
rect 18970 15600 18972 15609
rect 19024 15600 19026 15609
rect 18970 15535 19026 15544
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18892 14929 18920 15438
rect 19076 15178 19104 17614
rect 19260 17066 19288 17734
rect 19156 17060 19208 17066
rect 19156 17002 19208 17008
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 18984 15150 19104 15178
rect 18878 14920 18934 14929
rect 18878 14855 18934 14864
rect 18878 14784 18934 14793
rect 18878 14719 18934 14728
rect 18892 13569 18920 14719
rect 18878 13560 18934 13569
rect 18878 13495 18934 13504
rect 18800 13348 18920 13376
rect 18616 13280 18736 13308
rect 18432 13144 18552 13172
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18420 12708 18472 12714
rect 18420 12650 18472 12656
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17960 12368 18012 12374
rect 17960 12310 18012 12316
rect 17828 12260 17908 12288
rect 17776 12242 17828 12248
rect 17866 12064 17922 12073
rect 17866 11999 17922 12008
rect 17774 11928 17830 11937
rect 17684 11892 17736 11898
rect 17774 11863 17776 11872
rect 17684 11834 17736 11840
rect 17828 11863 17830 11872
rect 17776 11834 17828 11840
rect 17774 11792 17830 11801
rect 17774 11727 17830 11736
rect 17682 11656 17738 11665
rect 17682 11591 17738 11600
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17500 10668 17552 10674
rect 17552 10628 17632 10656
rect 17500 10610 17552 10616
rect 17314 10568 17370 10577
rect 17132 10532 17184 10538
rect 17314 10503 17316 10512
rect 17132 10474 17184 10480
rect 17368 10503 17370 10512
rect 17316 10474 17368 10480
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 17144 10130 17172 10474
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17314 10296 17370 10305
rect 17314 10231 17370 10240
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17224 10056 17276 10062
rect 17222 10024 17224 10033
rect 17276 10024 17278 10033
rect 17222 9959 17278 9968
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 17052 9586 17080 9862
rect 17222 9616 17278 9625
rect 17040 9580 17092 9586
rect 17222 9551 17278 9560
rect 17040 9522 17092 9528
rect 17052 9489 17080 9522
rect 17038 9480 17094 9489
rect 17038 9415 17094 9424
rect 16946 9344 17002 9353
rect 16946 9279 17002 9288
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16856 8424 16908 8430
rect 16762 8392 16818 8401
rect 16856 8366 16908 8372
rect 16762 8327 16818 8336
rect 16854 7848 16910 7857
rect 16854 7783 16910 7792
rect 16868 7546 16896 7783
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16868 7410 16896 7482
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16856 6996 16908 7002
rect 16856 6938 16908 6944
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 16500 2990 16528 3470
rect 16488 2984 16540 2990
rect 16488 2926 16540 2932
rect 16488 2848 16540 2854
rect 16540 2796 16620 2802
rect 16488 2790 16620 2796
rect 16500 2774 16620 2790
rect 16396 2576 16448 2582
rect 16396 2518 16448 2524
rect 16304 2304 16356 2310
rect 16304 2246 16356 2252
rect 16212 2100 16264 2106
rect 16212 2042 16264 2048
rect 16316 2009 16344 2246
rect 16592 2106 16620 2774
rect 16580 2100 16632 2106
rect 16580 2042 16632 2048
rect 16302 2000 16358 2009
rect 16684 1986 16712 3878
rect 16302 1935 16358 1944
rect 16500 1958 16712 1986
rect 16212 1624 16264 1630
rect 16212 1566 16264 1572
rect 16224 480 16252 1566
rect 16500 513 16528 1958
rect 16776 1442 16804 6598
rect 16868 5778 16896 6938
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16868 5370 16896 5714
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16868 3670 16896 4558
rect 16960 4185 16988 8978
rect 17052 8412 17080 9415
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17144 8566 17172 8910
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17052 8384 17172 8412
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 17052 7002 17080 7822
rect 17040 6996 17092 7002
rect 17040 6938 17092 6944
rect 17038 5944 17094 5953
rect 17038 5879 17094 5888
rect 17052 5778 17080 5879
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 17052 5370 17080 5714
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 16946 4176 17002 4185
rect 16946 4111 17002 4120
rect 16946 4040 17002 4049
rect 16946 3975 17002 3984
rect 16960 3942 16988 3975
rect 17052 3942 17080 4558
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 16856 3664 16908 3670
rect 16856 3606 16908 3612
rect 17052 3194 17080 3878
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 16948 3120 17000 3126
rect 17144 3074 17172 8384
rect 17236 7206 17264 9551
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17224 6928 17276 6934
rect 17224 6870 17276 6876
rect 17236 4826 17264 6870
rect 17328 6633 17356 10231
rect 17420 8129 17448 10406
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17512 10062 17540 10202
rect 17604 10062 17632 10628
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17500 9648 17552 9654
rect 17500 9590 17552 9596
rect 17590 9616 17646 9625
rect 17512 9160 17540 9590
rect 17590 9551 17646 9560
rect 17604 9518 17632 9551
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17512 9132 17632 9160
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17406 8120 17462 8129
rect 17406 8055 17462 8064
rect 17408 6656 17460 6662
rect 17314 6624 17370 6633
rect 17408 6598 17460 6604
rect 17314 6559 17370 6568
rect 17420 6322 17448 6598
rect 17512 6458 17540 8978
rect 17604 8294 17632 9132
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17696 8090 17724 11591
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17604 6662 17632 7890
rect 17788 7546 17816 11727
rect 17880 11393 17908 11999
rect 17972 11694 18000 12310
rect 18432 12209 18460 12650
rect 18418 12200 18474 12209
rect 18418 12135 18474 12144
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 18420 11620 18472 11626
rect 18420 11562 18472 11568
rect 17958 11520 18014 11529
rect 17958 11455 18014 11464
rect 17866 11384 17922 11393
rect 17866 11319 17922 11328
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17880 10538 17908 11086
rect 17868 10532 17920 10538
rect 17868 10474 17920 10480
rect 17866 10432 17922 10441
rect 17972 10418 18000 11455
rect 18144 11280 18196 11286
rect 18142 11248 18144 11257
rect 18196 11248 18198 11257
rect 18142 11183 18198 11192
rect 18432 11082 18460 11562
rect 18524 11354 18552 13144
rect 18602 13152 18658 13161
rect 18602 13087 18658 13096
rect 18616 12850 18644 13087
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18708 12220 18736 13280
rect 18788 13252 18840 13258
rect 18788 13194 18840 13200
rect 18800 13161 18828 13194
rect 18786 13152 18842 13161
rect 18786 13087 18842 13096
rect 18892 12968 18920 13348
rect 18800 12940 18920 12968
rect 18800 12850 18828 12940
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18880 12776 18932 12782
rect 18786 12744 18842 12753
rect 18880 12718 18932 12724
rect 18786 12679 18842 12688
rect 18616 12192 18736 12220
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18420 11076 18472 11082
rect 18420 11018 18472 11024
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18418 10704 18474 10713
rect 18418 10639 18474 10648
rect 18144 10600 18196 10606
rect 18196 10560 18276 10588
rect 18144 10542 18196 10548
rect 18248 10554 18276 10560
rect 18248 10526 18368 10554
rect 17922 10390 18000 10418
rect 17866 10367 17922 10376
rect 17972 10282 18000 10390
rect 17972 10254 18092 10282
rect 18064 10146 18092 10254
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 17972 10118 18092 10146
rect 18248 10130 18276 10202
rect 18236 10124 18288 10130
rect 17972 9602 18000 10118
rect 18236 10066 18288 10072
rect 18340 10062 18368 10526
rect 18432 10130 18460 10639
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18340 9908 18368 9998
rect 18340 9880 18552 9908
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18144 9648 18196 9654
rect 17972 9574 18092 9602
rect 18144 9590 18196 9596
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17880 7546 17908 9318
rect 17958 9072 18014 9081
rect 17958 9007 17960 9016
rect 18012 9007 18014 9016
rect 17960 8978 18012 8984
rect 18064 8888 18092 9574
rect 18156 9518 18184 9590
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18156 8906 18184 9114
rect 18524 9081 18552 9880
rect 18616 9110 18644 12192
rect 18694 12064 18750 12073
rect 18694 11999 18750 12008
rect 18604 9104 18656 9110
rect 18326 9072 18382 9081
rect 18326 9007 18328 9016
rect 18380 9007 18382 9016
rect 18510 9072 18566 9081
rect 18604 9046 18656 9052
rect 18510 9007 18566 9016
rect 18328 8978 18380 8984
rect 17972 8860 18092 8888
rect 18144 8900 18196 8906
rect 17972 7936 18000 8860
rect 18144 8842 18196 8848
rect 18510 8800 18566 8809
rect 18116 8732 18412 8752
rect 18510 8735 18566 8744
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 18524 8634 18552 8735
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18420 8492 18472 8498
rect 18472 8452 18552 8480
rect 18420 8434 18472 8440
rect 18052 7948 18104 7954
rect 17972 7908 18052 7936
rect 18052 7890 18104 7896
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 18524 7546 18552 8452
rect 18616 7750 18644 9046
rect 18708 8430 18736 11999
rect 18800 9994 18828 12679
rect 18892 12442 18920 12718
rect 18984 12442 19012 15150
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 19076 13462 19104 14758
rect 19064 13456 19116 13462
rect 19064 13398 19116 13404
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 19076 12782 19104 13262
rect 19064 12776 19116 12782
rect 19062 12744 19064 12753
rect 19116 12744 19118 12753
rect 19062 12679 19118 12688
rect 19076 12653 19104 12679
rect 19062 12608 19118 12617
rect 19062 12543 19118 12552
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 18892 11694 18920 12378
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18878 11520 18934 11529
rect 18878 11455 18934 11464
rect 18892 10554 18920 11455
rect 18984 11354 19012 12242
rect 19076 11393 19104 12543
rect 19062 11384 19118 11393
rect 18972 11348 19024 11354
rect 19062 11319 19118 11328
rect 18972 11290 19024 11296
rect 18972 11212 19024 11218
rect 18972 11154 19024 11160
rect 18984 10656 19012 11154
rect 19076 10810 19104 11319
rect 19064 10804 19116 10810
rect 19064 10746 19116 10752
rect 18984 10628 19104 10656
rect 18892 10526 19012 10554
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 18788 9988 18840 9994
rect 18788 9930 18840 9936
rect 18788 9580 18840 9586
rect 18892 9568 18920 10406
rect 18840 9540 18920 9568
rect 18788 9522 18840 9528
rect 18800 8498 18828 9522
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18708 8265 18736 8366
rect 18694 8256 18750 8265
rect 18694 8191 18750 8200
rect 18786 8120 18842 8129
rect 18892 8090 18920 8434
rect 18786 8055 18842 8064
rect 18880 8084 18932 8090
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 17960 7472 18012 7478
rect 17960 7414 18012 7420
rect 18234 7440 18290 7449
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17696 6866 17724 7346
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 17684 6860 17736 6866
rect 17684 6802 17736 6808
rect 17684 6724 17736 6730
rect 17684 6666 17736 6672
rect 17592 6656 17644 6662
rect 17592 6598 17644 6604
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17604 6338 17632 6598
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17512 6310 17632 6338
rect 17512 5574 17540 6310
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 17604 5556 17632 6190
rect 17696 5953 17724 6666
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17682 5944 17738 5953
rect 17682 5879 17738 5888
rect 17788 5642 17816 6054
rect 17776 5636 17828 5642
rect 17776 5578 17828 5584
rect 17684 5568 17736 5574
rect 17604 5528 17684 5556
rect 17498 4992 17554 5001
rect 17498 4927 17554 4936
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 17408 4480 17460 4486
rect 17408 4422 17460 4428
rect 16948 3062 17000 3068
rect 16856 2576 16908 2582
rect 16854 2544 16856 2553
rect 16908 2544 16910 2553
rect 16854 2479 16910 2488
rect 16592 1414 16804 1442
rect 16486 504 16542 513
rect 6090 439 6146 448
rect 6182 0 6238 480
rect 6550 0 6606 480
rect 6918 0 6974 480
rect 7286 0 7342 480
rect 7654 0 7710 480
rect 8022 0 8078 480
rect 8390 0 8446 480
rect 8758 0 8814 480
rect 9126 0 9182 480
rect 9494 0 9550 480
rect 9862 0 9918 480
rect 10230 0 10286 480
rect 10598 0 10654 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12162 0 12218 480
rect 12530 0 12586 480
rect 12898 0 12954 480
rect 13266 0 13322 480
rect 13634 0 13690 480
rect 14002 0 14058 480
rect 14370 0 14426 480
rect 14738 0 14794 480
rect 15106 0 15162 480
rect 15474 0 15530 480
rect 15842 0 15898 480
rect 16210 0 16266 480
rect 16592 480 16620 1414
rect 16960 480 16988 3062
rect 17052 3046 17172 3074
rect 17224 3052 17276 3058
rect 17052 2514 17080 3046
rect 17224 2994 17276 3000
rect 17130 2680 17186 2689
rect 17130 2615 17132 2624
rect 17184 2615 17186 2624
rect 17132 2586 17184 2592
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17236 1630 17264 2994
rect 17328 2310 17356 4422
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17224 1624 17276 1630
rect 17224 1566 17276 1572
rect 17420 480 17448 4422
rect 17512 2650 17540 4927
rect 17604 3670 17632 5528
rect 17880 5522 17908 6938
rect 17972 6322 18000 7414
rect 18234 7375 18290 7384
rect 18248 7002 18276 7375
rect 18326 7032 18382 7041
rect 18236 6996 18288 7002
rect 18326 6967 18328 6976
rect 18236 6938 18288 6944
rect 18380 6967 18382 6976
rect 18512 6996 18564 7002
rect 18328 6938 18380 6944
rect 18512 6938 18564 6944
rect 18524 6905 18552 6938
rect 18510 6896 18566 6905
rect 18510 6831 18566 6840
rect 18328 6792 18380 6798
rect 18326 6760 18328 6769
rect 18380 6760 18382 6769
rect 18326 6695 18382 6704
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 17684 5510 17736 5516
rect 17788 5494 17908 5522
rect 17788 4826 17816 5494
rect 17972 5370 18000 6122
rect 18340 6118 18368 6258
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 18328 6112 18380 6118
rect 18328 6054 18380 6060
rect 18064 5914 18092 6054
rect 18142 5944 18198 5953
rect 18052 5908 18104 5914
rect 18142 5879 18198 5888
rect 18052 5850 18104 5856
rect 18156 5710 18184 5879
rect 18326 5808 18382 5817
rect 18326 5743 18328 5752
rect 18380 5743 18382 5752
rect 18328 5714 18380 5720
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 18512 5024 18564 5030
rect 18512 4966 18564 4972
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 17684 4208 17736 4214
rect 17684 4150 17736 4156
rect 17592 3664 17644 3670
rect 17592 3606 17644 3612
rect 17696 3126 17724 4150
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 17592 2576 17644 2582
rect 17592 2518 17644 2524
rect 17604 1562 17632 2518
rect 17684 2508 17736 2514
rect 17684 2450 17736 2456
rect 17696 2417 17724 2450
rect 17682 2408 17738 2417
rect 17682 2343 17738 2352
rect 17592 1556 17644 1562
rect 17592 1498 17644 1504
rect 17788 480 17816 4218
rect 18050 4176 18106 4185
rect 17960 4140 18012 4146
rect 18050 4111 18052 4120
rect 17960 4082 18012 4088
rect 18104 4111 18106 4120
rect 18052 4082 18104 4088
rect 17972 3670 18000 4082
rect 18064 3738 18092 4082
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 17960 3664 18012 3670
rect 17960 3606 18012 3612
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 17868 3392 17920 3398
rect 18248 3380 18276 3538
rect 17868 3334 17920 3340
rect 17972 3352 18276 3380
rect 17880 3126 17908 3334
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 17972 2854 18000 3352
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 17960 2508 18012 2514
rect 17880 2468 17960 2496
rect 17880 1698 17908 2468
rect 17960 2450 18012 2456
rect 17960 2372 18012 2378
rect 17960 2314 18012 2320
rect 17868 1692 17920 1698
rect 17868 1634 17920 1640
rect 17972 1170 18000 2314
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1142 18184 1170
rect 18156 480 18184 1142
rect 18524 480 18552 4966
rect 18616 2446 18644 7686
rect 18800 7528 18828 8055
rect 18880 8026 18932 8032
rect 18800 7500 18920 7528
rect 18892 7410 18920 7500
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18786 7168 18842 7177
rect 18708 7002 18736 7142
rect 18786 7103 18842 7112
rect 18800 7002 18828 7103
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 18892 6882 18920 7346
rect 18800 6854 18920 6882
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18708 4758 18736 5510
rect 18800 5098 18828 6854
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18892 5166 18920 6190
rect 18880 5160 18932 5166
rect 18880 5102 18932 5108
rect 18788 5092 18840 5098
rect 18788 5034 18840 5040
rect 18696 4752 18748 4758
rect 18696 4694 18748 4700
rect 18788 4684 18840 4690
rect 18788 4626 18840 4632
rect 18696 3664 18748 3670
rect 18800 3641 18828 4626
rect 18892 4185 18920 5102
rect 18878 4176 18934 4185
rect 18878 4111 18934 4120
rect 18696 3606 18748 3612
rect 18786 3632 18842 3641
rect 18708 3058 18736 3606
rect 18984 3602 19012 10526
rect 19076 10130 19104 10628
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 19076 8634 19104 9862
rect 19168 9654 19196 17002
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19260 16697 19288 16730
rect 19246 16688 19302 16697
rect 19246 16623 19302 16632
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19260 16046 19288 16526
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19246 15872 19302 15881
rect 19246 15807 19302 15816
rect 19260 13734 19288 15807
rect 19352 15042 19380 18838
rect 19536 17649 19564 22320
rect 19904 21978 19932 22320
rect 19812 21950 19932 21978
rect 19616 20324 19668 20330
rect 19616 20266 19668 20272
rect 19628 19922 19656 20266
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19628 19360 19656 19858
rect 19628 19332 19748 19360
rect 19616 19236 19668 19242
rect 19616 19178 19668 19184
rect 19522 17640 19578 17649
rect 19522 17575 19578 17584
rect 19524 17536 19576 17542
rect 19524 17478 19576 17484
rect 19536 16697 19564 17478
rect 19628 16794 19656 19178
rect 19720 17814 19748 19332
rect 19812 19310 19840 21950
rect 19890 21856 19946 21865
rect 19890 21791 19946 21800
rect 19904 19990 19932 21791
rect 20364 20330 20392 22320
rect 20352 20324 20404 20330
rect 20352 20266 20404 20272
rect 20350 20224 20406 20233
rect 20350 20159 20406 20168
rect 19892 19984 19944 19990
rect 19892 19926 19944 19932
rect 20364 19922 20392 20159
rect 20640 19990 20668 22607
rect 20718 22320 20774 22800
rect 21086 22320 21142 22800
rect 21454 22320 21510 22800
rect 21822 22320 21878 22800
rect 22190 22320 22246 22800
rect 22558 22320 22614 22800
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 20352 19916 20404 19922
rect 20352 19858 20404 19864
rect 20444 19372 20496 19378
rect 20444 19314 20496 19320
rect 19800 19304 19852 19310
rect 19800 19246 19852 19252
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 19800 18760 19852 18766
rect 19800 18702 19852 18708
rect 19708 17808 19760 17814
rect 19708 17750 19760 17756
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 19522 16688 19578 16697
rect 19522 16623 19578 16632
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 19444 15337 19472 15846
rect 19430 15328 19486 15337
rect 19430 15263 19486 15272
rect 19430 15192 19486 15201
rect 19430 15127 19432 15136
rect 19484 15127 19486 15136
rect 19432 15098 19484 15104
rect 19352 15014 19472 15042
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19352 14657 19380 14758
rect 19338 14648 19394 14657
rect 19338 14583 19394 14592
rect 19338 14512 19394 14521
rect 19338 14447 19394 14456
rect 19352 14346 19380 14447
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19444 14249 19472 15014
rect 19430 14240 19486 14249
rect 19430 14175 19486 14184
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 19246 13560 19302 13569
rect 19246 13495 19302 13504
rect 19260 13025 19288 13495
rect 19352 13326 19380 13874
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19246 13016 19302 13025
rect 19246 12951 19302 12960
rect 19352 12918 19380 13126
rect 19248 12912 19300 12918
rect 19248 12854 19300 12860
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19260 12374 19288 12854
rect 19340 12776 19392 12782
rect 19338 12744 19340 12753
rect 19392 12744 19394 12753
rect 19338 12679 19394 12688
rect 19340 12640 19392 12646
rect 19338 12608 19340 12617
rect 19392 12608 19394 12617
rect 19338 12543 19394 12552
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19260 11762 19288 12038
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19260 10606 19288 11698
rect 19248 10600 19300 10606
rect 19248 10542 19300 10548
rect 19352 10452 19380 12378
rect 19444 11558 19472 13942
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19260 10424 19380 10452
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 19156 8832 19208 8838
rect 19156 8774 19208 8780
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 19168 8430 19196 8774
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 19064 7812 19116 7818
rect 19064 7754 19116 7760
rect 19076 5370 19104 7754
rect 19168 6905 19196 8366
rect 19154 6896 19210 6905
rect 19260 6866 19288 10424
rect 19444 9586 19472 10678
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19352 7342 19380 8910
rect 19444 8566 19472 9318
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 19536 8378 19564 15846
rect 19628 15706 19656 16390
rect 19720 16289 19748 17138
rect 19706 16280 19762 16289
rect 19706 16215 19762 16224
rect 19708 16108 19760 16114
rect 19708 16050 19760 16056
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19720 15586 19748 16050
rect 19628 15558 19748 15586
rect 19628 15502 19656 15558
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19628 10198 19656 15438
rect 19708 15020 19760 15026
rect 19708 14962 19760 14968
rect 19720 14414 19748 14962
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19708 14272 19760 14278
rect 19708 14214 19760 14220
rect 19720 13530 19748 14214
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19720 12186 19748 13262
rect 19812 12481 19840 18702
rect 19892 18148 19944 18154
rect 19892 18090 19944 18096
rect 19904 13326 19932 18090
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 19996 16572 20024 17274
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 20088 16697 20116 16934
rect 20180 16794 20208 19110
rect 20456 18766 20484 19314
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20456 18272 20484 18702
rect 20548 18698 20576 19110
rect 20536 18692 20588 18698
rect 20536 18634 20588 18640
rect 20536 18284 20588 18290
rect 20456 18244 20536 18272
rect 20536 18226 20588 18232
rect 20352 17808 20404 17814
rect 20352 17750 20404 17756
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20168 16788 20220 16794
rect 20168 16730 20220 16736
rect 20074 16688 20130 16697
rect 20074 16623 20130 16632
rect 19996 16544 20116 16572
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19892 13184 19944 13190
rect 19892 13126 19944 13132
rect 19904 12986 19932 13126
rect 19892 12980 19944 12986
rect 19892 12922 19944 12928
rect 19890 12608 19946 12617
rect 19890 12543 19946 12552
rect 19798 12472 19854 12481
rect 19798 12407 19854 12416
rect 19720 12158 19840 12186
rect 19708 12096 19760 12102
rect 19708 12038 19760 12044
rect 19720 11830 19748 12038
rect 19708 11824 19760 11830
rect 19708 11766 19760 11772
rect 19708 11280 19760 11286
rect 19708 11222 19760 11228
rect 19616 10192 19668 10198
rect 19616 10134 19668 10140
rect 19628 9178 19656 10134
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19614 8936 19670 8945
rect 19614 8871 19670 8880
rect 19444 8350 19564 8378
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19154 6831 19210 6840
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19168 6254 19196 6734
rect 19260 6458 19288 6802
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 19154 5128 19210 5137
rect 19154 5063 19210 5072
rect 19168 4060 19196 5063
rect 19352 4842 19380 6938
rect 19444 5001 19472 8350
rect 19628 7818 19656 8871
rect 19720 8634 19748 11222
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19720 7886 19748 8570
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19616 7812 19668 7818
rect 19616 7754 19668 7760
rect 19720 7410 19748 7822
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19524 6928 19576 6934
rect 19524 6870 19576 6876
rect 19536 5710 19564 6870
rect 19812 5914 19840 12158
rect 19904 10674 19932 12543
rect 19892 10668 19944 10674
rect 19892 10610 19944 10616
rect 19904 10305 19932 10610
rect 19890 10296 19946 10305
rect 19890 10231 19946 10240
rect 19892 10124 19944 10130
rect 19892 10066 19944 10072
rect 19904 9654 19932 10066
rect 19892 9648 19944 9654
rect 19892 9590 19944 9596
rect 19890 9344 19946 9353
rect 19890 9279 19946 9288
rect 19904 8838 19932 9279
rect 19996 9042 20024 15846
rect 20088 15065 20116 16544
rect 20168 16448 20220 16454
rect 20168 16390 20220 16396
rect 20074 15056 20130 15065
rect 20074 14991 20130 15000
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 20088 14618 20116 14826
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 20180 14249 20208 16390
rect 20166 14240 20222 14249
rect 20166 14175 20222 14184
rect 20168 13864 20220 13870
rect 20166 13832 20168 13841
rect 20220 13832 20222 13841
rect 20166 13767 20222 13776
rect 20076 13728 20128 13734
rect 20272 13682 20300 17682
rect 20076 13670 20128 13676
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 20088 8090 20116 13670
rect 20180 13654 20300 13682
rect 20180 10266 20208 13654
rect 20364 13546 20392 17750
rect 20548 17678 20576 18226
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20548 17202 20576 17614
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20548 16232 20576 16934
rect 20640 16454 20668 18022
rect 20732 17338 20760 22320
rect 21100 17354 21128 22320
rect 21468 20398 21496 22320
rect 21456 20392 21508 20398
rect 21456 20334 21508 20340
rect 21836 18358 21864 22320
rect 22204 19854 22232 22320
rect 22572 20058 22600 22320
rect 22560 20052 22612 20058
rect 22560 19994 22612 20000
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 21824 18352 21876 18358
rect 21824 18294 21876 18300
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 21008 17326 21128 17354
rect 21272 17332 21324 17338
rect 20902 17096 20958 17105
rect 20902 17031 20958 17040
rect 20628 16448 20680 16454
rect 20628 16390 20680 16396
rect 20548 16204 20760 16232
rect 20444 16176 20496 16182
rect 20548 16153 20576 16204
rect 20444 16118 20496 16124
rect 20534 16144 20590 16153
rect 20456 15570 20484 16118
rect 20534 16079 20590 16088
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20548 15638 20576 15846
rect 20536 15632 20588 15638
rect 20536 15574 20588 15580
rect 20444 15564 20496 15570
rect 20444 15506 20496 15512
rect 20442 15056 20498 15065
rect 20442 14991 20498 15000
rect 20536 15020 20588 15026
rect 20456 13716 20484 14991
rect 20536 14962 20588 14968
rect 20548 13841 20576 14962
rect 20534 13832 20590 13841
rect 20534 13767 20590 13776
rect 20456 13688 20576 13716
rect 20272 13518 20392 13546
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 20180 9897 20208 10202
rect 20166 9888 20222 9897
rect 20166 9823 20222 9832
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 20180 8242 20208 9454
rect 20272 8362 20300 13518
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 20364 12617 20392 13330
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20350 12608 20406 12617
rect 20350 12543 20406 12552
rect 20456 12238 20484 12786
rect 20548 12306 20576 13688
rect 20536 12300 20588 12306
rect 20536 12242 20588 12248
rect 20444 12232 20496 12238
rect 20444 12174 20496 12180
rect 20456 11898 20484 12174
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20536 11552 20588 11558
rect 20536 11494 20588 11500
rect 20548 11354 20576 11494
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20640 11218 20668 16050
rect 20732 13870 20760 16204
rect 20810 15600 20866 15609
rect 20810 15535 20866 15544
rect 20824 14618 20852 15535
rect 20812 14612 20864 14618
rect 20812 14554 20864 14560
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20824 13716 20852 14350
rect 20916 14074 20944 17031
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 20732 13688 20852 13716
rect 20902 13696 20958 13705
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 20444 11008 20496 11014
rect 20444 10950 20496 10956
rect 20456 10606 20484 10950
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 20456 9586 20484 10542
rect 20444 9580 20496 9586
rect 20364 9540 20444 9568
rect 20364 8498 20392 9540
rect 20444 9522 20496 9528
rect 20548 9518 20576 11086
rect 20640 10266 20668 11154
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 20626 10024 20682 10033
rect 20626 9959 20682 9968
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20456 8634 20484 9318
rect 20444 8628 20496 8634
rect 20444 8570 20496 8576
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20260 8356 20312 8362
rect 20260 8298 20312 8304
rect 20180 8214 20300 8242
rect 20076 8084 20128 8090
rect 20076 8026 20128 8032
rect 20076 7948 20128 7954
rect 20076 7890 20128 7896
rect 19890 5944 19946 5953
rect 19800 5908 19852 5914
rect 19890 5879 19946 5888
rect 19800 5850 19852 5856
rect 19904 5846 19932 5879
rect 19892 5840 19944 5846
rect 19892 5782 19944 5788
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 20088 5166 20116 7890
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20180 7546 20208 7822
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 20272 6662 20300 8214
rect 20548 7478 20576 9318
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 20640 7274 20668 9959
rect 20732 9081 20760 13688
rect 20902 13631 20958 13640
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20824 11830 20852 12582
rect 20916 12374 20944 13631
rect 20904 12368 20956 12374
rect 20904 12310 20956 12316
rect 20812 11824 20864 11830
rect 20812 11766 20864 11772
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 20718 9072 20774 9081
rect 20718 9007 20774 9016
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20732 8430 20760 8774
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20628 7268 20680 7274
rect 20628 7210 20680 7216
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20456 6254 20484 7142
rect 20444 6248 20496 6254
rect 20444 6190 20496 6196
rect 20260 6180 20312 6186
rect 20260 6122 20312 6128
rect 20272 5370 20300 6122
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20076 5160 20128 5166
rect 20076 5102 20128 5108
rect 19708 5092 19760 5098
rect 19708 5034 19760 5040
rect 19430 4992 19486 5001
rect 19430 4927 19486 4936
rect 19260 4814 19380 4842
rect 19260 4185 19288 4814
rect 19524 4684 19576 4690
rect 19524 4626 19576 4632
rect 19246 4176 19302 4185
rect 19246 4111 19302 4120
rect 19168 4032 19288 4060
rect 19260 3670 19288 4032
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19248 3664 19300 3670
rect 19248 3606 19300 3612
rect 18786 3567 18842 3576
rect 18972 3596 19024 3602
rect 18972 3538 19024 3544
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 18800 3108 18828 3470
rect 18892 3176 18920 3470
rect 18984 3346 19012 3538
rect 19352 3534 19380 3878
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 18984 3318 19104 3346
rect 18892 3148 19012 3176
rect 18800 3080 18920 3108
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 18708 2446 18736 2994
rect 18788 2576 18840 2582
rect 18788 2518 18840 2524
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 18602 2272 18658 2281
rect 18602 2207 18658 2216
rect 18616 2106 18644 2207
rect 18800 2106 18828 2518
rect 18604 2100 18656 2106
rect 18604 2042 18656 2048
rect 18788 2100 18840 2106
rect 18788 2042 18840 2048
rect 18892 1834 18920 3080
rect 18984 2378 19012 3148
rect 18972 2372 19024 2378
rect 18972 2314 19024 2320
rect 19076 2145 19104 3318
rect 19260 3058 19288 3470
rect 19536 3194 19564 4626
rect 19720 4622 19748 5034
rect 19800 4684 19852 4690
rect 19800 4626 19852 4632
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19708 4616 19760 4622
rect 19708 4558 19760 4564
rect 19628 3466 19656 4558
rect 19720 3942 19748 4558
rect 19812 4078 19840 4626
rect 19892 4616 19944 4622
rect 19892 4558 19944 4564
rect 19800 4072 19852 4078
rect 19800 4014 19852 4020
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19616 3460 19668 3466
rect 19616 3402 19668 3408
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 19246 2952 19302 2961
rect 19246 2887 19302 2896
rect 19430 2952 19486 2961
rect 19430 2887 19486 2896
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 19062 2136 19118 2145
rect 19062 2071 19118 2080
rect 18880 1828 18932 1834
rect 18880 1770 18932 1776
rect 18878 1728 18934 1737
rect 18878 1663 18934 1672
rect 18892 480 18920 1663
rect 19168 1329 19196 2790
rect 19154 1320 19210 1329
rect 19154 1255 19210 1264
rect 19260 480 19288 2887
rect 19444 2106 19472 2887
rect 19720 2650 19748 3334
rect 19904 2990 19932 4558
rect 20168 4548 20220 4554
rect 20168 4490 20220 4496
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 19982 4176 20038 4185
rect 19982 4111 19984 4120
rect 20036 4111 20038 4120
rect 19984 4082 20036 4088
rect 20088 3942 20116 4422
rect 20180 4060 20208 4490
rect 20272 4214 20300 5306
rect 20260 4208 20312 4214
rect 20260 4150 20312 4156
rect 20180 4032 20300 4060
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 19892 2984 19944 2990
rect 19892 2926 19944 2932
rect 19708 2644 19760 2650
rect 19708 2586 19760 2592
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 19432 2100 19484 2106
rect 19432 2042 19484 2048
rect 19904 1902 19932 2450
rect 19996 2446 20024 3878
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20088 3058 20116 3470
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 20272 2666 20300 4032
rect 20352 4004 20404 4010
rect 20352 3946 20404 3952
rect 20364 3777 20392 3946
rect 20350 3768 20406 3777
rect 20350 3703 20406 3712
rect 20352 3664 20404 3670
rect 20350 3632 20352 3641
rect 20404 3632 20406 3641
rect 20350 3567 20406 3576
rect 20272 2638 20392 2666
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 19892 1896 19944 1902
rect 19892 1838 19944 1844
rect 19616 1624 19668 1630
rect 19616 1566 19668 1572
rect 19628 480 19656 1566
rect 19996 480 20024 2246
rect 20364 480 20392 2638
rect 20456 2310 20484 5714
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20548 4282 20576 5102
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20548 2650 20576 4014
rect 20640 3210 20668 5850
rect 20732 3369 20760 8366
rect 20824 6118 20852 11630
rect 20902 11248 20958 11257
rect 20902 11183 20958 11192
rect 20916 9110 20944 11183
rect 21008 10169 21036 17326
rect 21272 17274 21324 17280
rect 21088 17060 21140 17066
rect 21088 17002 21140 17008
rect 20994 10160 21050 10169
rect 20994 10095 21050 10104
rect 20904 9104 20956 9110
rect 20904 9046 20956 9052
rect 20994 8528 21050 8537
rect 20994 8463 21050 8472
rect 20812 6112 20864 6118
rect 20812 6054 20864 6060
rect 20904 4208 20956 4214
rect 20902 4176 20904 4185
rect 20956 4176 20958 4185
rect 20902 4111 20958 4120
rect 20718 3360 20774 3369
rect 20718 3295 20774 3304
rect 20640 3182 20852 3210
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 20536 2644 20588 2650
rect 20536 2586 20588 2592
rect 20640 2582 20668 2790
rect 20628 2576 20680 2582
rect 20628 2518 20680 2524
rect 20444 2304 20496 2310
rect 20824 2281 20852 3182
rect 21008 2972 21036 8463
rect 21100 6866 21128 17002
rect 21178 16280 21234 16289
rect 21178 16215 21234 16224
rect 21192 11898 21220 16215
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21284 11121 21312 17274
rect 21548 17196 21600 17202
rect 21548 17138 21600 17144
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21376 14550 21404 15302
rect 21364 14544 21416 14550
rect 21364 14486 21416 14492
rect 21560 11150 21588 17138
rect 21548 11144 21600 11150
rect 21270 11112 21326 11121
rect 21548 11086 21600 11092
rect 21270 11047 21326 11056
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 21272 5840 21324 5846
rect 21272 5782 21324 5788
rect 21178 3768 21234 3777
rect 21178 3703 21234 3712
rect 20916 2944 21036 2972
rect 20916 2666 20944 2944
rect 21192 2825 21220 3703
rect 21178 2816 21234 2825
rect 21178 2751 21234 2760
rect 20916 2638 21128 2666
rect 20444 2246 20496 2252
rect 20810 2272 20866 2281
rect 20810 2207 20866 2216
rect 20720 1828 20772 1834
rect 20720 1770 20772 1776
rect 20732 480 20760 1770
rect 20824 1737 20852 2207
rect 20810 1728 20866 1737
rect 20810 1663 20866 1672
rect 21100 480 21128 2638
rect 21284 921 21312 5782
rect 21376 2961 21404 8230
rect 21822 4720 21878 4729
rect 21822 4655 21878 4664
rect 21362 2952 21418 2961
rect 21362 2887 21418 2896
rect 21456 1964 21508 1970
rect 21456 1906 21508 1912
rect 21270 912 21326 921
rect 21270 847 21326 856
rect 21468 480 21496 1906
rect 21836 480 21864 4655
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 22204 480 22232 2858
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 22572 480 22600 2790
rect 16486 439 16542 448
rect 16578 0 16634 480
rect 16946 0 17002 480
rect 17406 0 17462 480
rect 17774 0 17830 480
rect 18142 0 18198 480
rect 18510 0 18566 480
rect 18878 0 18934 480
rect 19246 0 19302 480
rect 19614 0 19670 480
rect 19982 0 20038 480
rect 20350 0 20406 480
rect 20718 0 20774 480
rect 21086 0 21142 480
rect 21454 0 21510 480
rect 21822 0 21878 480
rect 22190 0 22246 480
rect 22558 0 22614 480
<< via2 >>
rect 3514 22616 3570 22672
rect 1950 20576 2006 20632
rect 1858 19352 1914 19408
rect 1582 18944 1638 19000
rect 1490 17856 1546 17912
rect 1122 16224 1178 16280
rect 2870 20984 2926 21040
rect 2778 19796 2780 19816
rect 2780 19796 2832 19816
rect 2832 19796 2834 19816
rect 2778 19760 2834 19796
rect 1950 18672 2006 18728
rect 1858 17856 1914 17912
rect 1582 17448 1638 17504
rect 1306 13232 1362 13288
rect 1214 12416 1270 12472
rect 1306 9968 1362 10024
rect 1582 14320 1638 14376
rect 1766 13504 1822 13560
rect 1674 11736 1730 11792
rect 1582 11192 1638 11248
rect 1490 8608 1546 8664
rect 2318 18400 2374 18456
rect 2502 18672 2558 18728
rect 2410 17720 2466 17776
rect 2318 17176 2374 17232
rect 3054 19080 3110 19136
rect 3054 17040 3110 17096
rect 2318 15952 2374 16008
rect 2594 15680 2650 15736
rect 2042 10104 2098 10160
rect 1582 6296 1638 6352
rect 1766 7112 1822 7168
rect 1766 6724 1822 6760
rect 1766 6704 1768 6724
rect 1768 6704 1820 6724
rect 1820 6704 1822 6724
rect 1674 5480 1730 5536
rect 1674 4936 1730 4992
rect 1122 3848 1178 3904
rect 938 3576 994 3632
rect 1122 2896 1178 2952
rect 2594 13776 2650 13832
rect 2870 13096 2926 13152
rect 3146 12280 3202 12336
rect 3054 11872 3110 11928
rect 2778 8472 2834 8528
rect 3422 16652 3478 16688
rect 3422 16632 3424 16652
rect 3424 16632 3476 16652
rect 3476 16632 3478 16652
rect 3330 16496 3386 16552
rect 20626 22616 20682 22672
rect 3882 22208 3938 22264
rect 3698 21800 3754 21856
rect 3606 18264 3662 18320
rect 3698 17992 3754 18048
rect 3790 17584 3846 17640
rect 3606 17040 3662 17096
rect 3698 16768 3754 16824
rect 3422 14728 3478 14784
rect 4066 21412 4122 21448
rect 4066 21392 4068 21412
rect 4068 21392 4120 21412
rect 4120 21392 4122 21412
rect 4066 20204 4068 20224
rect 4068 20204 4120 20224
rect 4120 20204 4122 20224
rect 4066 20168 4122 20204
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4434 18808 4490 18864
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4802 18536 4858 18592
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 5078 19352 5134 19408
rect 4986 18128 5042 18184
rect 4710 17040 4766 17096
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4066 15816 4122 15872
rect 3238 9968 3294 10024
rect 3514 11192 3570 11248
rect 2778 3712 2834 3768
rect 1766 2760 1822 2816
rect 2686 2760 2742 2816
rect 2410 2624 2466 2680
rect 1950 2508 2006 2544
rect 1950 2488 1952 2508
rect 1952 2488 2004 2508
rect 2004 2488 2006 2508
rect 3698 9288 3754 9344
rect 3882 15408 3938 15464
rect 3974 15136 4030 15192
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4894 15544 4950 15600
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4250 13912 4306 13968
rect 3882 11600 3938 11656
rect 3698 9016 3754 9072
rect 3422 6704 3478 6760
rect 3606 6704 3662 6760
rect 3422 5752 3478 5808
rect 3238 3168 3294 3224
rect 2962 2080 3018 2136
rect 3054 1672 3110 1728
rect 3698 3984 3754 4040
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4066 12688 4122 12744
rect 5078 14728 5134 14784
rect 5630 19080 5686 19136
rect 5262 17856 5318 17912
rect 5538 17620 5540 17640
rect 5540 17620 5592 17640
rect 5592 17620 5594 17640
rect 5538 17584 5594 17620
rect 6366 18944 6422 19000
rect 6366 17992 6422 18048
rect 6366 17584 6422 17640
rect 5354 15272 5410 15328
rect 5262 15156 5318 15192
rect 5262 15136 5264 15156
rect 5264 15136 5316 15156
rect 5316 15136 5318 15156
rect 5354 14320 5410 14376
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4894 11636 4896 11656
rect 4896 11636 4948 11656
rect 4948 11636 4950 11656
rect 4894 11600 4950 11636
rect 4802 11464 4858 11520
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4894 10240 4950 10296
rect 4802 9424 4858 9480
rect 4710 8880 4766 8936
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4250 8608 4306 8664
rect 3974 7656 4030 7712
rect 3974 6604 3976 6624
rect 3976 6604 4028 6624
rect 4028 6604 4030 6624
rect 3974 6568 4030 6604
rect 4434 7792 4490 7848
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 5078 9560 5134 9616
rect 4986 8608 5042 8664
rect 4710 7384 4766 7440
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4250 6452 4306 6488
rect 4250 6432 4252 6452
rect 4252 6432 4304 6452
rect 4304 6432 4306 6452
rect 4710 5888 4766 5944
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 5354 11872 5410 11928
rect 5538 10920 5594 10976
rect 5354 10648 5410 10704
rect 5170 9288 5226 9344
rect 5170 7656 5226 7712
rect 5078 6160 5134 6216
rect 4986 5616 5042 5672
rect 4894 5480 4950 5536
rect 4802 4936 4858 4992
rect 4986 4936 5042 4992
rect 3790 3848 3846 3904
rect 3882 3168 3938 3224
rect 3790 3032 3846 3088
rect 3698 2896 3754 2952
rect 3698 1808 3754 1864
rect 3606 856 3662 912
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4342 4120 4398 4176
rect 4158 3460 4214 3496
rect 4158 3440 4160 3460
rect 4160 3440 4212 3460
rect 4212 3440 4214 3460
rect 4342 3440 4398 3496
rect 4250 3304 4306 3360
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4250 2760 4306 2816
rect 4158 2488 4214 2544
rect 4158 1264 4214 1320
rect 4342 2372 4398 2408
rect 4342 2352 4344 2372
rect 4344 2352 4396 2372
rect 4396 2352 4398 2372
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 5354 8880 5410 8936
rect 5262 5208 5318 5264
rect 5262 3712 5318 3768
rect 5078 3440 5134 3496
rect 5630 10648 5686 10704
rect 5446 6568 5502 6624
rect 5446 5480 5502 5536
rect 5538 5344 5594 5400
rect 5906 15680 5962 15736
rect 6458 15680 6514 15736
rect 6090 14048 6146 14104
rect 6182 13912 6238 13968
rect 5906 12688 5962 12744
rect 5906 11736 5962 11792
rect 5906 10412 5908 10432
rect 5908 10412 5960 10432
rect 5960 10412 5962 10432
rect 5906 10376 5962 10412
rect 6090 10648 6146 10704
rect 6090 10240 6146 10296
rect 6366 13368 6422 13424
rect 6826 18264 6882 18320
rect 6734 17856 6790 17912
rect 6642 15408 6698 15464
rect 6734 13640 6790 13696
rect 6458 11192 6514 11248
rect 6274 9424 6330 9480
rect 6182 7928 6238 7984
rect 6642 11872 6698 11928
rect 6642 9560 6698 9616
rect 6458 8200 6514 8256
rect 6458 7928 6514 7984
rect 6182 7520 6238 7576
rect 6366 7248 6422 7304
rect 5722 6432 5778 6488
rect 5722 6160 5778 6216
rect 5446 4256 5502 4312
rect 5538 3984 5594 4040
rect 5354 3032 5410 3088
rect 6642 6976 6698 7032
rect 7378 22208 7434 22264
rect 7194 17992 7250 18048
rect 7286 17448 7342 17504
rect 7010 12552 7066 12608
rect 7286 15000 7342 15056
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7470 15680 7526 15736
rect 7562 14456 7618 14512
rect 8298 19896 8354 19952
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 8206 18944 8262 19000
rect 7746 18536 7802 18592
rect 8022 18400 8078 18456
rect 8482 18672 8538 18728
rect 8666 19488 8722 19544
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 8022 17040 8078 17096
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7930 15272 7986 15328
rect 7746 15000 7802 15056
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7930 14476 7986 14512
rect 7930 14456 7932 14476
rect 7932 14456 7984 14476
rect 7984 14456 7986 14476
rect 8114 14048 8170 14104
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7102 12280 7158 12336
rect 6826 10240 6882 10296
rect 7010 10240 7066 10296
rect 6642 6060 6644 6080
rect 6644 6060 6696 6080
rect 6696 6060 6698 6080
rect 6642 6024 6698 6060
rect 6550 5888 6606 5944
rect 5998 4256 6054 4312
rect 5998 4004 6054 4040
rect 5998 3984 6000 4004
rect 6000 3984 6052 4004
rect 6052 3984 6054 4004
rect 6458 3440 6514 3496
rect 6366 1944 6422 2000
rect 6826 5888 6882 5944
rect 7286 12688 7342 12744
rect 7378 12436 7434 12472
rect 7378 12416 7380 12436
rect 7380 12416 7432 12436
rect 7432 12416 7434 12436
rect 7654 12280 7710 12336
rect 7470 12008 7526 12064
rect 7194 9016 7250 9072
rect 7470 9988 7526 10024
rect 7470 9968 7472 9988
rect 7472 9968 7524 9988
rect 7524 9968 7526 9988
rect 7470 9560 7526 9616
rect 7470 8608 7526 8664
rect 7286 7384 7342 7440
rect 7194 5888 7250 5944
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7930 12280 7986 12336
rect 8298 17856 8354 17912
rect 8666 17992 8722 18048
rect 8482 16088 8538 16144
rect 8482 15136 8538 15192
rect 8850 19080 8906 19136
rect 8850 18400 8906 18456
rect 9218 19352 9274 19408
rect 9034 17856 9090 17912
rect 8850 15952 8906 16008
rect 8758 15816 8814 15872
rect 8942 13232 8998 13288
rect 8298 11736 8354 11792
rect 7838 11636 7840 11656
rect 7840 11636 7892 11656
rect 7892 11636 7894 11656
rect 7838 11600 7894 11636
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 8574 12044 8576 12064
rect 8576 12044 8628 12064
rect 8628 12044 8630 12064
rect 8574 12008 8630 12044
rect 7746 11056 7802 11112
rect 8206 11056 8262 11112
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 8390 10376 8446 10432
rect 7838 10104 7894 10160
rect 8022 9424 8078 9480
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 8390 9152 8446 9208
rect 8298 8608 8354 8664
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 8666 10376 8722 10432
rect 8574 10240 8630 10296
rect 9034 12280 9090 12336
rect 8850 11328 8906 11384
rect 8942 11192 8998 11248
rect 8850 10648 8906 10704
rect 8574 8608 8630 8664
rect 7654 7792 7710 7848
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 6182 1536 6238 1592
rect 3974 176 4030 232
rect 6090 448 6146 504
rect 7378 3612 7380 3632
rect 7380 3612 7432 3632
rect 7432 3612 7434 3632
rect 7010 3304 7066 3360
rect 7378 3576 7434 3612
rect 7654 6432 7710 6488
rect 7930 6296 7986 6352
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7838 5072 7894 5128
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7470 3168 7526 3224
rect 7102 2624 7158 2680
rect 7378 2080 7434 2136
rect 7286 1672 7342 1728
rect 9034 10376 9090 10432
rect 9402 18400 9458 18456
rect 9678 18808 9734 18864
rect 9770 18400 9826 18456
rect 9494 17448 9550 17504
rect 9862 17856 9918 17912
rect 9678 16904 9734 16960
rect 9678 15700 9734 15736
rect 9678 15680 9680 15700
rect 9680 15680 9732 15700
rect 9732 15680 9734 15700
rect 9402 13640 9458 13696
rect 9310 12416 9366 12472
rect 9310 12144 9366 12200
rect 9586 12416 9642 12472
rect 10138 18264 10194 18320
rect 10046 16768 10102 16824
rect 9402 11328 9458 11384
rect 9218 10784 9274 10840
rect 9218 10512 9274 10568
rect 9402 10376 9458 10432
rect 8942 9424 8998 9480
rect 9034 8744 9090 8800
rect 8574 6316 8630 6352
rect 8574 6296 8576 6316
rect 8576 6296 8628 6316
rect 8628 6296 8630 6316
rect 8574 6180 8630 6216
rect 8574 6160 8576 6180
rect 8576 6160 8628 6180
rect 8628 6160 8630 6180
rect 8574 5908 8630 5944
rect 8574 5888 8576 5908
rect 8576 5888 8628 5908
rect 8628 5888 8630 5908
rect 8574 4392 8630 4448
rect 8298 3168 8354 3224
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 8482 3440 8538 3496
rect 8022 1536 8078 1592
rect 8850 7520 8906 7576
rect 8850 7248 8906 7304
rect 8850 4936 8906 4992
rect 9310 7792 9366 7848
rect 9494 8064 9550 8120
rect 9954 12416 10010 12472
rect 10322 16632 10378 16688
rect 10322 13252 10378 13288
rect 10322 13232 10324 13252
rect 10324 13232 10376 13252
rect 10376 13232 10378 13252
rect 10782 19488 10838 19544
rect 10874 19352 10930 19408
rect 10690 18536 10746 18592
rect 10782 18400 10838 18456
rect 10782 18264 10838 18320
rect 10690 16904 10746 16960
rect 10690 16396 10692 16416
rect 10692 16396 10744 16416
rect 10744 16396 10746 16416
rect 10690 16360 10746 16396
rect 10506 12980 10562 13016
rect 10506 12960 10508 12980
rect 10508 12960 10560 12980
rect 10560 12960 10562 12980
rect 10138 12416 10194 12472
rect 10046 12144 10102 12200
rect 10046 11600 10102 11656
rect 9862 9696 9918 9752
rect 9402 7520 9458 7576
rect 9402 6296 9458 6352
rect 8850 4120 8906 4176
rect 8850 3032 8906 3088
rect 9126 3304 9182 3360
rect 9586 6024 9642 6080
rect 9402 5344 9458 5400
rect 10138 10784 10194 10840
rect 9678 5072 9734 5128
rect 9862 5072 9918 5128
rect 10138 4664 10194 4720
rect 10414 12280 10470 12336
rect 11058 19760 11114 19816
rect 11058 18944 11114 19000
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 12254 19896 12310 19952
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11978 18148 12034 18184
rect 11978 18128 11980 18148
rect 11980 18128 12032 18148
rect 12032 18128 12034 18148
rect 12162 18128 12218 18184
rect 11794 17856 11850 17912
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 10598 11736 10654 11792
rect 10782 12824 10838 12880
rect 10874 12552 10930 12608
rect 12438 19508 12494 19544
rect 12438 19488 12440 19508
rect 12440 19488 12492 19508
rect 12492 19488 12494 19508
rect 12162 17720 12218 17776
rect 12070 17584 12126 17640
rect 11978 17040 12034 17096
rect 12070 16632 12126 16688
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11150 15680 11206 15736
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11518 15000 11574 15056
rect 11426 14456 11482 14512
rect 12254 15308 12256 15328
rect 12256 15308 12308 15328
rect 12308 15308 12310 15328
rect 12254 15272 12310 15308
rect 12622 17040 12678 17096
rect 12438 16088 12494 16144
rect 12438 15680 12494 15736
rect 11518 14356 11520 14376
rect 11520 14356 11572 14376
rect 11572 14356 11574 14376
rect 11518 14320 11574 14356
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11426 13912 11482 13968
rect 11518 13524 11574 13560
rect 11518 13504 11520 13524
rect 11520 13504 11572 13524
rect 11572 13504 11574 13524
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11150 12416 11206 12472
rect 10966 12144 11022 12200
rect 10598 11464 10654 11520
rect 10690 10920 10746 10976
rect 10598 9832 10654 9888
rect 10506 9696 10562 9752
rect 10414 9424 10470 9480
rect 10506 9288 10562 9344
rect 10598 9152 10654 9208
rect 10690 8200 10746 8256
rect 10322 7520 10378 7576
rect 9310 3168 9366 3224
rect 9126 2760 9182 2816
rect 9126 2216 9182 2272
rect 10506 6024 10562 6080
rect 9770 2760 9826 2816
rect 10230 2896 10286 2952
rect 10322 2644 10378 2680
rect 10322 2624 10324 2644
rect 10324 2624 10376 2644
rect 10376 2624 10378 2644
rect 11702 12008 11758 12064
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11978 14456 12034 14512
rect 11886 12552 11942 12608
rect 12254 14320 12310 14376
rect 12254 13640 12310 13696
rect 12070 12416 12126 12472
rect 11886 12280 11942 12336
rect 12070 12280 12126 12336
rect 12254 12280 12310 12336
rect 11978 12144 12034 12200
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11794 11736 11850 11792
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11150 9152 11206 9208
rect 11518 9560 11574 9616
rect 11610 9288 11666 9344
rect 11334 8880 11390 8936
rect 11518 8880 11574 8936
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11150 8336 11206 8392
rect 11058 8064 11114 8120
rect 10966 7520 11022 7576
rect 11058 7384 11114 7440
rect 11242 7792 11298 7848
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11150 7248 11206 7304
rect 11518 7248 11574 7304
rect 11242 6840 11298 6896
rect 11058 6568 11114 6624
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 10782 6024 10838 6080
rect 10966 5072 11022 5128
rect 10690 4936 10746 4992
rect 10690 3304 10746 3360
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 12162 12008 12218 12064
rect 12070 10784 12126 10840
rect 12254 11736 12310 11792
rect 12254 11328 12310 11384
rect 12530 14184 12586 14240
rect 12438 14048 12494 14104
rect 12714 16088 12770 16144
rect 13174 17040 13230 17096
rect 12714 12960 12770 13016
rect 12530 11736 12586 11792
rect 12070 9868 12072 9888
rect 12072 9868 12124 9888
rect 12124 9868 12126 9888
rect 12070 9832 12126 9868
rect 11794 8880 11850 8936
rect 11794 8744 11850 8800
rect 11702 5072 11758 5128
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11978 9596 11980 9616
rect 11980 9596 12032 9616
rect 12032 9596 12034 9616
rect 11978 9560 12034 9596
rect 11978 8608 12034 8664
rect 11978 8336 12034 8392
rect 12622 11348 12678 11384
rect 12622 11328 12624 11348
rect 12624 11328 12676 11348
rect 12676 11328 12678 11348
rect 13082 14456 13138 14512
rect 12990 12280 13046 12336
rect 13174 13368 13230 13424
rect 13542 15680 13598 15736
rect 13358 13368 13414 13424
rect 13358 12824 13414 12880
rect 13726 13096 13782 13152
rect 13634 12824 13690 12880
rect 12990 11872 13046 11928
rect 12254 9696 12310 9752
rect 12438 10784 12494 10840
rect 12254 8608 12310 8664
rect 12622 8880 12678 8936
rect 12070 7248 12126 7304
rect 11886 6432 11942 6488
rect 11978 3984 12034 4040
rect 10966 3440 11022 3496
rect 11058 3304 11114 3360
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 11978 3576 12034 3632
rect 11794 3168 11850 3224
rect 11794 2760 11850 2816
rect 12806 11056 12862 11112
rect 12806 8336 12862 8392
rect 12438 6024 12494 6080
rect 12622 5888 12678 5944
rect 12438 5616 12494 5672
rect 12346 4936 12402 4992
rect 12622 4936 12678 4992
rect 12622 4004 12678 4040
rect 12622 3984 12624 4004
rect 12624 3984 12676 4004
rect 12676 3984 12678 4004
rect 12530 3440 12586 3496
rect 12990 10920 13046 10976
rect 12990 8744 13046 8800
rect 13082 7520 13138 7576
rect 12990 7248 13046 7304
rect 12898 6976 12954 7032
rect 12898 6876 12900 6896
rect 12900 6876 12952 6896
rect 12952 6876 12954 6896
rect 12898 6840 12954 6876
rect 13450 12280 13506 12336
rect 13358 11872 13414 11928
rect 13542 11192 13598 11248
rect 14186 19352 14242 19408
rect 14370 19080 14426 19136
rect 14002 18128 14058 18184
rect 14094 16904 14150 16960
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14554 18400 14610 18456
rect 14094 15680 14150 15736
rect 14094 15020 14150 15056
rect 14094 15000 14096 15020
rect 14096 15000 14148 15020
rect 14148 15000 14150 15020
rect 13542 10376 13598 10432
rect 13542 9968 13598 10024
rect 13450 9152 13506 9208
rect 13082 5752 13138 5808
rect 13082 5072 13138 5128
rect 13082 4800 13138 4856
rect 12806 4392 12862 4448
rect 12806 3712 12862 3768
rect 13358 5480 13414 5536
rect 13266 5344 13322 5400
rect 13266 4528 13322 4584
rect 13082 3848 13138 3904
rect 13266 3032 13322 3088
rect 12990 2760 13046 2816
rect 13082 2488 13138 2544
rect 14186 12416 14242 12472
rect 14186 11328 14242 11384
rect 14002 11192 14058 11248
rect 13910 11092 13912 11112
rect 13912 11092 13964 11112
rect 13964 11092 13966 11112
rect 13910 11056 13966 11092
rect 14002 10920 14058 10976
rect 13726 8472 13782 8528
rect 13910 9424 13966 9480
rect 14186 10920 14242 10976
rect 13910 8064 13966 8120
rect 13726 7656 13782 7712
rect 13634 6976 13690 7032
rect 14370 11328 14426 11384
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 15474 19352 15530 19408
rect 15382 18808 15438 18864
rect 15290 18400 15346 18456
rect 15198 17856 15254 17912
rect 15106 17720 15162 17776
rect 15014 17448 15070 17504
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14554 16632 14610 16688
rect 15198 16360 15254 16416
rect 15106 15816 15162 15872
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 15106 15680 15162 15736
rect 15014 15544 15070 15600
rect 15014 15000 15070 15056
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14646 14456 14702 14512
rect 14646 13812 14648 13832
rect 14648 13812 14700 13832
rect 14700 13812 14702 13832
rect 14646 13776 14702 13812
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14646 13096 14702 13152
rect 14830 13096 14886 13152
rect 14554 12688 14610 12744
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14554 12144 14610 12200
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14554 11056 14610 11112
rect 14462 10376 14518 10432
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14922 9560 14978 9616
rect 14370 9152 14426 9208
rect 14278 8200 14334 8256
rect 14094 7520 14150 7576
rect 13910 6024 13966 6080
rect 13634 4392 13690 4448
rect 14094 6296 14150 6352
rect 14002 5480 14058 5536
rect 13910 5344 13966 5400
rect 14094 4972 14096 4992
rect 14096 4972 14148 4992
rect 14148 4972 14150 4992
rect 14094 4936 14150 4972
rect 14094 4800 14150 4856
rect 13910 4120 13966 4176
rect 13818 3984 13874 4040
rect 13818 3712 13874 3768
rect 13634 1944 13690 2000
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 15198 14456 15254 14512
rect 15198 13912 15254 13968
rect 15198 12144 15254 12200
rect 15106 11500 15108 11520
rect 15108 11500 15160 11520
rect 15160 11500 15162 11520
rect 15106 11464 15162 11500
rect 15566 15444 15568 15464
rect 15568 15444 15620 15464
rect 15620 15444 15622 15464
rect 15566 15408 15622 15444
rect 16118 18400 16174 18456
rect 16026 17992 16082 18048
rect 16026 17620 16028 17640
rect 16028 17620 16080 17640
rect 16080 17620 16082 17640
rect 16026 17584 16082 17620
rect 15842 17448 15898 17504
rect 16026 16768 16082 16824
rect 15750 15544 15806 15600
rect 15842 15408 15898 15464
rect 15658 15136 15714 15192
rect 15382 15020 15438 15056
rect 15382 15000 15384 15020
rect 15384 15000 15436 15020
rect 15436 15000 15438 15020
rect 15474 14900 15476 14920
rect 15476 14900 15528 14920
rect 15528 14900 15530 14920
rect 15474 14864 15530 14900
rect 15566 14048 15622 14104
rect 15474 12552 15530 12608
rect 15474 12416 15530 12472
rect 15474 11736 15530 11792
rect 15566 11328 15622 11384
rect 15658 11056 15714 11112
rect 15382 10376 15438 10432
rect 15198 9172 15254 9208
rect 15198 9152 15200 9172
rect 15200 9152 15252 9172
rect 15252 9152 15254 9172
rect 14646 8472 14702 8528
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 16302 19488 16358 19544
rect 16394 18536 16450 18592
rect 16486 18128 16542 18184
rect 16210 16360 16266 16416
rect 16118 16088 16174 16144
rect 16026 15136 16082 15192
rect 15934 13504 15990 13560
rect 16026 12552 16082 12608
rect 15842 11892 15898 11928
rect 15842 11872 15844 11892
rect 15844 11872 15896 11892
rect 15896 11872 15898 11892
rect 16302 15000 16358 15056
rect 16302 13912 16358 13968
rect 16762 19624 16818 19680
rect 16486 14456 16542 14512
rect 16394 13232 16450 13288
rect 16210 12688 16266 12744
rect 16118 12416 16174 12472
rect 17038 18264 17094 18320
rect 17498 19760 17554 19816
rect 17590 19624 17646 19680
rect 17222 18808 17278 18864
rect 17222 17992 17278 18048
rect 17222 16904 17278 16960
rect 17038 16632 17094 16688
rect 16394 12552 16450 12608
rect 16302 12416 16358 12472
rect 16118 11464 16174 11520
rect 15658 10104 15714 10160
rect 15566 9288 15622 9344
rect 15566 9052 15568 9072
rect 15568 9052 15620 9072
rect 15620 9052 15622 9072
rect 15566 9016 15622 9052
rect 15566 8744 15622 8800
rect 15842 9580 15898 9616
rect 15842 9560 15844 9580
rect 15844 9560 15896 9580
rect 15896 9560 15898 9580
rect 15750 9016 15806 9072
rect 14370 7112 14426 7168
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14922 6568 14978 6624
rect 15106 6604 15108 6624
rect 15108 6604 15160 6624
rect 15160 6604 15162 6624
rect 15106 6568 15162 6604
rect 15290 7148 15292 7168
rect 15292 7148 15344 7168
rect 15344 7148 15346 7168
rect 15290 7112 15346 7148
rect 15198 6432 15254 6488
rect 14922 6296 14978 6352
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14738 4256 14794 4312
rect 14462 3848 14518 3904
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14830 3596 14886 3632
rect 14830 3576 14832 3596
rect 14832 3576 14884 3596
rect 14884 3576 14886 3596
rect 14462 3168 14518 3224
rect 14462 2372 14518 2408
rect 14462 2352 14464 2372
rect 14464 2352 14516 2372
rect 14516 2352 14518 2372
rect 14922 3052 14978 3088
rect 14922 3032 14924 3052
rect 14924 3032 14976 3052
rect 14976 3032 14978 3052
rect 14738 2916 14794 2952
rect 15106 4800 15162 4856
rect 15198 3984 15254 4040
rect 15474 5208 15530 5264
rect 15474 4120 15530 4176
rect 15106 3712 15162 3768
rect 15382 3848 15438 3904
rect 15198 3576 15254 3632
rect 14738 2896 14740 2916
rect 14740 2896 14792 2916
rect 14792 2896 14794 2916
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 15382 3168 15438 3224
rect 15382 2896 15438 2952
rect 15382 2216 15438 2272
rect 15750 7520 15806 7576
rect 15842 7248 15898 7304
rect 15658 3984 15714 4040
rect 15842 5616 15898 5672
rect 15842 5208 15898 5264
rect 16394 11872 16450 11928
rect 16578 11736 16634 11792
rect 16578 11600 16634 11656
rect 16486 11464 16542 11520
rect 16394 11328 16450 11384
rect 16302 10532 16358 10568
rect 16302 10512 16304 10532
rect 16304 10512 16356 10532
rect 16356 10512 16358 10532
rect 16210 10104 16266 10160
rect 16026 9560 16082 9616
rect 16118 9424 16174 9480
rect 16394 9560 16450 9616
rect 16302 9444 16358 9480
rect 16302 9424 16304 9444
rect 16304 9424 16356 9444
rect 16356 9424 16358 9444
rect 16394 9288 16450 9344
rect 16302 8744 16358 8800
rect 16210 7148 16212 7168
rect 16212 7148 16264 7168
rect 16264 7148 16266 7168
rect 16210 7112 16266 7148
rect 16578 9152 16634 9208
rect 16486 9016 16542 9072
rect 16486 8472 16542 8528
rect 16210 6704 16266 6760
rect 16578 7928 16634 7984
rect 16486 6704 16542 6760
rect 16578 5344 16634 5400
rect 16946 14320 17002 14376
rect 17038 13504 17094 13560
rect 16854 13096 16910 13152
rect 17314 16668 17316 16688
rect 17316 16668 17368 16688
rect 17368 16668 17370 16688
rect 17314 16632 17370 16668
rect 17498 19252 17500 19272
rect 17500 19252 17552 19272
rect 17552 19252 17554 19272
rect 17498 19216 17554 19252
rect 17590 19080 17646 19136
rect 17958 20984 18014 21040
rect 18142 21392 18198 21448
rect 18786 20576 18842 20632
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 17682 18808 17738 18864
rect 17682 18128 17738 18184
rect 17590 17720 17646 17776
rect 17590 16632 17646 16688
rect 17958 18808 18014 18864
rect 18142 18672 18198 18728
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 17958 18300 17960 18320
rect 17960 18300 18012 18320
rect 18012 18300 18014 18320
rect 17958 18264 18014 18300
rect 18602 18672 18658 18728
rect 17866 17312 17922 17368
rect 18418 18028 18420 18048
rect 18420 18028 18472 18048
rect 18472 18028 18474 18048
rect 18418 17992 18474 18028
rect 18050 17856 18106 17912
rect 18234 17856 18290 17912
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 17958 17176 18014 17232
rect 18602 17040 18658 17096
rect 17774 16088 17830 16144
rect 17590 14728 17646 14784
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 17866 15544 17922 15600
rect 16762 11872 16818 11928
rect 16762 10920 16818 10976
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18602 15952 18658 16008
rect 18602 15680 18658 15736
rect 18142 14728 18198 14784
rect 17682 14320 17738 14376
rect 17682 13912 17738 13968
rect 17590 12824 17646 12880
rect 16946 11736 17002 11792
rect 16762 8608 16818 8664
rect 18234 14476 18290 14512
rect 18234 14456 18236 14476
rect 18236 14456 18288 14476
rect 18288 14456 18290 14476
rect 18418 14884 18474 14920
rect 18418 14864 18420 14884
rect 18420 14864 18472 14884
rect 18472 14864 18474 14884
rect 18510 14456 18566 14512
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18050 13776 18106 13832
rect 18418 13504 18474 13560
rect 18234 13368 18290 13424
rect 18878 19760 18934 19816
rect 18878 17448 18934 17504
rect 18878 17040 18934 17096
rect 19246 22208 19302 22264
rect 19154 18944 19210 19000
rect 19154 18164 19156 18184
rect 19156 18164 19208 18184
rect 19208 18164 19210 18184
rect 19154 18128 19210 18164
rect 19154 18028 19156 18048
rect 19156 18028 19208 18048
rect 19208 18028 19210 18048
rect 19154 17992 19210 18028
rect 18694 13640 18750 13696
rect 18970 15580 18972 15600
rect 18972 15580 19024 15600
rect 19024 15580 19026 15600
rect 18970 15544 19026 15580
rect 18878 14864 18934 14920
rect 18878 14728 18934 14784
rect 18878 13504 18934 13560
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 17866 12008 17922 12064
rect 17774 11892 17830 11928
rect 17774 11872 17776 11892
rect 17776 11872 17828 11892
rect 17828 11872 17830 11892
rect 17774 11736 17830 11792
rect 17682 11600 17738 11656
rect 17314 10532 17370 10568
rect 17314 10512 17316 10532
rect 17316 10512 17368 10532
rect 17368 10512 17370 10532
rect 17314 10240 17370 10296
rect 17222 10004 17224 10024
rect 17224 10004 17276 10024
rect 17276 10004 17278 10024
rect 17222 9968 17278 10004
rect 17222 9560 17278 9616
rect 17038 9424 17094 9480
rect 16946 9288 17002 9344
rect 16762 8336 16818 8392
rect 16854 7792 16910 7848
rect 16302 1944 16358 2000
rect 17038 5888 17094 5944
rect 16946 4120 17002 4176
rect 16946 3984 17002 4040
rect 17590 9560 17646 9616
rect 17406 8064 17462 8120
rect 17314 6568 17370 6624
rect 18418 12144 18474 12200
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 17958 11464 18014 11520
rect 17866 11328 17922 11384
rect 17866 10376 17922 10432
rect 18142 11228 18144 11248
rect 18144 11228 18196 11248
rect 18196 11228 18198 11248
rect 18142 11192 18198 11228
rect 18602 13096 18658 13152
rect 18786 13096 18842 13152
rect 18786 12688 18842 12744
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18418 10648 18474 10704
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 17958 9036 18014 9072
rect 17958 9016 17960 9036
rect 17960 9016 18012 9036
rect 18012 9016 18014 9036
rect 18694 12008 18750 12064
rect 18326 9036 18382 9072
rect 18326 9016 18328 9036
rect 18328 9016 18380 9036
rect 18380 9016 18382 9036
rect 18510 9016 18566 9072
rect 18510 8744 18566 8800
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 19062 12724 19064 12744
rect 19064 12724 19116 12744
rect 19116 12724 19118 12744
rect 19062 12688 19118 12724
rect 19062 12552 19118 12608
rect 18878 11464 18934 11520
rect 19062 11328 19118 11384
rect 18694 8200 18750 8256
rect 18786 8064 18842 8120
rect 17682 5888 17738 5944
rect 17498 4936 17554 4992
rect 16854 2524 16856 2544
rect 16856 2524 16908 2544
rect 16908 2524 16910 2544
rect 16854 2488 16910 2524
rect 16486 448 16542 504
rect 17130 2644 17186 2680
rect 17130 2624 17132 2644
rect 17132 2624 17184 2644
rect 17184 2624 17186 2644
rect 18234 7384 18290 7440
rect 18326 6996 18382 7032
rect 18326 6976 18328 6996
rect 18328 6976 18380 6996
rect 18380 6976 18382 6996
rect 18510 6840 18566 6896
rect 18326 6740 18328 6760
rect 18328 6740 18380 6760
rect 18380 6740 18382 6760
rect 18326 6704 18382 6740
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18142 5888 18198 5944
rect 18326 5772 18382 5808
rect 18326 5752 18328 5772
rect 18328 5752 18380 5772
rect 18380 5752 18382 5772
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 17682 2352 17738 2408
rect 18050 4140 18106 4176
rect 18050 4120 18052 4140
rect 18052 4120 18104 4140
rect 18104 4120 18106 4140
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 18786 7112 18842 7168
rect 18878 4120 18934 4176
rect 18786 3576 18842 3632
rect 19246 16632 19302 16688
rect 19246 15816 19302 15872
rect 19522 17584 19578 17640
rect 19890 21800 19946 21856
rect 20350 20168 20406 20224
rect 19522 16632 19578 16688
rect 19430 15272 19486 15328
rect 19430 15156 19486 15192
rect 19430 15136 19432 15156
rect 19432 15136 19484 15156
rect 19484 15136 19486 15156
rect 19338 14592 19394 14648
rect 19338 14456 19394 14512
rect 19430 14184 19486 14240
rect 19246 13504 19302 13560
rect 19246 12960 19302 13016
rect 19338 12724 19340 12744
rect 19340 12724 19392 12744
rect 19392 12724 19394 12744
rect 19338 12688 19394 12724
rect 19338 12588 19340 12608
rect 19340 12588 19392 12608
rect 19392 12588 19394 12608
rect 19338 12552 19394 12588
rect 19154 6840 19210 6896
rect 19706 16224 19762 16280
rect 20074 16632 20130 16688
rect 19890 12552 19946 12608
rect 19798 12416 19854 12472
rect 19614 8880 19670 8936
rect 19154 5072 19210 5128
rect 19890 10240 19946 10296
rect 19890 9288 19946 9344
rect 20074 15000 20130 15056
rect 20166 14184 20222 14240
rect 20166 13812 20168 13832
rect 20168 13812 20220 13832
rect 20220 13812 20222 13832
rect 20166 13776 20222 13812
rect 20902 17040 20958 17096
rect 20534 16088 20590 16144
rect 20442 15000 20498 15056
rect 20534 13776 20590 13832
rect 20166 9832 20222 9888
rect 20350 12552 20406 12608
rect 20810 15544 20866 15600
rect 20626 9968 20682 10024
rect 19890 5888 19946 5944
rect 20902 13640 20958 13696
rect 20718 9016 20774 9072
rect 19430 4936 19486 4992
rect 19246 4120 19302 4176
rect 18602 2216 18658 2272
rect 19246 2896 19302 2952
rect 19430 2896 19486 2952
rect 19062 2080 19118 2136
rect 18878 1672 18934 1728
rect 19154 1264 19210 1320
rect 19982 4140 20038 4176
rect 19982 4120 19984 4140
rect 19984 4120 20036 4140
rect 20036 4120 20038 4140
rect 20350 3712 20406 3768
rect 20350 3612 20352 3632
rect 20352 3612 20404 3632
rect 20404 3612 20406 3632
rect 20350 3576 20406 3612
rect 20902 11192 20958 11248
rect 20994 10104 21050 10160
rect 20994 8472 21050 8528
rect 20902 4156 20904 4176
rect 20904 4156 20956 4176
rect 20956 4156 20958 4176
rect 20902 4120 20958 4156
rect 20718 3304 20774 3360
rect 21178 16224 21234 16280
rect 21270 11056 21326 11112
rect 21178 3712 21234 3768
rect 21178 2760 21234 2816
rect 20810 2216 20866 2272
rect 20810 1672 20866 1728
rect 21822 4664 21878 4720
rect 21362 2896 21418 2952
rect 21270 856 21326 912
<< metal3 >>
rect 0 22674 480 22704
rect 3509 22674 3575 22677
rect 0 22672 3575 22674
rect 0 22616 3514 22672
rect 3570 22616 3575 22672
rect 0 22614 3575 22616
rect 0 22584 480 22614
rect 3509 22611 3575 22614
rect 20621 22674 20687 22677
rect 22320 22674 22800 22704
rect 20621 22672 22800 22674
rect 20621 22616 20626 22672
rect 20682 22616 22800 22672
rect 20621 22614 22800 22616
rect 20621 22611 20687 22614
rect 22320 22584 22800 22614
rect 0 22266 480 22296
rect 3877 22266 3943 22269
rect 0 22264 3943 22266
rect 0 22208 3882 22264
rect 3938 22208 3943 22264
rect 0 22206 3943 22208
rect 0 22176 480 22206
rect 3877 22203 3943 22206
rect 7046 22204 7052 22268
rect 7116 22266 7122 22268
rect 7373 22266 7439 22269
rect 7116 22264 7439 22266
rect 7116 22208 7378 22264
rect 7434 22208 7439 22264
rect 7116 22206 7439 22208
rect 7116 22204 7122 22206
rect 7373 22203 7439 22206
rect 19241 22266 19307 22269
rect 22320 22266 22800 22296
rect 19241 22264 22800 22266
rect 19241 22208 19246 22264
rect 19302 22208 22800 22264
rect 19241 22206 22800 22208
rect 19241 22203 19307 22206
rect 22320 22176 22800 22206
rect 0 21858 480 21888
rect 3693 21858 3759 21861
rect 0 21856 3759 21858
rect 0 21800 3698 21856
rect 3754 21800 3759 21856
rect 0 21798 3759 21800
rect 0 21768 480 21798
rect 3693 21795 3759 21798
rect 19885 21858 19951 21861
rect 22320 21858 22800 21888
rect 19885 21856 22800 21858
rect 19885 21800 19890 21856
rect 19946 21800 22800 21856
rect 19885 21798 22800 21800
rect 19885 21795 19951 21798
rect 22320 21768 22800 21798
rect 0 21450 480 21480
rect 4061 21450 4127 21453
rect 0 21448 4127 21450
rect 0 21392 4066 21448
rect 4122 21392 4127 21448
rect 0 21390 4127 21392
rect 0 21360 480 21390
rect 4061 21387 4127 21390
rect 18137 21450 18203 21453
rect 22320 21450 22800 21480
rect 18137 21448 22800 21450
rect 18137 21392 18142 21448
rect 18198 21392 22800 21448
rect 18137 21390 22800 21392
rect 18137 21387 18203 21390
rect 22320 21360 22800 21390
rect 0 21042 480 21072
rect 2865 21042 2931 21045
rect 0 21040 2931 21042
rect 0 20984 2870 21040
rect 2926 20984 2931 21040
rect 0 20982 2931 20984
rect 0 20952 480 20982
rect 2865 20979 2931 20982
rect 17953 21042 18019 21045
rect 22320 21042 22800 21072
rect 17953 21040 22800 21042
rect 17953 20984 17958 21040
rect 18014 20984 22800 21040
rect 17953 20982 22800 20984
rect 17953 20979 18019 20982
rect 22320 20952 22800 20982
rect 0 20634 480 20664
rect 1945 20634 2011 20637
rect 0 20632 2011 20634
rect 0 20576 1950 20632
rect 2006 20576 2011 20632
rect 0 20574 2011 20576
rect 0 20544 480 20574
rect 1945 20571 2011 20574
rect 18781 20634 18847 20637
rect 22320 20634 22800 20664
rect 18781 20632 22800 20634
rect 18781 20576 18786 20632
rect 18842 20576 22800 20632
rect 18781 20574 22800 20576
rect 18781 20571 18847 20574
rect 22320 20544 22800 20574
rect 0 20226 480 20256
rect 4061 20226 4127 20229
rect 0 20224 4127 20226
rect 0 20168 4066 20224
rect 4122 20168 4127 20224
rect 0 20166 4127 20168
rect 0 20136 480 20166
rect 4061 20163 4127 20166
rect 20345 20226 20411 20229
rect 22320 20226 22800 20256
rect 20345 20224 22800 20226
rect 20345 20168 20350 20224
rect 20406 20168 22800 20224
rect 20345 20166 22800 20168
rect 20345 20163 20411 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22320 20136 22800 20166
rect 14672 20095 14992 20096
rect 8293 19954 8359 19957
rect 12249 19954 12315 19957
rect 8293 19952 12315 19954
rect 8293 19896 8298 19952
rect 8354 19896 12254 19952
rect 12310 19896 12315 19952
rect 8293 19894 12315 19896
rect 8293 19891 8359 19894
rect 12249 19891 12315 19894
rect 0 19818 480 19848
rect 2773 19818 2839 19821
rect 0 19816 2839 19818
rect 0 19760 2778 19816
rect 2834 19760 2839 19816
rect 0 19758 2839 19760
rect 0 19728 480 19758
rect 2773 19755 2839 19758
rect 11053 19818 11119 19821
rect 17493 19818 17559 19821
rect 11053 19816 17559 19818
rect 11053 19760 11058 19816
rect 11114 19760 17498 19816
rect 17554 19760 17559 19816
rect 11053 19758 17559 19760
rect 11053 19755 11119 19758
rect 17493 19755 17559 19758
rect 18873 19818 18939 19821
rect 22320 19818 22800 19848
rect 18873 19816 22800 19818
rect 18873 19760 18878 19816
rect 18934 19760 22800 19816
rect 18873 19758 22800 19760
rect 18873 19755 18939 19758
rect 22320 19728 22800 19758
rect 16757 19682 16823 19685
rect 17585 19682 17651 19685
rect 11654 19680 17651 19682
rect 11654 19624 16762 19680
rect 16818 19624 17590 19680
rect 17646 19624 17651 19680
rect 11654 19622 17651 19624
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 8661 19546 8727 19549
rect 10777 19546 10843 19549
rect 8661 19544 10843 19546
rect 8661 19488 8666 19544
rect 8722 19488 10782 19544
rect 10838 19488 10843 19544
rect 8661 19486 10843 19488
rect 8661 19483 8727 19486
rect 10777 19483 10843 19486
rect 0 19410 480 19440
rect 1853 19410 1919 19413
rect 0 19408 1919 19410
rect 0 19352 1858 19408
rect 1914 19352 1919 19408
rect 0 19350 1919 19352
rect 0 19320 480 19350
rect 1853 19347 1919 19350
rect 5073 19410 5139 19413
rect 9213 19410 9279 19413
rect 5073 19408 9279 19410
rect 5073 19352 5078 19408
rect 5134 19352 9218 19408
rect 9274 19352 9279 19408
rect 5073 19350 9279 19352
rect 5073 19347 5139 19350
rect 9213 19347 9279 19350
rect 10869 19410 10935 19413
rect 11654 19410 11714 19622
rect 16757 19619 16823 19622
rect 17585 19619 17651 19622
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 12433 19546 12499 19549
rect 16297 19546 16363 19549
rect 12433 19544 16363 19546
rect 12433 19488 12438 19544
rect 12494 19488 16302 19544
rect 16358 19488 16363 19544
rect 12433 19486 16363 19488
rect 12433 19483 12499 19486
rect 16297 19483 16363 19486
rect 10869 19408 11714 19410
rect 10869 19352 10874 19408
rect 10930 19352 11714 19408
rect 10869 19350 11714 19352
rect 14181 19412 14247 19413
rect 14181 19408 14228 19412
rect 14292 19410 14298 19412
rect 15469 19410 15535 19413
rect 22320 19410 22800 19440
rect 14181 19352 14186 19408
rect 10869 19347 10935 19350
rect 14181 19348 14228 19352
rect 14292 19350 14338 19410
rect 15469 19408 22800 19410
rect 15469 19352 15474 19408
rect 15530 19352 22800 19408
rect 15469 19350 22800 19352
rect 14292 19348 14298 19350
rect 14181 19347 14247 19348
rect 15469 19347 15535 19350
rect 22320 19320 22800 19350
rect 17493 19274 17559 19277
rect 2868 19272 17559 19274
rect 2868 19216 17498 19272
rect 17554 19216 17559 19272
rect 2868 19214 17559 19216
rect 0 19138 480 19168
rect 2868 19138 2928 19214
rect 17493 19211 17559 19214
rect 0 19078 2928 19138
rect 3049 19138 3115 19141
rect 5625 19138 5691 19141
rect 3049 19136 5691 19138
rect 3049 19080 3054 19136
rect 3110 19080 5630 19136
rect 5686 19080 5691 19136
rect 3049 19078 5691 19080
rect 0 19048 480 19078
rect 3049 19075 3115 19078
rect 5625 19075 5691 19078
rect 8845 19138 8911 19141
rect 12198 19138 12204 19140
rect 8845 19136 12204 19138
rect 8845 19080 8850 19136
rect 8906 19080 12204 19136
rect 8845 19078 12204 19080
rect 8845 19075 8911 19078
rect 12198 19076 12204 19078
rect 12268 19138 12274 19140
rect 14365 19138 14431 19141
rect 12268 19136 14431 19138
rect 12268 19080 14370 19136
rect 14426 19080 14431 19136
rect 12268 19078 14431 19080
rect 12268 19076 12274 19078
rect 14365 19075 14431 19078
rect 17585 19138 17651 19141
rect 22320 19138 22800 19168
rect 17585 19136 22800 19138
rect 17585 19080 17590 19136
rect 17646 19080 22800 19136
rect 17585 19078 22800 19080
rect 17585 19075 17651 19078
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 22320 19048 22800 19078
rect 14672 19007 14992 19008
rect 1577 19002 1643 19005
rect 6361 19002 6427 19005
rect 1577 19000 6427 19002
rect 1577 18944 1582 19000
rect 1638 18944 6366 19000
rect 6422 18944 6427 19000
rect 1577 18942 6427 18944
rect 1577 18939 1643 18942
rect 6361 18939 6427 18942
rect 8201 19002 8267 19005
rect 11053 19002 11119 19005
rect 11830 19002 11836 19004
rect 8201 19000 11836 19002
rect 8201 18944 8206 19000
rect 8262 18944 11058 19000
rect 11114 18944 11836 19000
rect 8201 18942 11836 18944
rect 8201 18939 8267 18942
rect 11053 18939 11119 18942
rect 11830 18940 11836 18942
rect 11900 18940 11906 19004
rect 16430 18940 16436 19004
rect 16500 19002 16506 19004
rect 19149 19002 19215 19005
rect 16500 19000 19215 19002
rect 16500 18944 19154 19000
rect 19210 18944 19215 19000
rect 16500 18942 19215 18944
rect 16500 18940 16506 18942
rect 19149 18939 19215 18942
rect 4429 18866 4495 18869
rect 9673 18868 9739 18869
rect 4429 18864 8402 18866
rect 4429 18808 4434 18864
rect 4490 18808 8402 18864
rect 4429 18806 8402 18808
rect 4429 18803 4495 18806
rect 0 18730 480 18760
rect 1945 18730 2011 18733
rect 0 18728 2011 18730
rect 0 18672 1950 18728
rect 2006 18672 2011 18728
rect 0 18670 2011 18672
rect 0 18640 480 18670
rect 1945 18667 2011 18670
rect 2497 18730 2563 18733
rect 2497 18728 8218 18730
rect 2497 18672 2502 18728
rect 2558 18672 8218 18728
rect 2497 18670 8218 18672
rect 2497 18667 2563 18670
rect 4797 18594 4863 18597
rect 7741 18594 7807 18597
rect 4797 18592 7807 18594
rect 4797 18536 4802 18592
rect 4858 18536 7746 18592
rect 7802 18536 7807 18592
rect 4797 18534 7807 18536
rect 4797 18531 4863 18534
rect 7741 18531 7807 18534
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 2313 18458 2379 18461
rect 8017 18458 8083 18461
rect 2313 18456 4308 18458
rect 2313 18400 2318 18456
rect 2374 18400 4308 18456
rect 2313 18398 4308 18400
rect 2313 18395 2379 18398
rect 0 18322 480 18352
rect 3601 18322 3667 18325
rect 0 18320 3667 18322
rect 0 18264 3606 18320
rect 3662 18264 3667 18320
rect 0 18262 3667 18264
rect 4248 18322 4308 18398
rect 6686 18456 8083 18458
rect 6686 18400 8022 18456
rect 8078 18400 8083 18456
rect 6686 18398 8083 18400
rect 8158 18458 8218 18670
rect 8342 18594 8402 18806
rect 9622 18804 9628 18868
rect 9692 18866 9739 18868
rect 9692 18864 9784 18866
rect 9734 18808 9784 18864
rect 9692 18806 9784 18808
rect 9692 18804 9739 18806
rect 10542 18804 10548 18868
rect 10612 18866 10618 18868
rect 15377 18866 15443 18869
rect 10612 18864 15443 18866
rect 10612 18808 15382 18864
rect 15438 18808 15443 18864
rect 10612 18806 15443 18808
rect 10612 18804 10618 18806
rect 9673 18803 9739 18804
rect 15377 18803 15443 18806
rect 17217 18866 17283 18869
rect 17677 18866 17743 18869
rect 17953 18866 18019 18869
rect 17217 18864 18019 18866
rect 17217 18808 17222 18864
rect 17278 18808 17682 18864
rect 17738 18808 17958 18864
rect 18014 18808 18019 18864
rect 17217 18806 18019 18808
rect 17217 18803 17283 18806
rect 17677 18803 17743 18806
rect 17953 18803 18019 18806
rect 8477 18730 8543 18733
rect 8886 18730 8892 18732
rect 8477 18728 8892 18730
rect 8477 18672 8482 18728
rect 8538 18672 8892 18728
rect 8477 18670 8892 18672
rect 8477 18667 8543 18670
rect 8886 18668 8892 18670
rect 8956 18730 8962 18732
rect 8956 18670 11714 18730
rect 8956 18668 8962 18670
rect 10685 18594 10751 18597
rect 8342 18592 10751 18594
rect 8342 18536 10690 18592
rect 10746 18536 10751 18592
rect 8342 18534 10751 18536
rect 11654 18594 11714 18670
rect 12750 18668 12756 18732
rect 12820 18730 12826 18732
rect 18137 18730 18203 18733
rect 12820 18728 18203 18730
rect 12820 18672 18142 18728
rect 18198 18672 18203 18728
rect 12820 18670 18203 18672
rect 12820 18668 12826 18670
rect 18137 18667 18203 18670
rect 18597 18730 18663 18733
rect 22320 18730 22800 18760
rect 18597 18728 22800 18730
rect 18597 18672 18602 18728
rect 18658 18672 22800 18728
rect 18597 18670 22800 18672
rect 18597 18667 18663 18670
rect 22320 18640 22800 18670
rect 16389 18594 16455 18597
rect 11654 18592 16455 18594
rect 11654 18536 16394 18592
rect 16450 18536 16455 18592
rect 11654 18534 16455 18536
rect 10685 18531 10751 18534
rect 16389 18531 16455 18534
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 8845 18458 8911 18461
rect 8158 18456 8911 18458
rect 8158 18400 8850 18456
rect 8906 18400 8911 18456
rect 8158 18398 8911 18400
rect 6686 18322 6746 18398
rect 8017 18395 8083 18398
rect 8845 18395 8911 18398
rect 9397 18458 9463 18461
rect 9622 18458 9628 18460
rect 9397 18456 9628 18458
rect 9397 18400 9402 18456
rect 9458 18400 9628 18456
rect 9397 18398 9628 18400
rect 9397 18395 9463 18398
rect 9622 18396 9628 18398
rect 9692 18396 9698 18460
rect 9765 18458 9831 18461
rect 10777 18458 10843 18461
rect 9765 18456 10843 18458
rect 9765 18400 9770 18456
rect 9826 18400 10782 18456
rect 10838 18400 10843 18456
rect 9765 18398 10843 18400
rect 9765 18395 9831 18398
rect 10777 18395 10843 18398
rect 13854 18396 13860 18460
rect 13924 18458 13930 18460
rect 14549 18458 14615 18461
rect 13924 18456 14615 18458
rect 13924 18400 14554 18456
rect 14610 18400 14615 18456
rect 13924 18398 14615 18400
rect 13924 18396 13930 18398
rect 14549 18395 14615 18398
rect 15285 18458 15351 18461
rect 16113 18458 16179 18461
rect 15285 18456 16179 18458
rect 15285 18400 15290 18456
rect 15346 18400 16118 18456
rect 16174 18400 16179 18456
rect 15285 18398 16179 18400
rect 15285 18395 15351 18398
rect 16113 18395 16179 18398
rect 4248 18262 6746 18322
rect 6821 18322 6887 18325
rect 10133 18322 10199 18325
rect 6821 18320 10199 18322
rect 6821 18264 6826 18320
rect 6882 18264 10138 18320
rect 10194 18264 10199 18320
rect 6821 18262 10199 18264
rect 0 18232 480 18262
rect 3601 18259 3667 18262
rect 6821 18259 6887 18262
rect 10133 18259 10199 18262
rect 10777 18322 10843 18325
rect 17033 18322 17099 18325
rect 10777 18320 17099 18322
rect 10777 18264 10782 18320
rect 10838 18264 17038 18320
rect 17094 18264 17099 18320
rect 10777 18262 17099 18264
rect 10777 18259 10843 18262
rect 17033 18259 17099 18262
rect 17953 18322 18019 18325
rect 22320 18322 22800 18352
rect 17953 18320 22800 18322
rect 17953 18264 17958 18320
rect 18014 18264 22800 18320
rect 17953 18262 22800 18264
rect 17953 18259 18019 18262
rect 22320 18232 22800 18262
rect 4981 18186 5047 18189
rect 11973 18186 12039 18189
rect 4981 18184 12039 18186
rect 4981 18128 4986 18184
rect 5042 18128 11978 18184
rect 12034 18128 12039 18184
rect 4981 18126 12039 18128
rect 4981 18123 5047 18126
rect 11973 18123 12039 18126
rect 12157 18186 12223 18189
rect 13997 18186 14063 18189
rect 16481 18186 16547 18189
rect 12157 18184 14063 18186
rect 12157 18128 12162 18184
rect 12218 18128 14002 18184
rect 14058 18128 14063 18184
rect 12157 18126 14063 18128
rect 12157 18123 12223 18126
rect 13997 18123 14063 18126
rect 14414 18184 16547 18186
rect 14414 18128 16486 18184
rect 16542 18128 16547 18184
rect 14414 18126 16547 18128
rect 3693 18050 3759 18053
rect 6361 18050 6427 18053
rect 3693 18048 6427 18050
rect 3693 17992 3698 18048
rect 3754 17992 6366 18048
rect 6422 17992 6427 18048
rect 3693 17990 6427 17992
rect 3693 17987 3759 17990
rect 6361 17987 6427 17990
rect 7046 17988 7052 18052
rect 7116 18050 7122 18052
rect 7189 18050 7255 18053
rect 7116 18048 7255 18050
rect 7116 17992 7194 18048
rect 7250 17992 7255 18048
rect 7116 17990 7255 17992
rect 7116 17988 7122 17990
rect 7189 17987 7255 17990
rect 8518 17988 8524 18052
rect 8588 18050 8594 18052
rect 8661 18050 8727 18053
rect 8588 18048 8727 18050
rect 8588 17992 8666 18048
rect 8722 17992 8727 18048
rect 8588 17990 8727 17992
rect 8588 17988 8594 17990
rect 8661 17987 8727 17990
rect 10358 17988 10364 18052
rect 10428 18050 10434 18052
rect 14414 18050 14474 18126
rect 16481 18123 16547 18126
rect 17677 18186 17743 18189
rect 19149 18186 19215 18189
rect 17677 18184 19215 18186
rect 17677 18128 17682 18184
rect 17738 18128 19154 18184
rect 19210 18128 19215 18184
rect 17677 18126 19215 18128
rect 17677 18123 17743 18126
rect 19149 18123 19215 18126
rect 10428 17990 14474 18050
rect 10428 17988 10434 17990
rect 15142 17988 15148 18052
rect 15212 18050 15218 18052
rect 16021 18050 16087 18053
rect 15212 18048 16087 18050
rect 15212 17992 16026 18048
rect 16082 17992 16087 18048
rect 15212 17990 16087 17992
rect 15212 17988 15218 17990
rect 16021 17987 16087 17990
rect 17217 18050 17283 18053
rect 17350 18050 17356 18052
rect 17217 18048 17356 18050
rect 17217 17992 17222 18048
rect 17278 17992 17356 18048
rect 17217 17990 17356 17992
rect 17217 17987 17283 17990
rect 17350 17988 17356 17990
rect 17420 17988 17426 18052
rect 17902 17988 17908 18052
rect 17972 18050 17978 18052
rect 18413 18050 18479 18053
rect 17972 18048 18479 18050
rect 17972 17992 18418 18048
rect 18474 17992 18479 18048
rect 17972 17990 18479 17992
rect 17972 17988 17978 17990
rect 18413 17987 18479 17990
rect 18638 17988 18644 18052
rect 18708 18050 18714 18052
rect 19149 18050 19215 18053
rect 18708 18048 19215 18050
rect 18708 17992 19154 18048
rect 19210 17992 19215 18048
rect 18708 17990 19215 17992
rect 18708 17988 18714 17990
rect 19149 17987 19215 17990
rect 7808 17984 8128 17985
rect 0 17914 480 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 1485 17914 1551 17917
rect 0 17912 1551 17914
rect 0 17856 1490 17912
rect 1546 17856 1551 17912
rect 0 17854 1551 17856
rect 0 17824 480 17854
rect 1485 17851 1551 17854
rect 1853 17914 1919 17917
rect 5257 17914 5323 17917
rect 6729 17914 6795 17917
rect 1853 17912 6795 17914
rect 1853 17856 1858 17912
rect 1914 17856 5262 17912
rect 5318 17856 6734 17912
rect 6790 17856 6795 17912
rect 1853 17854 6795 17856
rect 1853 17851 1919 17854
rect 5257 17851 5323 17854
rect 6729 17851 6795 17854
rect 8293 17914 8359 17917
rect 9029 17914 9095 17917
rect 8293 17912 9095 17914
rect 8293 17856 8298 17912
rect 8354 17856 9034 17912
rect 9090 17856 9095 17912
rect 8293 17854 9095 17856
rect 8293 17851 8359 17854
rect 9029 17851 9095 17854
rect 9857 17914 9923 17917
rect 11789 17914 11855 17917
rect 9857 17912 11855 17914
rect 9857 17856 9862 17912
rect 9918 17856 11794 17912
rect 11850 17856 11855 17912
rect 9857 17854 11855 17856
rect 9857 17851 9923 17854
rect 11789 17851 11855 17854
rect 15193 17914 15259 17917
rect 18045 17914 18111 17917
rect 15193 17912 18111 17914
rect 15193 17856 15198 17912
rect 15254 17856 18050 17912
rect 18106 17856 18111 17912
rect 15193 17854 18111 17856
rect 15193 17851 15259 17854
rect 18045 17851 18111 17854
rect 18229 17914 18295 17917
rect 22320 17914 22800 17944
rect 18229 17912 22800 17914
rect 18229 17856 18234 17912
rect 18290 17856 22800 17912
rect 18229 17854 22800 17856
rect 18229 17851 18295 17854
rect 22320 17824 22800 17854
rect 2405 17778 2471 17781
rect 5758 17778 5764 17780
rect 2405 17776 5764 17778
rect 2405 17720 2410 17776
rect 2466 17720 5764 17776
rect 2405 17718 5764 17720
rect 2405 17715 2471 17718
rect 5758 17716 5764 17718
rect 5828 17778 5834 17780
rect 12157 17778 12223 17781
rect 5828 17776 12223 17778
rect 5828 17720 12162 17776
rect 12218 17720 12223 17776
rect 5828 17718 12223 17720
rect 5828 17716 5834 17718
rect 12157 17715 12223 17718
rect 15101 17778 15167 17781
rect 17585 17778 17651 17781
rect 15101 17776 17651 17778
rect 15101 17720 15106 17776
rect 15162 17720 17590 17776
rect 17646 17720 17651 17776
rect 15101 17718 17651 17720
rect 15101 17715 15167 17718
rect 17585 17715 17651 17718
rect 3785 17642 3851 17645
rect 5533 17642 5599 17645
rect 3785 17640 5599 17642
rect 3785 17584 3790 17640
rect 3846 17584 5538 17640
rect 5594 17584 5599 17640
rect 3785 17582 5599 17584
rect 3785 17579 3851 17582
rect 5533 17579 5599 17582
rect 6361 17642 6427 17645
rect 12065 17642 12131 17645
rect 16021 17642 16087 17645
rect 6361 17640 11944 17642
rect 6361 17584 6366 17640
rect 6422 17584 11944 17640
rect 6361 17582 11944 17584
rect 6361 17579 6427 17582
rect 0 17506 480 17536
rect 1577 17506 1643 17509
rect 0 17504 1643 17506
rect 0 17448 1582 17504
rect 1638 17448 1643 17504
rect 0 17446 1643 17448
rect 0 17416 480 17446
rect 1577 17443 1643 17446
rect 7281 17506 7347 17509
rect 9489 17506 9555 17509
rect 7281 17504 9555 17506
rect 7281 17448 7286 17504
rect 7342 17448 9494 17504
rect 9550 17448 9555 17504
rect 7281 17446 9555 17448
rect 7281 17443 7347 17446
rect 9489 17443 9555 17446
rect 4376 17440 4696 17441
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 11884 17370 11944 17582
rect 12065 17640 16087 17642
rect 12065 17584 12070 17640
rect 12126 17584 16026 17640
rect 16082 17584 16087 17640
rect 12065 17582 16087 17584
rect 12065 17579 12131 17582
rect 16021 17579 16087 17582
rect 16246 17580 16252 17644
rect 16316 17642 16322 17644
rect 19517 17642 19583 17645
rect 16316 17640 19583 17642
rect 16316 17584 19522 17640
rect 19578 17584 19583 17640
rect 16316 17582 19583 17584
rect 16316 17580 16322 17582
rect 19517 17579 19583 17582
rect 12382 17444 12388 17508
rect 12452 17506 12458 17508
rect 15009 17506 15075 17509
rect 12452 17504 15075 17506
rect 12452 17448 15014 17504
rect 15070 17448 15075 17504
rect 12452 17446 15075 17448
rect 12452 17444 12458 17446
rect 15009 17443 15075 17446
rect 15694 17444 15700 17508
rect 15764 17506 15770 17508
rect 15837 17506 15903 17509
rect 15764 17504 15903 17506
rect 15764 17448 15842 17504
rect 15898 17448 15903 17504
rect 15764 17446 15903 17448
rect 15764 17444 15770 17446
rect 15837 17443 15903 17446
rect 18873 17506 18939 17509
rect 22320 17506 22800 17536
rect 18873 17504 22800 17506
rect 18873 17448 18878 17504
rect 18934 17448 22800 17504
rect 18873 17446 22800 17448
rect 18873 17443 18939 17446
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 22320 17416 22800 17446
rect 18104 17375 18424 17376
rect 17861 17370 17927 17373
rect 11884 17368 17927 17370
rect 11884 17312 17866 17368
rect 17922 17312 17927 17368
rect 11884 17310 17927 17312
rect 17861 17307 17927 17310
rect 2313 17234 2379 17237
rect 5206 17234 5212 17236
rect 2313 17232 5212 17234
rect 2313 17176 2318 17232
rect 2374 17176 5212 17232
rect 2313 17174 5212 17176
rect 2313 17171 2379 17174
rect 5206 17172 5212 17174
rect 5276 17234 5282 17236
rect 17953 17234 18019 17237
rect 5276 17232 18019 17234
rect 5276 17176 17958 17232
rect 18014 17176 18019 17232
rect 5276 17174 18019 17176
rect 5276 17172 5282 17174
rect 17953 17171 18019 17174
rect 0 17098 480 17128
rect 3049 17098 3115 17101
rect 0 17096 3115 17098
rect 0 17040 3054 17096
rect 3110 17040 3115 17096
rect 0 17038 3115 17040
rect 0 17008 480 17038
rect 3049 17035 3115 17038
rect 3601 17098 3667 17101
rect 4705 17098 4771 17101
rect 3601 17096 4771 17098
rect 3601 17040 3606 17096
rect 3662 17040 4710 17096
rect 4766 17040 4771 17096
rect 3601 17038 4771 17040
rect 3601 17035 3667 17038
rect 4705 17035 4771 17038
rect 8017 17098 8083 17101
rect 11973 17100 12039 17101
rect 11646 17098 11652 17100
rect 8017 17096 11652 17098
rect 8017 17040 8022 17096
rect 8078 17040 11652 17096
rect 8017 17038 11652 17040
rect 8017 17035 8083 17038
rect 11646 17036 11652 17038
rect 11716 17036 11722 17100
rect 11973 17096 12020 17100
rect 12084 17098 12090 17100
rect 12617 17098 12683 17101
rect 12084 17096 12683 17098
rect 11973 17040 11978 17096
rect 12084 17040 12622 17096
rect 12678 17040 12683 17096
rect 11973 17036 12020 17040
rect 12084 17038 12683 17040
rect 12084 17036 12090 17038
rect 11973 17035 12039 17036
rect 12617 17035 12683 17038
rect 13169 17098 13235 17101
rect 18597 17098 18663 17101
rect 13169 17096 18663 17098
rect 13169 17040 13174 17096
rect 13230 17040 18602 17096
rect 18658 17040 18663 17096
rect 13169 17038 18663 17040
rect 13169 17035 13235 17038
rect 18597 17035 18663 17038
rect 18873 17096 18939 17101
rect 18873 17040 18878 17096
rect 18934 17040 18939 17096
rect 18873 17035 18939 17040
rect 20897 17098 20963 17101
rect 22320 17098 22800 17128
rect 20897 17096 22800 17098
rect 20897 17040 20902 17096
rect 20958 17040 22800 17096
rect 20897 17038 22800 17040
rect 20897 17035 20963 17038
rect 9070 16900 9076 16964
rect 9140 16962 9146 16964
rect 9673 16962 9739 16965
rect 9140 16960 9739 16962
rect 9140 16904 9678 16960
rect 9734 16904 9739 16960
rect 9140 16902 9739 16904
rect 9140 16900 9146 16902
rect 9673 16899 9739 16902
rect 10685 16962 10751 16965
rect 14089 16962 14155 16965
rect 10685 16960 14155 16962
rect 10685 16904 10690 16960
rect 10746 16904 14094 16960
rect 14150 16904 14155 16960
rect 10685 16902 14155 16904
rect 10685 16899 10751 16902
rect 14089 16899 14155 16902
rect 17217 16962 17283 16965
rect 18876 16962 18936 17035
rect 22320 17008 22800 17038
rect 17217 16960 18936 16962
rect 17217 16904 17222 16960
rect 17278 16904 18936 16960
rect 17217 16902 18936 16904
rect 17217 16899 17283 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 3693 16826 3759 16829
rect 1350 16824 3759 16826
rect 1350 16768 3698 16824
rect 3754 16768 3759 16824
rect 1350 16766 3759 16768
rect 0 16690 480 16720
rect 1350 16690 1410 16766
rect 3693 16763 3759 16766
rect 10041 16826 10107 16829
rect 16021 16826 16087 16829
rect 10041 16824 12772 16826
rect 10041 16768 10046 16824
rect 10102 16768 12772 16824
rect 10041 16766 12772 16768
rect 10041 16763 10107 16766
rect 0 16630 1410 16690
rect 3417 16690 3483 16693
rect 3550 16690 3556 16692
rect 3417 16688 3556 16690
rect 3417 16632 3422 16688
rect 3478 16632 3556 16688
rect 3417 16630 3556 16632
rect 0 16600 480 16630
rect 3417 16627 3483 16630
rect 3550 16628 3556 16630
rect 3620 16628 3626 16692
rect 10317 16690 10383 16693
rect 12065 16690 12131 16693
rect 10317 16688 12131 16690
rect 10317 16632 10322 16688
rect 10378 16632 12070 16688
rect 12126 16632 12131 16688
rect 10317 16630 12131 16632
rect 10317 16627 10383 16630
rect 12065 16627 12131 16630
rect 3325 16554 3391 16557
rect 4838 16554 4844 16556
rect 3325 16552 4844 16554
rect 3325 16496 3330 16552
rect 3386 16496 4844 16552
rect 3325 16494 4844 16496
rect 3325 16491 3391 16494
rect 4838 16492 4844 16494
rect 4908 16554 4914 16556
rect 12712 16554 12772 16766
rect 16021 16824 20362 16826
rect 16021 16768 16026 16824
rect 16082 16768 20362 16824
rect 16021 16766 20362 16768
rect 16021 16763 16087 16766
rect 14549 16690 14615 16693
rect 17033 16690 17099 16693
rect 17309 16690 17375 16693
rect 14549 16688 17099 16690
rect 14549 16632 14554 16688
rect 14610 16632 17038 16688
rect 17094 16632 17099 16688
rect 14549 16630 17099 16632
rect 14549 16627 14615 16630
rect 17033 16627 17099 16630
rect 17174 16688 17375 16690
rect 17174 16632 17314 16688
rect 17370 16632 17375 16688
rect 17174 16630 17375 16632
rect 17174 16554 17234 16630
rect 17309 16627 17375 16630
rect 17585 16690 17651 16693
rect 19241 16692 19307 16693
rect 17718 16690 17724 16692
rect 17585 16688 17724 16690
rect 17585 16632 17590 16688
rect 17646 16632 17724 16688
rect 17585 16630 17724 16632
rect 17585 16627 17651 16630
rect 17718 16628 17724 16630
rect 17788 16628 17794 16692
rect 19190 16690 19196 16692
rect 19150 16630 19196 16690
rect 19260 16688 19307 16692
rect 19302 16632 19307 16688
rect 19190 16628 19196 16630
rect 19260 16628 19307 16632
rect 19241 16627 19307 16628
rect 19517 16692 19583 16693
rect 20069 16692 20135 16693
rect 19517 16688 19564 16692
rect 19628 16690 19634 16692
rect 19517 16632 19522 16688
rect 19517 16628 19564 16632
rect 19628 16630 19674 16690
rect 20069 16688 20116 16692
rect 20180 16690 20186 16692
rect 20302 16690 20362 16766
rect 22320 16690 22800 16720
rect 20069 16632 20074 16688
rect 19628 16628 19634 16630
rect 20069 16628 20116 16632
rect 20180 16630 20226 16690
rect 20302 16630 22800 16690
rect 20180 16628 20186 16630
rect 19517 16627 19583 16628
rect 20069 16627 20135 16628
rect 22320 16600 22800 16630
rect 4908 16494 12496 16554
rect 12712 16494 17234 16554
rect 4908 16492 4914 16494
rect 10685 16418 10751 16421
rect 10910 16418 10916 16420
rect 10685 16416 10916 16418
rect 10685 16360 10690 16416
rect 10746 16360 10916 16416
rect 10685 16358 10916 16360
rect 10685 16355 10751 16358
rect 10910 16356 10916 16358
rect 10980 16356 10986 16420
rect 4376 16352 4696 16353
rect 0 16282 480 16312
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 1117 16282 1183 16285
rect 0 16280 1183 16282
rect 0 16224 1122 16280
rect 1178 16224 1183 16280
rect 0 16222 1183 16224
rect 12436 16282 12496 16494
rect 15193 16418 15259 16421
rect 16205 16418 16271 16421
rect 15193 16416 16271 16418
rect 15193 16360 15198 16416
rect 15254 16360 16210 16416
rect 16266 16360 16271 16416
rect 15193 16358 16271 16360
rect 15193 16355 15259 16358
rect 16205 16355 16271 16358
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 19701 16284 19767 16285
rect 12436 16222 17970 16282
rect 0 16192 480 16222
rect 1117 16219 1183 16222
rect 8477 16146 8543 16149
rect 12433 16146 12499 16149
rect 8477 16144 12499 16146
rect 8477 16088 8482 16144
rect 8538 16088 12438 16144
rect 12494 16088 12499 16144
rect 8477 16086 12499 16088
rect 8477 16083 8586 16086
rect 12433 16083 12499 16086
rect 12709 16146 12775 16149
rect 12934 16146 12940 16148
rect 12709 16144 12940 16146
rect 12709 16088 12714 16144
rect 12770 16088 12940 16144
rect 12709 16086 12940 16088
rect 12709 16083 12775 16086
rect 12934 16084 12940 16086
rect 13004 16084 13010 16148
rect 16113 16146 16179 16149
rect 17769 16146 17835 16149
rect 16113 16144 17835 16146
rect 16113 16088 16118 16144
rect 16174 16088 17774 16144
rect 17830 16088 17835 16144
rect 16113 16086 17835 16088
rect 17910 16146 17970 16222
rect 19701 16280 19748 16284
rect 19812 16282 19818 16284
rect 21173 16282 21239 16285
rect 22320 16282 22800 16312
rect 19701 16224 19706 16280
rect 19701 16220 19748 16224
rect 19812 16222 19858 16282
rect 21173 16280 22800 16282
rect 21173 16224 21178 16280
rect 21234 16224 22800 16280
rect 21173 16222 22800 16224
rect 19812 16220 19818 16222
rect 19701 16219 19767 16220
rect 21173 16219 21239 16222
rect 22320 16192 22800 16222
rect 20529 16146 20595 16149
rect 17910 16144 20595 16146
rect 17910 16088 20534 16144
rect 20590 16088 20595 16144
rect 17910 16086 20595 16088
rect 16113 16083 16179 16086
rect 17769 16083 17835 16086
rect 20529 16083 20595 16086
rect 2313 16010 2379 16013
rect 8334 16010 8340 16012
rect 2313 16008 8340 16010
rect 2313 15952 2318 16008
rect 2374 15952 8340 16008
rect 2313 15950 8340 15952
rect 2313 15947 2379 15950
rect 8334 15948 8340 15950
rect 8404 15948 8410 16012
rect 0 15874 480 15904
rect 4061 15874 4127 15877
rect 0 15872 4127 15874
rect 0 15816 4066 15872
rect 4122 15816 4127 15872
rect 0 15814 4127 15816
rect 8526 15874 8586 16083
rect 8845 16010 8911 16013
rect 16430 16010 16436 16012
rect 8845 16008 16436 16010
rect 8845 15952 8850 16008
rect 8906 15952 16436 16008
rect 8845 15950 16436 15952
rect 8845 15947 8911 15950
rect 16430 15948 16436 15950
rect 16500 15948 16506 16012
rect 18597 16010 18663 16013
rect 19006 16010 19012 16012
rect 18597 16008 19012 16010
rect 18597 15952 18602 16008
rect 18658 15952 19012 16008
rect 18597 15950 19012 15952
rect 18597 15947 18663 15950
rect 19006 15948 19012 15950
rect 19076 15948 19082 16012
rect 8753 15874 8819 15877
rect 8526 15872 8819 15874
rect 8526 15816 8758 15872
rect 8814 15816 8819 15872
rect 8526 15814 8819 15816
rect 0 15784 480 15814
rect 4061 15811 4127 15814
rect 8753 15811 8819 15814
rect 15101 15874 15167 15877
rect 15326 15874 15332 15876
rect 15101 15872 15332 15874
rect 15101 15816 15106 15872
rect 15162 15816 15332 15872
rect 15101 15814 15332 15816
rect 15101 15811 15167 15814
rect 15326 15812 15332 15814
rect 15396 15812 15402 15876
rect 19241 15874 19307 15877
rect 22320 15874 22800 15904
rect 19241 15872 22800 15874
rect 19241 15816 19246 15872
rect 19302 15816 22800 15872
rect 19241 15814 22800 15816
rect 19241 15811 19307 15814
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 22320 15784 22800 15814
rect 14672 15743 14992 15744
rect 2589 15738 2655 15741
rect 5901 15738 5967 15741
rect 2589 15736 5967 15738
rect 2589 15680 2594 15736
rect 2650 15680 5906 15736
rect 5962 15680 5967 15736
rect 2589 15678 5967 15680
rect 2589 15675 2655 15678
rect 5901 15675 5967 15678
rect 6453 15738 6519 15741
rect 7465 15738 7531 15741
rect 6453 15736 7531 15738
rect 6453 15680 6458 15736
rect 6514 15680 7470 15736
rect 7526 15680 7531 15736
rect 6453 15678 7531 15680
rect 6453 15675 6519 15678
rect 7465 15675 7531 15678
rect 9673 15738 9739 15741
rect 11145 15738 11211 15741
rect 9673 15736 11211 15738
rect 9673 15680 9678 15736
rect 9734 15680 11150 15736
rect 11206 15680 11211 15736
rect 9673 15678 11211 15680
rect 9673 15675 9739 15678
rect 11145 15675 11211 15678
rect 12433 15738 12499 15741
rect 12566 15738 12572 15740
rect 12433 15736 12572 15738
rect 12433 15680 12438 15736
rect 12494 15680 12572 15736
rect 12433 15678 12572 15680
rect 12433 15675 12499 15678
rect 12566 15676 12572 15678
rect 12636 15738 12642 15740
rect 13537 15738 13603 15741
rect 14089 15738 14155 15741
rect 12636 15736 14155 15738
rect 12636 15680 13542 15736
rect 13598 15680 14094 15736
rect 14150 15680 14155 15736
rect 12636 15678 14155 15680
rect 12636 15676 12642 15678
rect 13537 15675 13603 15678
rect 14089 15675 14155 15678
rect 15101 15738 15167 15741
rect 18597 15738 18663 15741
rect 15101 15736 18663 15738
rect 15101 15680 15106 15736
rect 15162 15680 18602 15736
rect 18658 15680 18663 15736
rect 15101 15678 18663 15680
rect 15101 15675 15167 15678
rect 18597 15675 18663 15678
rect 4889 15602 4955 15605
rect 15009 15602 15075 15605
rect 4889 15600 15075 15602
rect 4889 15544 4894 15600
rect 4950 15544 15014 15600
rect 15070 15544 15075 15600
rect 4889 15542 15075 15544
rect 4889 15539 4955 15542
rect 0 15466 480 15496
rect 3877 15466 3943 15469
rect 0 15464 3943 15466
rect 0 15408 3882 15464
rect 3938 15408 3943 15464
rect 0 15406 3943 15408
rect 0 15376 480 15406
rect 3877 15403 3943 15406
rect 4376 15264 4696 15265
rect 0 15194 480 15224
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 3969 15194 4035 15197
rect 0 15192 4035 15194
rect 0 15136 3974 15192
rect 4030 15136 4035 15192
rect 0 15134 4035 15136
rect 0 15104 480 15134
rect 3969 15131 4035 15134
rect 0 14786 480 14816
rect 5030 14789 5090 15542
rect 15009 15539 15075 15542
rect 15745 15602 15811 15605
rect 16430 15602 16436 15604
rect 15745 15600 16436 15602
rect 15745 15544 15750 15600
rect 15806 15544 16436 15600
rect 15745 15542 16436 15544
rect 15745 15539 15811 15542
rect 16430 15540 16436 15542
rect 16500 15540 16506 15604
rect 16982 15540 16988 15604
rect 17052 15602 17058 15604
rect 17861 15602 17927 15605
rect 17052 15600 17927 15602
rect 17052 15544 17866 15600
rect 17922 15544 17927 15600
rect 17052 15542 17927 15544
rect 17052 15540 17058 15542
rect 17861 15539 17927 15542
rect 18965 15602 19031 15605
rect 20805 15602 20871 15605
rect 18965 15600 20871 15602
rect 18965 15544 18970 15600
rect 19026 15544 20810 15600
rect 20866 15544 20871 15600
rect 18965 15542 20871 15544
rect 18965 15539 19031 15542
rect 20805 15539 20871 15542
rect 6637 15468 6703 15469
rect 6637 15464 6684 15468
rect 6748 15466 6754 15468
rect 6637 15408 6642 15464
rect 6637 15404 6684 15408
rect 6748 15406 6794 15466
rect 6748 15404 6754 15406
rect 13302 15404 13308 15468
rect 13372 15466 13378 15468
rect 15561 15466 15627 15469
rect 13372 15464 15627 15466
rect 13372 15408 15566 15464
rect 15622 15408 15627 15464
rect 13372 15406 15627 15408
rect 13372 15404 13378 15406
rect 6637 15403 6703 15404
rect 15561 15403 15627 15406
rect 15837 15466 15903 15469
rect 22320 15466 22800 15496
rect 15837 15464 22800 15466
rect 15837 15408 15842 15464
rect 15898 15408 22800 15464
rect 15837 15406 22800 15408
rect 15837 15403 15903 15406
rect 22320 15376 22800 15406
rect 5349 15330 5415 15333
rect 7925 15330 7991 15333
rect 5349 15328 7991 15330
rect 5349 15272 5354 15328
rect 5410 15272 7930 15328
rect 7986 15272 7991 15328
rect 5349 15270 7991 15272
rect 5349 15267 5415 15270
rect 7925 15267 7991 15270
rect 12249 15330 12315 15333
rect 19425 15332 19491 15333
rect 19374 15330 19380 15332
rect 12249 15328 16084 15330
rect 12249 15272 12254 15328
rect 12310 15272 16084 15328
rect 12249 15270 16084 15272
rect 19334 15270 19380 15330
rect 19444 15328 19491 15332
rect 19486 15272 19491 15328
rect 12249 15267 12315 15270
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 16024 15197 16084 15270
rect 19374 15268 19380 15270
rect 19444 15268 19491 15272
rect 19425 15267 19491 15268
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 5257 15194 5323 15197
rect 8477 15194 8543 15197
rect 15653 15194 15719 15197
rect 5257 15192 8543 15194
rect 5257 15136 5262 15192
rect 5318 15136 8482 15192
rect 8538 15136 8543 15192
rect 5257 15134 8543 15136
rect 5257 15131 5323 15134
rect 8477 15131 8543 15134
rect 12252 15192 15719 15194
rect 12252 15136 15658 15192
rect 15714 15136 15719 15192
rect 12252 15134 15719 15136
rect 7281 15058 7347 15061
rect 7741 15058 7807 15061
rect 7281 15056 7807 15058
rect 7281 15000 7286 15056
rect 7342 15000 7746 15056
rect 7802 15000 7807 15056
rect 7281 14998 7807 15000
rect 7281 14995 7347 14998
rect 7741 14995 7807 14998
rect 11513 15058 11579 15061
rect 12252 15058 12312 15134
rect 15653 15131 15719 15134
rect 16021 15192 16087 15197
rect 16021 15136 16026 15192
rect 16082 15136 16087 15192
rect 16021 15131 16087 15136
rect 18822 15132 18828 15196
rect 18892 15194 18898 15196
rect 19425 15194 19491 15197
rect 22320 15194 22800 15224
rect 18892 15192 19491 15194
rect 18892 15136 19430 15192
rect 19486 15136 19491 15192
rect 18892 15134 19491 15136
rect 18892 15132 18898 15134
rect 19425 15131 19491 15134
rect 19934 15134 22800 15194
rect 11513 15056 12312 15058
rect 11513 15000 11518 15056
rect 11574 15000 12312 15056
rect 11513 14998 12312 15000
rect 14089 15058 14155 15061
rect 15009 15058 15075 15061
rect 15377 15058 15443 15061
rect 14089 15056 15443 15058
rect 14089 15000 14094 15056
rect 14150 15000 15014 15056
rect 15070 15000 15382 15056
rect 15438 15000 15443 15056
rect 14089 14998 15443 15000
rect 11513 14995 11579 14998
rect 14089 14995 14155 14998
rect 15009 14995 15075 14998
rect 15377 14995 15443 14998
rect 16297 15058 16363 15061
rect 19934 15058 19994 15134
rect 22320 15104 22800 15134
rect 16297 15056 19994 15058
rect 16297 15000 16302 15056
rect 16358 15000 19994 15056
rect 16297 14998 19994 15000
rect 20069 15058 20135 15061
rect 20437 15058 20503 15061
rect 20069 15056 20503 15058
rect 20069 15000 20074 15056
rect 20130 15000 20442 15056
rect 20498 15000 20503 15056
rect 20069 14998 20503 15000
rect 16297 14995 16363 14998
rect 20069 14995 20135 14998
rect 20437 14995 20503 14998
rect 15469 14922 15535 14925
rect 18413 14922 18479 14925
rect 18873 14922 18939 14925
rect 15469 14920 18479 14922
rect 15469 14864 15474 14920
rect 15530 14864 18418 14920
rect 18474 14864 18479 14920
rect 15469 14862 18479 14864
rect 15469 14859 15535 14862
rect 18413 14859 18479 14862
rect 18600 14920 18939 14922
rect 18600 14864 18878 14920
rect 18934 14864 18939 14920
rect 18600 14862 18939 14864
rect 3417 14786 3483 14789
rect 0 14784 3483 14786
rect 0 14728 3422 14784
rect 3478 14728 3483 14784
rect 0 14726 3483 14728
rect 5030 14784 5139 14789
rect 5030 14728 5078 14784
rect 5134 14728 5139 14784
rect 5030 14726 5139 14728
rect 0 14696 480 14726
rect 3417 14723 3483 14726
rect 5073 14723 5139 14726
rect 17166 14724 17172 14788
rect 17236 14786 17242 14788
rect 17585 14786 17651 14789
rect 17236 14784 17651 14786
rect 17236 14728 17590 14784
rect 17646 14728 17651 14784
rect 17236 14726 17651 14728
rect 17236 14724 17242 14726
rect 17585 14723 17651 14726
rect 18137 14786 18203 14789
rect 18600 14786 18660 14862
rect 18873 14859 18939 14862
rect 18137 14784 18660 14786
rect 18137 14728 18142 14784
rect 18198 14728 18660 14784
rect 18137 14726 18660 14728
rect 18873 14786 18939 14789
rect 22320 14786 22800 14816
rect 18873 14784 22800 14786
rect 18873 14728 18878 14784
rect 18934 14728 22800 14784
rect 18873 14726 22800 14728
rect 18137 14723 18203 14726
rect 18873 14723 18939 14726
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 22320 14696 22800 14726
rect 14672 14655 14992 14656
rect 15694 14588 15700 14652
rect 15764 14650 15770 14652
rect 18822 14650 18828 14652
rect 15764 14590 18828 14650
rect 15764 14588 15770 14590
rect 18822 14588 18828 14590
rect 18892 14588 18898 14652
rect 19333 14650 19399 14653
rect 18968 14648 19399 14650
rect 18968 14592 19338 14648
rect 19394 14592 19399 14648
rect 18968 14590 19399 14592
rect 7557 14514 7623 14517
rect 7925 14514 7991 14517
rect 8334 14514 8340 14516
rect 7557 14512 8340 14514
rect 7557 14456 7562 14512
rect 7618 14456 7930 14512
rect 7986 14456 8340 14512
rect 7557 14454 8340 14456
rect 7557 14451 7623 14454
rect 7925 14451 7991 14454
rect 8334 14452 8340 14454
rect 8404 14452 8410 14516
rect 11421 14514 11487 14517
rect 11973 14514 12039 14517
rect 13077 14514 13143 14517
rect 11421 14512 13143 14514
rect 11421 14456 11426 14512
rect 11482 14456 11978 14512
rect 12034 14456 13082 14512
rect 13138 14456 13143 14512
rect 11421 14454 13143 14456
rect 11421 14451 11487 14454
rect 11973 14451 12039 14454
rect 13077 14451 13143 14454
rect 14641 14514 14707 14517
rect 15193 14514 15259 14517
rect 14641 14512 15259 14514
rect 14641 14456 14646 14512
rect 14702 14456 15198 14512
rect 15254 14456 15259 14512
rect 14641 14454 15259 14456
rect 14641 14451 14707 14454
rect 15193 14451 15259 14454
rect 16481 14514 16547 14517
rect 16614 14514 16620 14516
rect 16481 14512 16620 14514
rect 16481 14456 16486 14512
rect 16542 14456 16620 14512
rect 16481 14454 16620 14456
rect 16481 14451 16547 14454
rect 16614 14452 16620 14454
rect 16684 14452 16690 14516
rect 17534 14452 17540 14516
rect 17604 14514 17610 14516
rect 18229 14514 18295 14517
rect 17604 14512 18295 14514
rect 17604 14456 18234 14512
rect 18290 14456 18295 14512
rect 17604 14454 18295 14456
rect 17604 14452 17610 14454
rect 18229 14451 18295 14454
rect 18505 14514 18571 14517
rect 18968 14514 19028 14590
rect 19333 14587 19399 14590
rect 18505 14512 19028 14514
rect 18505 14456 18510 14512
rect 18566 14456 19028 14512
rect 18505 14454 19028 14456
rect 19333 14514 19399 14517
rect 19742 14514 19748 14516
rect 19333 14512 19748 14514
rect 19333 14456 19338 14512
rect 19394 14456 19748 14512
rect 19333 14454 19748 14456
rect 18505 14451 18571 14454
rect 19333 14451 19399 14454
rect 19742 14452 19748 14454
rect 19812 14452 19818 14516
rect 0 14378 480 14408
rect 1577 14378 1643 14381
rect 0 14376 1643 14378
rect 0 14320 1582 14376
rect 1638 14320 1643 14376
rect 0 14318 1643 14320
rect 0 14288 480 14318
rect 1577 14315 1643 14318
rect 5349 14378 5415 14381
rect 9070 14378 9076 14380
rect 5349 14376 9076 14378
rect 5349 14320 5354 14376
rect 5410 14320 9076 14376
rect 5349 14318 9076 14320
rect 5349 14315 5415 14318
rect 9070 14316 9076 14318
rect 9140 14316 9146 14380
rect 11094 14316 11100 14380
rect 11164 14378 11170 14380
rect 11513 14378 11579 14381
rect 11164 14376 11579 14378
rect 11164 14320 11518 14376
rect 11574 14320 11579 14376
rect 11164 14318 11579 14320
rect 11164 14316 11170 14318
rect 11513 14315 11579 14318
rect 12249 14378 12315 14381
rect 16941 14378 17007 14381
rect 12249 14376 17007 14378
rect 12249 14320 12254 14376
rect 12310 14320 16946 14376
rect 17002 14320 17007 14376
rect 12249 14318 17007 14320
rect 12249 14315 12315 14318
rect 16941 14315 17007 14318
rect 17677 14378 17743 14381
rect 22320 14378 22800 14408
rect 17677 14376 22800 14378
rect 17677 14320 17682 14376
rect 17738 14320 22800 14376
rect 17677 14318 22800 14320
rect 17677 14315 17743 14318
rect 22320 14288 22800 14318
rect 12525 14242 12591 14245
rect 16246 14242 16252 14244
rect 12525 14240 16252 14242
rect 12525 14184 12530 14240
rect 12586 14184 16252 14240
rect 12525 14182 16252 14184
rect 12525 14179 12591 14182
rect 16246 14180 16252 14182
rect 16316 14180 16322 14244
rect 18822 14180 18828 14244
rect 18892 14242 18898 14244
rect 19425 14242 19491 14245
rect 18892 14240 19491 14242
rect 18892 14184 19430 14240
rect 19486 14184 19491 14240
rect 18892 14182 19491 14184
rect 18892 14180 18898 14182
rect 19425 14179 19491 14182
rect 19742 14180 19748 14244
rect 19812 14242 19818 14244
rect 20161 14242 20227 14245
rect 19812 14240 20227 14242
rect 19812 14184 20166 14240
rect 20222 14184 20227 14240
rect 19812 14182 20227 14184
rect 19812 14180 19818 14182
rect 20161 14179 20227 14182
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 6085 14106 6151 14109
rect 8109 14106 8175 14109
rect 6085 14104 8175 14106
rect 6085 14048 6090 14104
rect 6146 14048 8114 14104
rect 8170 14048 8175 14104
rect 6085 14046 8175 14048
rect 6085 14043 6151 14046
rect 8109 14043 8175 14046
rect 12433 14106 12499 14109
rect 15561 14106 15627 14109
rect 12433 14104 15627 14106
rect 12433 14048 12438 14104
rect 12494 14048 15566 14104
rect 15622 14048 15627 14104
rect 12433 14046 15627 14048
rect 12433 14043 12499 14046
rect 15561 14043 15627 14046
rect 18646 14046 20362 14106
rect 0 13970 480 14000
rect 4245 13970 4311 13973
rect 0 13968 4311 13970
rect 0 13912 4250 13968
rect 4306 13912 4311 13968
rect 0 13910 4311 13912
rect 0 13880 480 13910
rect 4245 13907 4311 13910
rect 6177 13970 6243 13973
rect 11421 13970 11487 13973
rect 6177 13968 11487 13970
rect 6177 13912 6182 13968
rect 6238 13912 11426 13968
rect 11482 13912 11487 13968
rect 6177 13910 11487 13912
rect 6177 13907 6243 13910
rect 11421 13907 11487 13910
rect 15193 13970 15259 13973
rect 16297 13970 16363 13973
rect 15193 13968 16363 13970
rect 15193 13912 15198 13968
rect 15254 13912 16302 13968
rect 16358 13912 16363 13968
rect 15193 13910 16363 13912
rect 15193 13907 15259 13910
rect 16297 13907 16363 13910
rect 17677 13970 17743 13973
rect 18646 13970 18706 14046
rect 17677 13968 18706 13970
rect 17677 13912 17682 13968
rect 17738 13912 18706 13968
rect 17677 13910 18706 13912
rect 20302 13970 20362 14046
rect 22320 13970 22800 14000
rect 20302 13910 22800 13970
rect 17677 13907 17743 13910
rect 22320 13880 22800 13910
rect 2589 13834 2655 13837
rect 9438 13834 9444 13836
rect 2589 13832 9444 13834
rect 2589 13776 2594 13832
rect 2650 13776 9444 13832
rect 2589 13774 9444 13776
rect 2589 13771 2655 13774
rect 9438 13772 9444 13774
rect 9508 13772 9514 13836
rect 14641 13834 14707 13837
rect 18045 13834 18111 13837
rect 14641 13832 18111 13834
rect 14641 13776 14646 13832
rect 14702 13776 18050 13832
rect 18106 13776 18111 13832
rect 14641 13774 18111 13776
rect 14641 13771 14707 13774
rect 18045 13771 18111 13774
rect 20161 13834 20227 13837
rect 20529 13836 20595 13837
rect 20294 13834 20300 13836
rect 20161 13832 20300 13834
rect 20161 13776 20166 13832
rect 20222 13776 20300 13832
rect 20161 13774 20300 13776
rect 20161 13771 20227 13774
rect 20294 13772 20300 13774
rect 20364 13772 20370 13836
rect 20478 13834 20484 13836
rect 20438 13774 20484 13834
rect 20548 13832 20595 13836
rect 20590 13776 20595 13832
rect 20478 13772 20484 13774
rect 20548 13772 20595 13776
rect 20529 13771 20595 13772
rect 6729 13700 6795 13701
rect 6678 13636 6684 13700
rect 6748 13698 6795 13700
rect 9397 13698 9463 13701
rect 12249 13698 12315 13701
rect 6748 13696 6840 13698
rect 6790 13640 6840 13696
rect 6748 13638 6840 13640
rect 9397 13696 12315 13698
rect 9397 13640 9402 13696
rect 9458 13640 12254 13696
rect 12310 13640 12315 13696
rect 9397 13638 12315 13640
rect 6748 13636 6795 13638
rect 6729 13635 6795 13636
rect 9397 13635 9463 13638
rect 12249 13635 12315 13638
rect 18689 13698 18755 13701
rect 20897 13698 20963 13701
rect 18689 13696 20963 13698
rect 18689 13640 18694 13696
rect 18750 13640 20902 13696
rect 20958 13640 20963 13696
rect 18689 13638 20963 13640
rect 18689 13635 18755 13638
rect 20897 13635 20963 13638
rect 7808 13632 8128 13633
rect 0 13562 480 13592
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 1761 13562 1827 13565
rect 0 13560 1827 13562
rect 0 13504 1766 13560
rect 1822 13504 1827 13560
rect 0 13502 1827 13504
rect 0 13472 480 13502
rect 1761 13499 1827 13502
rect 11513 13562 11579 13565
rect 14406 13562 14412 13564
rect 11513 13560 14412 13562
rect 11513 13504 11518 13560
rect 11574 13504 14412 13560
rect 11513 13502 14412 13504
rect 11513 13499 11579 13502
rect 14406 13500 14412 13502
rect 14476 13500 14482 13564
rect 15929 13562 15995 13565
rect 16798 13562 16804 13564
rect 15929 13560 16804 13562
rect 15929 13504 15934 13560
rect 15990 13504 16804 13560
rect 15929 13502 16804 13504
rect 15929 13499 15995 13502
rect 16798 13500 16804 13502
rect 16868 13500 16874 13564
rect 17033 13560 17099 13565
rect 17033 13504 17038 13560
rect 17094 13504 17099 13560
rect 17033 13499 17099 13504
rect 18413 13562 18479 13565
rect 18873 13562 18939 13565
rect 18413 13560 18939 13562
rect 18413 13504 18418 13560
rect 18474 13504 18878 13560
rect 18934 13504 18939 13560
rect 18413 13502 18939 13504
rect 18413 13499 18479 13502
rect 18873 13499 18939 13502
rect 19241 13562 19307 13565
rect 22320 13562 22800 13592
rect 19241 13560 22800 13562
rect 19241 13504 19246 13560
rect 19302 13504 22800 13560
rect 19241 13502 22800 13504
rect 19241 13499 19307 13502
rect 6361 13426 6427 13429
rect 13169 13426 13235 13429
rect 6361 13424 13235 13426
rect 6361 13368 6366 13424
rect 6422 13368 13174 13424
rect 13230 13368 13235 13424
rect 6361 13366 13235 13368
rect 6361 13363 6427 13366
rect 13169 13363 13235 13366
rect 13353 13426 13419 13429
rect 17036 13426 17096 13499
rect 22320 13472 22800 13502
rect 18229 13426 18295 13429
rect 13353 13424 18295 13426
rect 13353 13368 13358 13424
rect 13414 13368 18234 13424
rect 18290 13368 18295 13424
rect 13353 13366 18295 13368
rect 13353 13363 13419 13366
rect 18229 13363 18295 13366
rect 1301 13290 1367 13293
rect 8937 13290 9003 13293
rect 1301 13288 9003 13290
rect 1301 13232 1306 13288
rect 1362 13232 8942 13288
rect 8998 13232 9003 13288
rect 1301 13230 9003 13232
rect 1301 13227 1367 13230
rect 8937 13227 9003 13230
rect 10317 13290 10383 13293
rect 16389 13290 16455 13293
rect 19742 13290 19748 13292
rect 10317 13288 16455 13290
rect 10317 13232 10322 13288
rect 10378 13232 16394 13288
rect 16450 13232 16455 13288
rect 10317 13230 16455 13232
rect 10317 13227 10383 13230
rect 16389 13227 16455 13230
rect 18646 13230 19748 13290
rect 0 13154 480 13184
rect 18646 13157 18706 13230
rect 19742 13228 19748 13230
rect 19812 13228 19818 13292
rect 2865 13154 2931 13157
rect 0 13152 2931 13154
rect 0 13096 2870 13152
rect 2926 13096 2931 13152
rect 0 13094 2931 13096
rect 0 13064 480 13094
rect 2865 13091 2931 13094
rect 13721 13154 13787 13157
rect 14641 13154 14707 13157
rect 13721 13152 14707 13154
rect 13721 13096 13726 13152
rect 13782 13096 14646 13152
rect 14702 13096 14707 13152
rect 13721 13094 14707 13096
rect 13721 13091 13787 13094
rect 14641 13091 14707 13094
rect 14825 13154 14891 13157
rect 15510 13154 15516 13156
rect 14825 13152 15516 13154
rect 14825 13096 14830 13152
rect 14886 13096 15516 13152
rect 14825 13094 15516 13096
rect 14825 13091 14891 13094
rect 15510 13092 15516 13094
rect 15580 13154 15586 13156
rect 16849 13154 16915 13157
rect 15580 13152 16915 13154
rect 15580 13096 16854 13152
rect 16910 13096 16915 13152
rect 15580 13094 16915 13096
rect 15580 13092 15586 13094
rect 16849 13091 16915 13094
rect 18597 13152 18706 13157
rect 18597 13096 18602 13152
rect 18658 13096 18706 13152
rect 18597 13094 18706 13096
rect 18781 13154 18847 13157
rect 22320 13154 22800 13184
rect 18781 13152 22800 13154
rect 18781 13096 18786 13152
rect 18842 13096 22800 13152
rect 18781 13094 22800 13096
rect 18597 13091 18663 13094
rect 18781 13091 18847 13094
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 22320 13064 22800 13094
rect 18104 13023 18424 13024
rect 10501 13018 10567 13021
rect 10726 13018 10732 13020
rect 10501 13016 10732 13018
rect 10501 12960 10506 13016
rect 10562 12960 10732 13016
rect 10501 12958 10732 12960
rect 10501 12955 10567 12958
rect 10726 12956 10732 12958
rect 10796 12956 10802 13020
rect 12709 13018 12775 13021
rect 16614 13018 16620 13020
rect 12709 13016 16620 13018
rect 12709 12960 12714 13016
rect 12770 12960 16620 13016
rect 12709 12958 16620 12960
rect 12709 12955 12775 12958
rect 16614 12956 16620 12958
rect 16684 12956 16690 13020
rect 19241 13016 19307 13021
rect 19241 12960 19246 13016
rect 19302 12960 19307 13016
rect 19241 12955 19307 12960
rect 10777 12882 10843 12885
rect 13353 12882 13419 12885
rect 10777 12880 13419 12882
rect 10777 12824 10782 12880
rect 10838 12824 13358 12880
rect 13414 12824 13419 12880
rect 10777 12822 13419 12824
rect 10777 12819 10843 12822
rect 13353 12819 13419 12822
rect 13629 12882 13695 12885
rect 17585 12884 17651 12885
rect 17534 12882 17540 12884
rect 13629 12880 17540 12882
rect 17604 12880 17651 12884
rect 19244 12882 19304 12955
rect 13629 12824 13634 12880
rect 13690 12824 17540 12880
rect 17646 12824 17651 12880
rect 13629 12822 17540 12824
rect 13629 12819 13695 12822
rect 17534 12820 17540 12822
rect 17604 12820 17651 12824
rect 17585 12819 17651 12820
rect 18784 12822 19304 12882
rect 0 12746 480 12776
rect 18784 12749 18844 12822
rect 4061 12746 4127 12749
rect 0 12744 4127 12746
rect 0 12688 4066 12744
rect 4122 12688 4127 12744
rect 0 12686 4127 12688
rect 0 12656 480 12686
rect 4061 12683 4127 12686
rect 5574 12684 5580 12748
rect 5644 12746 5650 12748
rect 5901 12746 5967 12749
rect 5644 12744 5967 12746
rect 5644 12688 5906 12744
rect 5962 12688 5967 12744
rect 5644 12686 5967 12688
rect 5644 12684 5650 12686
rect 5901 12683 5967 12686
rect 7281 12746 7347 12749
rect 14038 12746 14044 12748
rect 7281 12744 14044 12746
rect 7281 12688 7286 12744
rect 7342 12688 14044 12744
rect 7281 12686 14044 12688
rect 7281 12683 7347 12686
rect 14038 12684 14044 12686
rect 14108 12684 14114 12748
rect 14549 12746 14615 12749
rect 15832 12746 15838 12748
rect 14549 12744 15838 12746
rect 14549 12688 14554 12744
rect 14610 12688 15838 12744
rect 14549 12686 15838 12688
rect 14549 12683 14615 12686
rect 15832 12684 15838 12686
rect 15902 12684 15908 12748
rect 16205 12746 16271 12749
rect 16205 12744 17418 12746
rect 16205 12688 16210 12744
rect 16266 12688 17418 12744
rect 16205 12686 17418 12688
rect 16205 12683 16271 12686
rect 7005 12610 7071 12613
rect 7230 12610 7236 12612
rect 7005 12608 7236 12610
rect 7005 12552 7010 12608
rect 7066 12552 7236 12608
rect 7005 12550 7236 12552
rect 7005 12547 7071 12550
rect 7230 12548 7236 12550
rect 7300 12548 7306 12612
rect 10869 12608 10935 12613
rect 11881 12612 11947 12613
rect 10869 12552 10874 12608
rect 10930 12552 10935 12608
rect 10869 12547 10935 12552
rect 11830 12548 11836 12612
rect 11900 12610 11947 12612
rect 15469 12610 15535 12613
rect 16021 12610 16087 12613
rect 11900 12608 11992 12610
rect 11942 12552 11992 12608
rect 11900 12550 11992 12552
rect 15469 12608 16087 12610
rect 15469 12552 15474 12608
rect 15530 12552 16026 12608
rect 16082 12552 16087 12608
rect 15469 12550 16087 12552
rect 11900 12548 11947 12550
rect 11881 12547 11947 12548
rect 15469 12547 15535 12550
rect 16021 12547 16087 12550
rect 16246 12548 16252 12612
rect 16316 12610 16322 12612
rect 16389 12610 16455 12613
rect 16316 12608 16455 12610
rect 16316 12552 16394 12608
rect 16450 12552 16455 12608
rect 16316 12550 16455 12552
rect 17358 12610 17418 12686
rect 17534 12684 17540 12748
rect 17604 12746 17610 12748
rect 18638 12746 18644 12748
rect 17604 12686 18644 12746
rect 17604 12684 17610 12686
rect 18638 12684 18644 12686
rect 18708 12684 18714 12748
rect 18781 12744 18847 12749
rect 18781 12688 18786 12744
rect 18842 12688 18847 12744
rect 18781 12683 18847 12688
rect 19057 12746 19123 12749
rect 19333 12746 19399 12749
rect 22320 12746 22800 12776
rect 19057 12744 19399 12746
rect 19057 12688 19062 12744
rect 19118 12688 19338 12744
rect 19394 12688 19399 12744
rect 19057 12686 19399 12688
rect 19057 12683 19123 12686
rect 19333 12683 19399 12686
rect 19520 12686 22800 12746
rect 18638 12610 18644 12612
rect 17358 12550 18644 12610
rect 16316 12548 16322 12550
rect 16389 12547 16455 12550
rect 18638 12548 18644 12550
rect 18708 12548 18714 12612
rect 19057 12610 19123 12613
rect 19333 12610 19399 12613
rect 19057 12608 19399 12610
rect 19057 12552 19062 12608
rect 19118 12552 19338 12608
rect 19394 12552 19399 12608
rect 19057 12550 19399 12552
rect 19057 12547 19123 12550
rect 19333 12547 19399 12550
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 1209 12474 1275 12477
rect 7373 12474 7439 12477
rect 1209 12472 7439 12474
rect 1209 12416 1214 12472
rect 1270 12416 7378 12472
rect 7434 12416 7439 12472
rect 1209 12414 7439 12416
rect 1209 12411 1275 12414
rect 7373 12411 7439 12414
rect 8702 12412 8708 12476
rect 8772 12474 8778 12476
rect 9305 12474 9371 12477
rect 9581 12476 9647 12477
rect 9581 12474 9628 12476
rect 8772 12472 9371 12474
rect 8772 12416 9310 12472
rect 9366 12416 9371 12472
rect 8772 12414 9371 12416
rect 9540 12472 9628 12474
rect 9692 12474 9698 12476
rect 9540 12416 9586 12472
rect 9540 12414 9628 12416
rect 8772 12412 8778 12414
rect 9305 12411 9371 12414
rect 9581 12412 9628 12414
rect 9692 12414 9738 12474
rect 9692 12412 9698 12414
rect 9806 12412 9812 12476
rect 9876 12474 9882 12476
rect 9949 12474 10015 12477
rect 9876 12472 10015 12474
rect 9876 12416 9954 12472
rect 10010 12416 10015 12472
rect 9876 12414 10015 12416
rect 9876 12412 9882 12414
rect 9581 12411 9647 12412
rect 9949 12411 10015 12414
rect 10133 12476 10199 12477
rect 10133 12472 10180 12476
rect 10244 12474 10250 12476
rect 10133 12416 10138 12472
rect 10133 12412 10180 12416
rect 10244 12414 10290 12474
rect 10244 12412 10250 12414
rect 10133 12411 10199 12412
rect 0 12338 480 12368
rect 3141 12338 3207 12341
rect 7097 12338 7163 12341
rect 0 12336 3207 12338
rect 0 12280 3146 12336
rect 3202 12280 3207 12336
rect 0 12278 3207 12280
rect 0 12248 480 12278
rect 3141 12275 3207 12278
rect 7054 12336 7163 12338
rect 7054 12280 7102 12336
rect 7158 12280 7163 12336
rect 7054 12275 7163 12280
rect 7230 12276 7236 12340
rect 7300 12338 7306 12340
rect 7649 12338 7715 12341
rect 7300 12336 7715 12338
rect 7300 12280 7654 12336
rect 7710 12280 7715 12336
rect 7300 12278 7715 12280
rect 7300 12276 7306 12278
rect 7649 12275 7715 12278
rect 7925 12338 7991 12341
rect 9029 12338 9095 12341
rect 7925 12336 9095 12338
rect 7925 12280 7930 12336
rect 7986 12280 9034 12336
rect 9090 12280 9095 12336
rect 7925 12278 9095 12280
rect 7925 12275 7991 12278
rect 9029 12275 9095 12278
rect 10409 12338 10475 12341
rect 10872 12338 10932 12547
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 11145 12474 11211 12477
rect 12065 12474 12131 12477
rect 14181 12474 14247 12477
rect 11145 12472 12131 12474
rect 11145 12416 11150 12472
rect 11206 12416 12070 12472
rect 12126 12416 12131 12472
rect 11145 12414 12131 12416
rect 11145 12411 11211 12414
rect 12065 12411 12131 12414
rect 12252 12472 14247 12474
rect 12252 12416 14186 12472
rect 14242 12416 14247 12472
rect 12252 12414 14247 12416
rect 12252 12341 12312 12414
rect 14181 12411 14247 12414
rect 15469 12474 15535 12477
rect 16113 12474 16179 12477
rect 15469 12472 16179 12474
rect 15469 12416 15474 12472
rect 15530 12416 16118 12472
rect 16174 12416 16179 12472
rect 15469 12414 16179 12416
rect 15469 12411 15535 12414
rect 16113 12411 16179 12414
rect 16297 12474 16363 12477
rect 19520 12474 19580 12686
rect 22320 12656 22800 12686
rect 19885 12610 19951 12613
rect 20345 12610 20411 12613
rect 19885 12608 20411 12610
rect 19885 12552 19890 12608
rect 19946 12552 20350 12608
rect 20406 12552 20411 12608
rect 19885 12550 20411 12552
rect 19885 12547 19951 12550
rect 20345 12547 20411 12550
rect 19793 12476 19859 12477
rect 19742 12474 19748 12476
rect 16297 12472 19580 12474
rect 16297 12416 16302 12472
rect 16358 12416 19580 12472
rect 16297 12414 19580 12416
rect 19702 12414 19748 12474
rect 19812 12472 19859 12476
rect 19854 12416 19859 12472
rect 16297 12411 16363 12414
rect 19742 12412 19748 12414
rect 19812 12412 19859 12416
rect 19793 12411 19859 12412
rect 10409 12336 10932 12338
rect 10409 12280 10414 12336
rect 10470 12280 10932 12336
rect 10409 12278 10932 12280
rect 11881 12338 11947 12341
rect 12065 12338 12131 12341
rect 11881 12336 12131 12338
rect 11881 12280 11886 12336
rect 11942 12280 12070 12336
rect 12126 12280 12131 12336
rect 11881 12278 12131 12280
rect 10409 12275 10475 12278
rect 11881 12275 11947 12278
rect 12065 12275 12131 12278
rect 12249 12336 12315 12341
rect 12249 12280 12254 12336
rect 12310 12280 12315 12336
rect 12249 12275 12315 12280
rect 12985 12338 13051 12341
rect 13118 12338 13124 12340
rect 12985 12336 13124 12338
rect 12985 12280 12990 12336
rect 13046 12280 13124 12336
rect 12985 12278 13124 12280
rect 12985 12275 13051 12278
rect 13118 12276 13124 12278
rect 13188 12276 13194 12340
rect 13445 12338 13511 12341
rect 22320 12338 22800 12368
rect 13445 12336 22800 12338
rect 13445 12280 13450 12336
rect 13506 12280 22800 12336
rect 13445 12278 22800 12280
rect 13445 12275 13511 12278
rect 7054 12202 7114 12275
rect 22320 12248 22800 12278
rect 9305 12202 9371 12205
rect 7054 12200 9371 12202
rect 7054 12144 9310 12200
rect 9366 12144 9371 12200
rect 7054 12142 9371 12144
rect 9305 12139 9371 12142
rect 10041 12202 10107 12205
rect 10174 12202 10180 12204
rect 10041 12200 10180 12202
rect 10041 12144 10046 12200
rect 10102 12144 10180 12200
rect 10041 12142 10180 12144
rect 10041 12139 10107 12142
rect 10174 12140 10180 12142
rect 10244 12140 10250 12204
rect 10961 12202 11027 12205
rect 11830 12202 11836 12204
rect 10961 12200 11836 12202
rect 10961 12144 10966 12200
rect 11022 12144 11836 12200
rect 10961 12142 11836 12144
rect 10961 12139 11027 12142
rect 11830 12140 11836 12142
rect 11900 12140 11906 12204
rect 11973 12202 12039 12205
rect 14549 12202 14615 12205
rect 11973 12200 14615 12202
rect 11973 12144 11978 12200
rect 12034 12144 14554 12200
rect 14610 12144 14615 12200
rect 11973 12142 14615 12144
rect 11973 12139 12039 12142
rect 14549 12139 14615 12142
rect 15193 12202 15259 12205
rect 18413 12202 18479 12205
rect 15193 12200 18479 12202
rect 15193 12144 15198 12200
rect 15254 12144 18418 12200
rect 18474 12144 18479 12200
rect 15193 12142 18479 12144
rect 15193 12139 15259 12142
rect 18413 12139 18479 12142
rect 7465 12066 7531 12069
rect 8334 12066 8340 12068
rect 7465 12064 8340 12066
rect 7465 12008 7470 12064
rect 7526 12008 8340 12064
rect 7465 12006 8340 12008
rect 7465 12003 7531 12006
rect 8334 12004 8340 12006
rect 8404 12066 8410 12068
rect 8569 12066 8635 12069
rect 8404 12064 8635 12066
rect 8404 12008 8574 12064
rect 8630 12008 8635 12064
rect 8404 12006 8635 12008
rect 8404 12004 8410 12006
rect 8569 12003 8635 12006
rect 4376 12000 4696 12001
rect 0 11930 480 11960
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 3049 11930 3115 11933
rect 5349 11932 5415 11933
rect 5349 11930 5396 11932
rect 0 11928 3115 11930
rect 0 11872 3054 11928
rect 3110 11872 3115 11928
rect 0 11870 3115 11872
rect 5304 11928 5396 11930
rect 5304 11872 5354 11928
rect 5304 11870 5396 11872
rect 0 11840 480 11870
rect 3049 11867 3115 11870
rect 5349 11868 5396 11870
rect 5460 11868 5466 11932
rect 6637 11930 6703 11933
rect 10964 11930 11024 12139
rect 11697 12066 11763 12069
rect 11654 12064 11763 12066
rect 11654 12008 11702 12064
rect 11758 12008 11763 12064
rect 11654 12003 11763 12008
rect 12157 12066 12223 12069
rect 15326 12066 15332 12068
rect 12157 12064 15332 12066
rect 12157 12008 12162 12064
rect 12218 12008 15332 12064
rect 12157 12006 15332 12008
rect 12157 12003 12223 12006
rect 15326 12004 15332 12006
rect 15396 12066 15402 12068
rect 17861 12066 17927 12069
rect 15396 12064 17927 12066
rect 15396 12008 17866 12064
rect 17922 12008 17927 12064
rect 15396 12006 17927 12008
rect 15396 12004 15402 12006
rect 17861 12003 17927 12006
rect 18689 12066 18755 12069
rect 18822 12066 18828 12068
rect 18689 12064 18828 12066
rect 18689 12008 18694 12064
rect 18750 12008 18828 12064
rect 18689 12006 18828 12008
rect 18689 12003 18755 12006
rect 18822 12004 18828 12006
rect 18892 12004 18898 12068
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 6637 11928 11024 11930
rect 6637 11872 6642 11928
rect 6698 11872 11024 11928
rect 6637 11870 11024 11872
rect 5349 11867 5415 11868
rect 6637 11867 6703 11870
rect 1669 11794 1735 11797
rect 5901 11794 5967 11797
rect 1669 11792 5967 11794
rect 1669 11736 1674 11792
rect 1730 11736 5906 11792
rect 5962 11736 5967 11792
rect 1669 11734 5967 11736
rect 1669 11731 1735 11734
rect 5901 11731 5967 11734
rect 8293 11796 8359 11797
rect 8293 11792 8340 11796
rect 8404 11794 8410 11796
rect 10593 11794 10659 11797
rect 11654 11794 11714 12003
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 12985 11930 13051 11933
rect 11792 11928 13051 11930
rect 11792 11872 12990 11928
rect 13046 11872 13051 11928
rect 11792 11870 13051 11872
rect 11792 11797 11852 11870
rect 12985 11867 13051 11870
rect 13353 11930 13419 11933
rect 15694 11930 15700 11932
rect 13353 11928 15700 11930
rect 13353 11872 13358 11928
rect 13414 11872 15700 11928
rect 13353 11870 15700 11872
rect 13353 11867 13419 11870
rect 15694 11868 15700 11870
rect 15764 11930 15770 11932
rect 15837 11930 15903 11933
rect 15764 11928 15903 11930
rect 15764 11872 15842 11928
rect 15898 11872 15903 11928
rect 15764 11870 15903 11872
rect 15764 11868 15770 11870
rect 15837 11867 15903 11870
rect 16389 11930 16455 11933
rect 16614 11930 16620 11932
rect 16389 11928 16620 11930
rect 16389 11872 16394 11928
rect 16450 11872 16620 11928
rect 16389 11870 16620 11872
rect 16389 11867 16455 11870
rect 16614 11868 16620 11870
rect 16684 11868 16690 11932
rect 16757 11930 16823 11933
rect 16982 11930 16988 11932
rect 16757 11928 16988 11930
rect 16757 11872 16762 11928
rect 16818 11872 16988 11928
rect 16757 11870 16988 11872
rect 16757 11867 16823 11870
rect 16982 11868 16988 11870
rect 17052 11930 17058 11932
rect 17769 11930 17835 11933
rect 22320 11930 22800 11960
rect 17052 11928 17835 11930
rect 17052 11872 17774 11928
rect 17830 11872 17835 11928
rect 17052 11870 17835 11872
rect 17052 11868 17058 11870
rect 17769 11867 17835 11870
rect 18876 11870 22800 11930
rect 8293 11736 8298 11792
rect 8293 11732 8340 11736
rect 8404 11734 8450 11794
rect 10593 11792 11714 11794
rect 10593 11736 10598 11792
rect 10654 11736 11714 11792
rect 10593 11734 11714 11736
rect 11789 11792 11855 11797
rect 11789 11736 11794 11792
rect 11850 11736 11855 11792
rect 8404 11732 8410 11734
rect 8293 11731 8359 11732
rect 10593 11731 10659 11734
rect 11789 11731 11855 11736
rect 12249 11794 12315 11797
rect 12525 11794 12591 11797
rect 15469 11794 15535 11797
rect 12249 11792 15535 11794
rect 12249 11736 12254 11792
rect 12310 11736 12530 11792
rect 12586 11736 15474 11792
rect 15530 11736 15535 11792
rect 12249 11734 15535 11736
rect 12249 11731 12315 11734
rect 12525 11731 12591 11734
rect 15469 11731 15535 11734
rect 16573 11794 16639 11797
rect 16941 11794 17007 11797
rect 16573 11792 17007 11794
rect 16573 11736 16578 11792
rect 16634 11736 16946 11792
rect 17002 11736 17007 11792
rect 16573 11734 17007 11736
rect 16573 11731 16639 11734
rect 16941 11731 17007 11734
rect 17769 11794 17835 11797
rect 18876 11794 18936 11870
rect 22320 11840 22800 11870
rect 17769 11792 18936 11794
rect 17769 11736 17774 11792
rect 17830 11736 18936 11792
rect 17769 11734 18936 11736
rect 17769 11731 17835 11734
rect 0 11658 480 11688
rect 3877 11658 3943 11661
rect 0 11656 3943 11658
rect 0 11600 3882 11656
rect 3938 11600 3943 11656
rect 0 11598 3943 11600
rect 0 11568 480 11598
rect 3877 11595 3943 11598
rect 4889 11658 4955 11661
rect 7833 11658 7899 11661
rect 10041 11658 10107 11661
rect 13118 11658 13124 11660
rect 4889 11656 8264 11658
rect 4889 11600 4894 11656
rect 4950 11600 7838 11656
rect 7894 11600 8264 11656
rect 4889 11598 8264 11600
rect 4889 11595 4955 11598
rect 7833 11595 7899 11598
rect 4797 11524 4863 11525
rect 4797 11522 4844 11524
rect 4752 11520 4844 11522
rect 4752 11464 4802 11520
rect 4752 11462 4844 11464
rect 4797 11460 4844 11462
rect 4908 11460 4914 11524
rect 8204 11522 8264 11598
rect 10041 11656 13124 11658
rect 10041 11600 10046 11656
rect 10102 11600 13124 11656
rect 10041 11598 13124 11600
rect 10041 11595 10107 11598
rect 13118 11596 13124 11598
rect 13188 11596 13194 11660
rect 16573 11658 16639 11661
rect 14552 11656 16639 11658
rect 14552 11600 16578 11656
rect 16634 11600 16639 11656
rect 14552 11598 16639 11600
rect 10593 11522 10659 11525
rect 8204 11520 10659 11522
rect 8204 11464 10598 11520
rect 10654 11464 10659 11520
rect 8204 11462 10659 11464
rect 4797 11459 4863 11460
rect 10593 11459 10659 11462
rect 10726 11460 10732 11524
rect 10796 11522 10802 11524
rect 14552 11522 14612 11598
rect 16573 11595 16639 11598
rect 17677 11658 17743 11661
rect 22320 11658 22800 11688
rect 17677 11656 22800 11658
rect 17677 11600 17682 11656
rect 17738 11600 22800 11656
rect 17677 11598 22800 11600
rect 17677 11595 17743 11598
rect 22320 11568 22800 11598
rect 10796 11462 14612 11522
rect 15101 11522 15167 11525
rect 16113 11524 16179 11525
rect 15326 11522 15332 11524
rect 15101 11520 15332 11522
rect 15101 11464 15106 11520
rect 15162 11464 15332 11520
rect 15101 11462 15332 11464
rect 10796 11460 10802 11462
rect 15101 11459 15167 11462
rect 15326 11460 15332 11462
rect 15396 11460 15402 11524
rect 16062 11522 16068 11524
rect 16022 11462 16068 11522
rect 16132 11520 16179 11524
rect 16174 11464 16179 11520
rect 16062 11460 16068 11462
rect 16132 11460 16179 11464
rect 16246 11460 16252 11524
rect 16316 11522 16322 11524
rect 16481 11522 16547 11525
rect 16316 11520 16547 11522
rect 16316 11464 16486 11520
rect 16542 11464 16547 11520
rect 16316 11462 16547 11464
rect 16316 11460 16322 11462
rect 16113 11459 16179 11460
rect 16481 11459 16547 11462
rect 16798 11460 16804 11524
rect 16868 11522 16874 11524
rect 17953 11522 18019 11525
rect 16868 11520 18019 11522
rect 16868 11464 17958 11520
rect 18014 11464 18019 11520
rect 16868 11462 18019 11464
rect 16868 11460 16874 11462
rect 17953 11459 18019 11462
rect 18873 11522 18939 11525
rect 19926 11522 19932 11524
rect 18873 11520 19932 11522
rect 18873 11464 18878 11520
rect 18934 11464 19932 11520
rect 18873 11462 19932 11464
rect 18873 11459 18939 11462
rect 19926 11460 19932 11462
rect 19996 11460 20002 11524
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 8845 11386 8911 11389
rect 9254 11386 9260 11388
rect 8845 11384 9260 11386
rect 8845 11328 8850 11384
rect 8906 11328 9260 11384
rect 8845 11326 9260 11328
rect 8845 11323 8911 11326
rect 9254 11324 9260 11326
rect 9324 11324 9330 11388
rect 9397 11386 9463 11389
rect 12249 11386 12315 11389
rect 9397 11384 12315 11386
rect 9397 11328 9402 11384
rect 9458 11328 12254 11384
rect 12310 11328 12315 11384
rect 9397 11326 12315 11328
rect 9397 11323 9463 11326
rect 12249 11323 12315 11326
rect 12617 11386 12683 11389
rect 12750 11386 12756 11388
rect 12617 11384 12756 11386
rect 12617 11328 12622 11384
rect 12678 11328 12756 11384
rect 12617 11326 12756 11328
rect 12617 11323 12683 11326
rect 12750 11324 12756 11326
rect 12820 11324 12826 11388
rect 13670 11324 13676 11388
rect 13740 11386 13746 11388
rect 14181 11386 14247 11389
rect 14365 11386 14431 11389
rect 13740 11384 14431 11386
rect 13740 11328 14186 11384
rect 14242 11328 14370 11384
rect 14426 11328 14431 11384
rect 13740 11326 14431 11328
rect 13740 11324 13746 11326
rect 14181 11323 14247 11326
rect 14365 11323 14431 11326
rect 15561 11386 15627 11389
rect 16389 11386 16455 11389
rect 15561 11384 16455 11386
rect 15561 11328 15566 11384
rect 15622 11328 16394 11384
rect 16450 11328 16455 11384
rect 15561 11326 16455 11328
rect 15561 11323 15627 11326
rect 16389 11323 16455 11326
rect 17861 11386 17927 11389
rect 19057 11386 19123 11389
rect 17861 11384 19123 11386
rect 17861 11328 17866 11384
rect 17922 11328 19062 11384
rect 19118 11328 19123 11384
rect 17861 11326 19123 11328
rect 17861 11323 17927 11326
rect 19057 11323 19123 11326
rect 0 11250 480 11280
rect 1577 11250 1643 11253
rect 0 11248 1643 11250
rect 0 11192 1582 11248
rect 1638 11192 1643 11248
rect 0 11190 1643 11192
rect 0 11160 480 11190
rect 1577 11187 1643 11190
rect 3509 11250 3575 11253
rect 6453 11250 6519 11253
rect 3509 11248 6519 11250
rect 3509 11192 3514 11248
rect 3570 11192 6458 11248
rect 6514 11192 6519 11248
rect 3509 11190 6519 11192
rect 3509 11187 3575 11190
rect 6453 11187 6519 11190
rect 8937 11250 9003 11253
rect 13537 11250 13603 11253
rect 13997 11250 14063 11253
rect 18137 11250 18203 11253
rect 8937 11248 13603 11250
rect 8937 11192 8942 11248
rect 8998 11192 13542 11248
rect 13598 11192 13603 11248
rect 8937 11190 13603 11192
rect 8937 11187 9003 11190
rect 13537 11187 13603 11190
rect 13724 11248 14063 11250
rect 13724 11192 14002 11248
rect 14058 11192 14063 11248
rect 14414 11248 18203 11250
rect 14414 11216 18142 11248
rect 13724 11190 14063 11192
rect 2998 11052 3004 11116
rect 3068 11114 3074 11116
rect 7741 11114 7807 11117
rect 8201 11114 8267 11117
rect 12382 11114 12388 11116
rect 3068 11112 8034 11114
rect 3068 11056 7746 11112
rect 7802 11056 8034 11112
rect 3068 11054 8034 11056
rect 3068 11052 3074 11054
rect 7741 11051 7807 11054
rect 5533 10980 5599 10981
rect 5533 10978 5580 10980
rect 5488 10976 5580 10978
rect 5488 10920 5538 10976
rect 5488 10918 5580 10920
rect 5533 10916 5580 10918
rect 5644 10916 5650 10980
rect 7974 10978 8034 11054
rect 8201 11112 12388 11114
rect 8201 11056 8206 11112
rect 8262 11056 12388 11112
rect 8201 11054 12388 11056
rect 8201 11051 8267 11054
rect 12382 11052 12388 11054
rect 12452 11052 12458 11116
rect 12801 11114 12867 11117
rect 13724 11114 13784 11190
rect 13997 11187 14063 11190
rect 14230 11192 18142 11216
rect 18198 11192 18203 11248
rect 14230 11190 18203 11192
rect 14230 11156 14474 11190
rect 18137 11187 18203 11190
rect 20897 11250 20963 11253
rect 22320 11250 22800 11280
rect 20897 11248 22800 11250
rect 20897 11192 20902 11248
rect 20958 11192 22800 11248
rect 20897 11190 22800 11192
rect 20897 11187 20963 11190
rect 22320 11160 22800 11190
rect 12801 11112 13784 11114
rect 12801 11056 12806 11112
rect 12862 11056 13784 11112
rect 12801 11054 13784 11056
rect 13905 11114 13971 11117
rect 14230 11114 14290 11156
rect 13905 11112 14290 11114
rect 13905 11056 13910 11112
rect 13966 11056 14290 11112
rect 13905 11054 14290 11056
rect 14549 11114 14615 11117
rect 15653 11114 15719 11117
rect 21265 11114 21331 11117
rect 14549 11112 15719 11114
rect 14549 11056 14554 11112
rect 14610 11056 15658 11112
rect 15714 11056 15719 11112
rect 14549 11054 15719 11056
rect 12801 11051 12867 11054
rect 13905 11051 13971 11054
rect 14549 11051 14615 11054
rect 15653 11051 15719 11054
rect 16944 11112 21331 11114
rect 16944 11056 21270 11112
rect 21326 11056 21331 11112
rect 16944 11054 21331 11056
rect 10685 10978 10751 10981
rect 7974 10976 10751 10978
rect 7974 10920 10690 10976
rect 10746 10920 10751 10976
rect 7974 10918 10751 10920
rect 5533 10915 5599 10916
rect 10685 10915 10751 10918
rect 12985 10978 13051 10981
rect 13997 10978 14063 10981
rect 12985 10976 14063 10978
rect 12985 10920 12990 10976
rect 13046 10920 14002 10976
rect 14058 10920 14063 10976
rect 12985 10918 14063 10920
rect 12985 10915 13051 10918
rect 13997 10915 14063 10918
rect 14181 10978 14247 10981
rect 16757 10978 16823 10981
rect 14181 10976 16823 10978
rect 14181 10920 14186 10976
rect 14242 10920 16762 10976
rect 16818 10920 16823 10976
rect 14181 10918 16823 10920
rect 14181 10915 14247 10918
rect 16757 10915 16823 10918
rect 4376 10912 4696 10913
rect 0 10842 480 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 9213 10842 9279 10845
rect 0 10782 4216 10842
rect 0 10752 480 10782
rect 4156 10706 4216 10782
rect 4800 10840 9279 10842
rect 4800 10784 9218 10840
rect 9274 10784 9279 10840
rect 4800 10782 9279 10784
rect 4800 10706 4860 10782
rect 9213 10779 9279 10782
rect 10133 10844 10199 10845
rect 10133 10840 10180 10844
rect 10244 10842 10250 10844
rect 12065 10842 12131 10845
rect 12198 10842 12204 10844
rect 10133 10784 10138 10840
rect 10133 10780 10180 10784
rect 10244 10782 10290 10842
rect 12065 10840 12204 10842
rect 12065 10784 12070 10840
rect 12126 10784 12204 10840
rect 12065 10782 12204 10784
rect 10244 10780 10250 10782
rect 10133 10779 10199 10780
rect 12065 10779 12131 10782
rect 12198 10780 12204 10782
rect 12268 10780 12274 10844
rect 12433 10842 12499 10845
rect 16944 10842 17004 11054
rect 21265 11051 21331 11054
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 12433 10840 17004 10842
rect 12433 10784 12438 10840
rect 12494 10784 17004 10840
rect 12433 10782 17004 10784
rect 12433 10779 12499 10782
rect 18638 10780 18644 10844
rect 18708 10842 18714 10844
rect 22320 10842 22800 10872
rect 18708 10782 22800 10842
rect 18708 10780 18714 10782
rect 22320 10752 22800 10782
rect 4156 10646 4860 10706
rect 5206 10644 5212 10708
rect 5276 10706 5282 10708
rect 5349 10706 5415 10709
rect 5276 10704 5415 10706
rect 5276 10648 5354 10704
rect 5410 10648 5415 10704
rect 5276 10646 5415 10648
rect 5276 10644 5282 10646
rect 5349 10643 5415 10646
rect 5625 10706 5691 10709
rect 5758 10706 5764 10708
rect 5625 10704 5764 10706
rect 5625 10648 5630 10704
rect 5686 10648 5764 10704
rect 5625 10646 5764 10648
rect 5625 10643 5691 10646
rect 5758 10644 5764 10646
rect 5828 10644 5834 10708
rect 6085 10706 6151 10709
rect 8845 10706 8911 10709
rect 17534 10706 17540 10708
rect 6085 10704 8911 10706
rect 6085 10648 6090 10704
rect 6146 10648 8850 10704
rect 8906 10648 8911 10704
rect 6085 10646 8911 10648
rect 6085 10643 6151 10646
rect 8845 10643 8911 10646
rect 9078 10646 17540 10706
rect 3550 10508 3556 10572
rect 3620 10570 3626 10572
rect 9078 10570 9138 10646
rect 17534 10644 17540 10646
rect 17604 10706 17610 10708
rect 18413 10706 18479 10709
rect 17604 10704 18479 10706
rect 17604 10648 18418 10704
rect 18474 10648 18479 10704
rect 17604 10646 18479 10648
rect 17604 10644 17610 10646
rect 18413 10643 18479 10646
rect 3620 10510 9138 10570
rect 9213 10570 9279 10573
rect 16297 10570 16363 10573
rect 9213 10568 16363 10570
rect 9213 10512 9218 10568
rect 9274 10512 16302 10568
rect 16358 10512 16363 10568
rect 9213 10510 16363 10512
rect 3620 10508 3626 10510
rect 9213 10507 9279 10510
rect 16297 10507 16363 10510
rect 17309 10570 17375 10573
rect 19742 10570 19748 10572
rect 17309 10568 19748 10570
rect 17309 10512 17314 10568
rect 17370 10512 19748 10568
rect 17309 10510 19748 10512
rect 17309 10507 17375 10510
rect 19742 10508 19748 10510
rect 19812 10508 19818 10572
rect 0 10434 480 10464
rect 5901 10434 5967 10437
rect 8385 10436 8451 10437
rect 0 10432 5967 10434
rect 0 10376 5906 10432
rect 5962 10376 5967 10432
rect 0 10374 5967 10376
rect 0 10344 480 10374
rect 5901 10371 5967 10374
rect 8334 10372 8340 10436
rect 8404 10434 8451 10436
rect 8661 10436 8727 10437
rect 9029 10436 9095 10437
rect 8661 10434 8708 10436
rect 8404 10432 8496 10434
rect 8446 10376 8496 10432
rect 8404 10374 8496 10376
rect 8616 10432 8708 10434
rect 8616 10376 8666 10432
rect 8616 10374 8708 10376
rect 8404 10372 8451 10374
rect 8385 10371 8451 10372
rect 8661 10372 8708 10374
rect 8772 10372 8778 10436
rect 9029 10432 9076 10436
rect 9140 10434 9146 10436
rect 9397 10434 9463 10437
rect 9622 10434 9628 10436
rect 9029 10376 9034 10432
rect 9029 10372 9076 10376
rect 9140 10374 9186 10434
rect 9397 10432 9628 10434
rect 9397 10376 9402 10432
rect 9458 10376 9628 10432
rect 9397 10374 9628 10376
rect 9140 10372 9146 10374
rect 8661 10371 8727 10372
rect 9029 10371 9095 10372
rect 9397 10371 9463 10374
rect 9622 10372 9628 10374
rect 9692 10372 9698 10436
rect 12198 10372 12204 10436
rect 12268 10434 12274 10436
rect 12934 10434 12940 10436
rect 12268 10374 12940 10434
rect 12268 10372 12274 10374
rect 12934 10372 12940 10374
rect 13004 10372 13010 10436
rect 13537 10434 13603 10437
rect 14457 10434 14523 10437
rect 13537 10432 14523 10434
rect 13537 10376 13542 10432
rect 13598 10376 14462 10432
rect 14518 10376 14523 10432
rect 13537 10374 14523 10376
rect 13537 10371 13603 10374
rect 14457 10371 14523 10374
rect 15377 10434 15443 10437
rect 15510 10434 15516 10436
rect 15377 10432 15516 10434
rect 15377 10376 15382 10432
rect 15438 10376 15516 10432
rect 15377 10374 15516 10376
rect 15377 10371 15443 10374
rect 15510 10372 15516 10374
rect 15580 10372 15586 10436
rect 17861 10434 17927 10437
rect 22320 10434 22800 10464
rect 17861 10432 22800 10434
rect 17861 10376 17866 10432
rect 17922 10376 22800 10432
rect 17861 10374 22800 10376
rect 17861 10371 17927 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 22320 10344 22800 10374
rect 14672 10303 14992 10304
rect 4889 10300 4955 10301
rect 4838 10298 4844 10300
rect 4798 10238 4844 10298
rect 4908 10296 4955 10300
rect 4950 10240 4955 10296
rect 4838 10236 4844 10238
rect 4908 10236 4955 10240
rect 4889 10235 4955 10236
rect 6085 10298 6151 10301
rect 6821 10298 6887 10301
rect 7005 10300 7071 10301
rect 7005 10298 7052 10300
rect 6085 10296 6887 10298
rect 6085 10240 6090 10296
rect 6146 10240 6826 10296
rect 6882 10240 6887 10296
rect 6085 10238 6887 10240
rect 6960 10296 7052 10298
rect 6960 10240 7010 10296
rect 6960 10238 7052 10240
rect 6085 10235 6151 10238
rect 6821 10235 6887 10238
rect 7005 10236 7052 10238
rect 7116 10236 7122 10300
rect 8569 10298 8635 10301
rect 17309 10298 17375 10301
rect 19885 10298 19951 10301
rect 8569 10296 13876 10298
rect 8569 10240 8574 10296
rect 8630 10240 13876 10296
rect 8569 10238 13876 10240
rect 7005 10235 7071 10236
rect 8569 10235 8635 10238
rect 2037 10162 2103 10165
rect 7833 10162 7899 10165
rect 13816 10162 13876 10238
rect 17309 10296 19951 10298
rect 17309 10240 17314 10296
rect 17370 10240 19890 10296
rect 19946 10240 19951 10296
rect 17309 10238 19951 10240
rect 17309 10235 17375 10238
rect 19885 10235 19951 10238
rect 15653 10162 15719 10165
rect 2037 10160 7666 10162
rect 2037 10104 2042 10160
rect 2098 10104 7666 10160
rect 2037 10102 7666 10104
rect 2037 10099 2103 10102
rect 0 10026 480 10056
rect 1301 10026 1367 10029
rect 0 10024 1367 10026
rect 0 9968 1306 10024
rect 1362 9968 1367 10024
rect 0 9966 1367 9968
rect 0 9936 480 9966
rect 1301 9963 1367 9966
rect 3233 10026 3299 10029
rect 7465 10026 7531 10029
rect 3233 10024 7531 10026
rect 3233 9968 3238 10024
rect 3294 9968 7470 10024
rect 7526 9968 7531 10024
rect 3233 9966 7531 9968
rect 7606 10026 7666 10102
rect 7833 10160 13738 10162
rect 7833 10104 7838 10160
rect 7894 10104 13738 10160
rect 7833 10102 13738 10104
rect 13816 10160 15719 10162
rect 13816 10104 15658 10160
rect 15714 10104 15719 10160
rect 13816 10102 15719 10104
rect 7833 10099 7899 10102
rect 13537 10026 13603 10029
rect 7606 10024 13603 10026
rect 7606 9968 13542 10024
rect 13598 9968 13603 10024
rect 7606 9966 13603 9968
rect 13678 10026 13738 10102
rect 15653 10099 15719 10102
rect 16205 10162 16271 10165
rect 16430 10162 16436 10164
rect 16205 10160 16436 10162
rect 16205 10104 16210 10160
rect 16266 10104 16436 10160
rect 16205 10102 16436 10104
rect 16205 10099 16271 10102
rect 16430 10100 16436 10102
rect 16500 10100 16506 10164
rect 20989 10162 21055 10165
rect 17358 10160 21055 10162
rect 17358 10104 20994 10160
rect 21050 10104 21055 10160
rect 17358 10102 21055 10104
rect 17217 10026 17283 10029
rect 13678 10024 17283 10026
rect 13678 9968 17222 10024
rect 17278 9968 17283 10024
rect 13678 9966 17283 9968
rect 3233 9963 3299 9966
rect 7465 9963 7531 9966
rect 13537 9963 13603 9966
rect 17217 9963 17283 9966
rect 7230 9828 7236 9892
rect 7300 9890 7306 9892
rect 9806 9890 9812 9892
rect 7300 9830 9812 9890
rect 7300 9828 7306 9830
rect 9806 9828 9812 9830
rect 9876 9828 9882 9892
rect 10593 9890 10659 9893
rect 11094 9890 11100 9892
rect 10593 9888 11100 9890
rect 10593 9832 10598 9888
rect 10654 9832 11100 9888
rect 10593 9830 11100 9832
rect 10593 9827 10659 9830
rect 11094 9828 11100 9830
rect 11164 9828 11170 9892
rect 12065 9890 12131 9893
rect 17358 9890 17418 10102
rect 20989 10099 21055 10102
rect 20621 10026 20687 10029
rect 22320 10026 22800 10056
rect 12065 9888 17418 9890
rect 12065 9832 12070 9888
rect 12126 9832 17418 9888
rect 12065 9830 17418 9832
rect 17496 10024 22800 10026
rect 17496 9968 20626 10024
rect 20682 9968 22800 10024
rect 17496 9966 22800 9968
rect 12065 9827 12131 9830
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 9857 9754 9923 9757
rect 4846 9752 9923 9754
rect 4846 9696 9862 9752
rect 9918 9696 9923 9752
rect 4846 9694 9923 9696
rect 0 9618 480 9648
rect 4846 9618 4906 9694
rect 9857 9691 9923 9694
rect 10174 9692 10180 9756
rect 10244 9754 10250 9756
rect 10501 9754 10567 9757
rect 12014 9754 12020 9756
rect 10244 9752 10567 9754
rect 10244 9696 10506 9752
rect 10562 9696 10567 9752
rect 10244 9694 10567 9696
rect 10244 9692 10250 9694
rect 10501 9691 10567 9694
rect 11654 9694 12020 9754
rect 5073 9618 5139 9621
rect 0 9558 4906 9618
rect 5030 9616 5139 9618
rect 5030 9560 5078 9616
rect 5134 9560 5139 9616
rect 0 9528 480 9558
rect 5030 9555 5139 9560
rect 6637 9618 6703 9621
rect 7230 9618 7236 9620
rect 6637 9616 7236 9618
rect 6637 9560 6642 9616
rect 6698 9560 7236 9616
rect 6637 9558 7236 9560
rect 6637 9555 6703 9558
rect 7230 9556 7236 9558
rect 7300 9556 7306 9620
rect 7465 9618 7531 9621
rect 11513 9618 11579 9621
rect 11654 9618 11714 9694
rect 12014 9692 12020 9694
rect 12084 9692 12090 9756
rect 12249 9754 12315 9757
rect 17496 9754 17556 9966
rect 20621 9963 20687 9966
rect 22320 9936 22800 9966
rect 18822 9828 18828 9892
rect 18892 9890 18898 9892
rect 20161 9890 20227 9893
rect 18892 9888 20227 9890
rect 18892 9832 20166 9888
rect 20222 9832 20227 9888
rect 18892 9830 20227 9832
rect 18892 9828 18898 9830
rect 20161 9827 20227 9830
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 12249 9752 17556 9754
rect 12249 9696 12254 9752
rect 12310 9696 17556 9752
rect 12249 9694 17556 9696
rect 12249 9691 12315 9694
rect 7465 9616 11714 9618
rect 7465 9560 7470 9616
rect 7526 9560 11518 9616
rect 11574 9560 11714 9616
rect 7465 9558 11714 9560
rect 11973 9618 12039 9621
rect 13854 9618 13860 9620
rect 11973 9616 13860 9618
rect 11973 9560 11978 9616
rect 12034 9560 13860 9616
rect 11973 9558 13860 9560
rect 7465 9555 7531 9558
rect 11513 9555 11579 9558
rect 11973 9555 12039 9558
rect 13854 9556 13860 9558
rect 13924 9556 13930 9620
rect 14917 9618 14983 9621
rect 15837 9618 15903 9621
rect 16021 9618 16087 9621
rect 14917 9616 16087 9618
rect 14917 9560 14922 9616
rect 14978 9560 15842 9616
rect 15898 9560 16026 9616
rect 16082 9560 16087 9616
rect 14917 9558 16087 9560
rect 14917 9555 14983 9558
rect 15837 9555 15903 9558
rect 16021 9555 16087 9558
rect 16389 9618 16455 9621
rect 17217 9618 17283 9621
rect 16389 9616 17283 9618
rect 16389 9560 16394 9616
rect 16450 9560 17222 9616
rect 17278 9560 17283 9616
rect 16389 9558 17283 9560
rect 16389 9555 16455 9558
rect 17217 9555 17283 9558
rect 17585 9618 17651 9621
rect 22320 9618 22800 9648
rect 17585 9616 22800 9618
rect 17585 9560 17590 9616
rect 17646 9560 22800 9616
rect 17585 9558 22800 9560
rect 17585 9555 17651 9558
rect 4797 9482 4863 9485
rect 5030 9482 5090 9555
rect 22320 9528 22800 9558
rect 4797 9480 5090 9482
rect 4797 9424 4802 9480
rect 4858 9424 5090 9480
rect 4797 9422 5090 9424
rect 6269 9484 6335 9485
rect 6269 9480 6316 9484
rect 6380 9482 6386 9484
rect 6269 9424 6274 9480
rect 4797 9419 4863 9422
rect 6269 9420 6316 9424
rect 6380 9422 6426 9482
rect 6380 9420 6386 9422
rect 6862 9420 6868 9484
rect 6932 9482 6938 9484
rect 8017 9482 8083 9485
rect 8937 9482 9003 9485
rect 6932 9480 9003 9482
rect 6932 9424 8022 9480
rect 8078 9424 8942 9480
rect 8998 9424 9003 9480
rect 6932 9422 9003 9424
rect 6932 9420 6938 9422
rect 6269 9419 6335 9420
rect 8017 9419 8083 9422
rect 8937 9419 9003 9422
rect 10174 9420 10180 9484
rect 10244 9482 10250 9484
rect 10409 9482 10475 9485
rect 13486 9482 13492 9484
rect 10244 9480 10475 9482
rect 10244 9424 10414 9480
rect 10470 9424 10475 9480
rect 10244 9422 10475 9424
rect 10244 9420 10250 9422
rect 10409 9419 10475 9422
rect 10550 9422 13492 9482
rect 10550 9349 10610 9422
rect 13486 9420 13492 9422
rect 13556 9420 13562 9484
rect 13905 9482 13971 9485
rect 16113 9482 16179 9485
rect 13905 9480 16179 9482
rect 13905 9424 13910 9480
rect 13966 9424 16118 9480
rect 16174 9424 16179 9480
rect 13905 9422 16179 9424
rect 13905 9419 13971 9422
rect 16113 9419 16179 9422
rect 16297 9482 16363 9485
rect 17033 9482 17099 9485
rect 16297 9480 17099 9482
rect 16297 9424 16302 9480
rect 16358 9424 17038 9480
rect 17094 9424 17099 9480
rect 16297 9422 17099 9424
rect 16297 9419 16363 9422
rect 17033 9419 17099 9422
rect 3693 9346 3759 9349
rect 3918 9346 3924 9348
rect 3693 9344 3924 9346
rect 3693 9288 3698 9344
rect 3754 9288 3924 9344
rect 3693 9286 3924 9288
rect 3693 9283 3759 9286
rect 3918 9284 3924 9286
rect 3988 9284 3994 9348
rect 5165 9346 5231 9349
rect 4064 9344 5231 9346
rect 4064 9288 5170 9344
rect 5226 9288 5231 9344
rect 4064 9286 5231 9288
rect 0 9210 480 9240
rect 4064 9210 4124 9286
rect 5165 9283 5231 9286
rect 10501 9344 10610 9349
rect 10501 9288 10506 9344
rect 10562 9288 10610 9344
rect 10501 9286 10610 9288
rect 11605 9346 11671 9349
rect 13670 9346 13676 9348
rect 11605 9344 13676 9346
rect 11605 9288 11610 9344
rect 11666 9288 13676 9344
rect 11605 9286 13676 9288
rect 10501 9283 10567 9286
rect 11605 9283 11671 9286
rect 13670 9284 13676 9286
rect 13740 9284 13746 9348
rect 15561 9346 15627 9349
rect 16389 9346 16455 9349
rect 15561 9344 16455 9346
rect 15561 9288 15566 9344
rect 15622 9288 16394 9344
rect 16450 9288 16455 9344
rect 15561 9286 16455 9288
rect 15561 9283 15627 9286
rect 16389 9283 16455 9286
rect 16941 9346 17007 9349
rect 19885 9346 19951 9349
rect 16941 9344 19951 9346
rect 16941 9288 16946 9344
rect 17002 9288 19890 9344
rect 19946 9288 19951 9344
rect 16941 9286 19951 9288
rect 16941 9283 17007 9286
rect 19885 9283 19951 9286
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 0 9150 4124 9210
rect 8385 9210 8451 9213
rect 10593 9210 10659 9213
rect 8385 9208 10659 9210
rect 8385 9152 8390 9208
rect 8446 9152 10598 9208
rect 10654 9152 10659 9208
rect 8385 9150 10659 9152
rect 0 9120 480 9150
rect 8385 9147 8451 9150
rect 10593 9147 10659 9150
rect 11145 9210 11211 9213
rect 12198 9210 12204 9212
rect 11145 9208 12204 9210
rect 11145 9152 11150 9208
rect 11206 9152 12204 9208
rect 11145 9150 12204 9152
rect 11145 9147 11211 9150
rect 12198 9148 12204 9150
rect 12268 9148 12274 9212
rect 13445 9210 13511 9213
rect 14365 9210 14431 9213
rect 13445 9208 14431 9210
rect 13445 9152 13450 9208
rect 13506 9152 14370 9208
rect 14426 9152 14431 9208
rect 13445 9150 14431 9152
rect 13445 9147 13511 9150
rect 14365 9147 14431 9150
rect 15193 9210 15259 9213
rect 16573 9210 16639 9213
rect 22320 9210 22800 9240
rect 15193 9208 16498 9210
rect 15193 9152 15198 9208
rect 15254 9152 16498 9208
rect 15193 9150 16498 9152
rect 15193 9147 15259 9150
rect 16438 9077 16498 9150
rect 16573 9208 22800 9210
rect 16573 9152 16578 9208
rect 16634 9152 22800 9208
rect 16573 9150 22800 9152
rect 16573 9147 16639 9150
rect 22320 9120 22800 9150
rect 3693 9074 3759 9077
rect 7189 9074 7255 9077
rect 15561 9074 15627 9077
rect 15745 9074 15811 9077
rect 3693 9072 7068 9074
rect 3693 9016 3698 9072
rect 3754 9016 7068 9072
rect 3693 9014 7068 9016
rect 3693 9011 3759 9014
rect 4705 8938 4771 8941
rect 4156 8936 4771 8938
rect 4156 8880 4710 8936
rect 4766 8880 4771 8936
rect 4156 8878 4771 8880
rect 0 8802 480 8832
rect 4156 8802 4216 8878
rect 4705 8875 4771 8878
rect 5349 8938 5415 8941
rect 5574 8938 5580 8940
rect 5349 8936 5580 8938
rect 5349 8880 5354 8936
rect 5410 8880 5580 8936
rect 5349 8878 5580 8880
rect 5349 8875 5415 8878
rect 5574 8876 5580 8878
rect 5644 8876 5650 8940
rect 7008 8938 7068 9014
rect 7189 9072 15811 9074
rect 7189 9016 7194 9072
rect 7250 9016 15566 9072
rect 15622 9016 15750 9072
rect 15806 9016 15811 9072
rect 7189 9014 15811 9016
rect 16438 9072 16547 9077
rect 16438 9016 16486 9072
rect 16542 9016 16547 9072
rect 16438 9014 16547 9016
rect 7189 9011 7255 9014
rect 15561 9011 15627 9014
rect 15745 9011 15811 9014
rect 16481 9011 16547 9014
rect 17953 9074 18019 9077
rect 18321 9074 18387 9077
rect 18505 9074 18571 9077
rect 20713 9074 20779 9077
rect 17953 9072 18571 9074
rect 17953 9016 17958 9072
rect 18014 9016 18326 9072
rect 18382 9016 18510 9072
rect 18566 9016 18571 9072
rect 17953 9014 18571 9016
rect 17953 9011 18019 9014
rect 18321 9011 18387 9014
rect 18505 9011 18571 9014
rect 20670 9072 20779 9074
rect 20670 9016 20718 9072
rect 20774 9016 20779 9072
rect 20670 9011 20779 9016
rect 9070 8938 9076 8940
rect 7008 8878 9076 8938
rect 9070 8876 9076 8878
rect 9140 8938 9146 8940
rect 11329 8938 11395 8941
rect 9140 8936 11395 8938
rect 9140 8880 11334 8936
rect 11390 8880 11395 8936
rect 9140 8878 11395 8880
rect 9140 8876 9146 8878
rect 11329 8875 11395 8878
rect 11513 8938 11579 8941
rect 11789 8938 11855 8941
rect 12617 8938 12683 8941
rect 12934 8938 12940 8940
rect 11513 8936 11714 8938
rect 11513 8880 11518 8936
rect 11574 8880 11714 8936
rect 11513 8878 11714 8880
rect 11513 8875 11579 8878
rect 9029 8802 9095 8805
rect 0 8742 4216 8802
rect 4984 8800 9095 8802
rect 4984 8744 9034 8800
rect 9090 8744 9095 8800
rect 4984 8742 9095 8744
rect 0 8712 480 8742
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 4984 8669 5044 8742
rect 9029 8739 9095 8742
rect 9438 8740 9444 8804
rect 9508 8802 9514 8804
rect 11094 8802 11100 8804
rect 9508 8742 11100 8802
rect 9508 8740 9514 8742
rect 11094 8740 11100 8742
rect 11164 8740 11170 8804
rect 11654 8802 11714 8878
rect 11789 8936 12036 8938
rect 11789 8880 11794 8936
rect 11850 8880 12036 8936
rect 11789 8878 12036 8880
rect 11789 8875 11855 8878
rect 11789 8802 11855 8805
rect 11654 8800 11855 8802
rect 11654 8744 11794 8800
rect 11850 8744 11855 8800
rect 11654 8742 11855 8744
rect 11976 8802 12036 8878
rect 12617 8936 12940 8938
rect 12617 8880 12622 8936
rect 12678 8880 12940 8936
rect 12617 8878 12940 8880
rect 12617 8875 12683 8878
rect 12934 8876 12940 8878
rect 13004 8938 13010 8940
rect 19609 8938 19675 8941
rect 20670 8938 20730 9011
rect 13004 8936 20730 8938
rect 13004 8880 19614 8936
rect 19670 8880 20730 8936
rect 13004 8878 20730 8880
rect 13004 8876 13010 8878
rect 19609 8875 19675 8878
rect 12985 8802 13051 8805
rect 11976 8800 13051 8802
rect 11976 8744 12990 8800
rect 13046 8744 13051 8800
rect 11976 8742 13051 8744
rect 11789 8739 11855 8742
rect 12985 8739 13051 8742
rect 15561 8802 15627 8805
rect 16297 8802 16363 8805
rect 15561 8800 16363 8802
rect 15561 8744 15566 8800
rect 15622 8744 16302 8800
rect 16358 8744 16363 8800
rect 15561 8742 16363 8744
rect 15561 8739 15627 8742
rect 16297 8739 16363 8742
rect 18505 8802 18571 8805
rect 22320 8802 22800 8832
rect 18505 8800 22800 8802
rect 18505 8744 18510 8800
rect 18566 8744 22800 8800
rect 18505 8742 22800 8744
rect 18505 8739 18571 8742
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 22320 8712 22800 8742
rect 18104 8671 18424 8672
rect 1485 8666 1551 8669
rect 4245 8666 4311 8669
rect 1485 8664 4311 8666
rect 1485 8608 1490 8664
rect 1546 8608 4250 8664
rect 4306 8608 4311 8664
rect 1485 8606 4311 8608
rect 1485 8603 1551 8606
rect 4245 8603 4311 8606
rect 4981 8664 5047 8669
rect 4981 8608 4986 8664
rect 5042 8608 5047 8664
rect 4981 8603 5047 8608
rect 7465 8666 7531 8669
rect 8293 8666 8359 8669
rect 7465 8664 8359 8666
rect 7465 8608 7470 8664
rect 7526 8608 8298 8664
rect 8354 8608 8359 8664
rect 7465 8606 8359 8608
rect 7465 8603 7531 8606
rect 8293 8603 8359 8606
rect 8569 8666 8635 8669
rect 8886 8666 8892 8668
rect 8569 8664 8892 8666
rect 8569 8608 8574 8664
rect 8630 8608 8892 8664
rect 8569 8606 8892 8608
rect 8569 8603 8635 8606
rect 8886 8604 8892 8606
rect 8956 8604 8962 8668
rect 11973 8666 12039 8669
rect 12249 8666 12315 8669
rect 16757 8666 16823 8669
rect 11973 8664 16823 8666
rect 11973 8608 11978 8664
rect 12034 8608 12254 8664
rect 12310 8608 16762 8664
rect 16818 8608 16823 8664
rect 11973 8606 16823 8608
rect 11973 8603 12039 8606
rect 12249 8603 12315 8606
rect 16757 8603 16823 8606
rect 2773 8530 2839 8533
rect 13721 8530 13787 8533
rect 14641 8530 14707 8533
rect 2773 8528 14707 8530
rect 2773 8472 2778 8528
rect 2834 8472 13726 8528
rect 13782 8472 14646 8528
rect 14702 8472 14707 8528
rect 2773 8470 14707 8472
rect 2773 8467 2839 8470
rect 13721 8467 13787 8470
rect 14641 8467 14707 8470
rect 16481 8530 16547 8533
rect 20989 8530 21055 8533
rect 16481 8528 21055 8530
rect 16481 8472 16486 8528
rect 16542 8472 20994 8528
rect 21050 8472 21055 8528
rect 16481 8470 21055 8472
rect 16481 8467 16547 8470
rect 20989 8467 21055 8470
rect 0 8394 480 8424
rect 11145 8394 11211 8397
rect 0 8392 11211 8394
rect 0 8336 11150 8392
rect 11206 8336 11211 8392
rect 0 8334 11211 8336
rect 0 8304 480 8334
rect 11145 8331 11211 8334
rect 11973 8396 12039 8397
rect 11973 8392 12020 8396
rect 12084 8394 12090 8396
rect 12801 8394 12867 8397
rect 16062 8394 16068 8396
rect 11973 8336 11978 8392
rect 11973 8332 12020 8336
rect 12084 8334 12130 8394
rect 12801 8392 16068 8394
rect 12801 8336 12806 8392
rect 12862 8336 16068 8392
rect 12801 8334 16068 8336
rect 12084 8332 12090 8334
rect 11973 8331 12039 8332
rect 12801 8331 12867 8334
rect 16062 8332 16068 8334
rect 16132 8332 16138 8396
rect 16757 8394 16823 8397
rect 22320 8394 22800 8424
rect 16757 8392 22800 8394
rect 16757 8336 16762 8392
rect 16818 8336 22800 8392
rect 16757 8334 22800 8336
rect 16757 8331 16823 8334
rect 22320 8304 22800 8334
rect 5390 8196 5396 8260
rect 5460 8258 5466 8260
rect 6453 8258 6519 8261
rect 5460 8256 6519 8258
rect 5460 8200 6458 8256
rect 6514 8200 6519 8256
rect 5460 8198 6519 8200
rect 5460 8196 5466 8198
rect 6453 8195 6519 8198
rect 8334 8196 8340 8260
rect 8404 8258 8410 8260
rect 10685 8258 10751 8261
rect 14273 8258 14339 8261
rect 18689 8260 18755 8261
rect 8404 8256 10751 8258
rect 8404 8200 10690 8256
rect 10746 8200 10751 8256
rect 8404 8198 10751 8200
rect 8404 8196 8410 8198
rect 10685 8195 10751 8198
rect 10872 8256 14339 8258
rect 10872 8200 14278 8256
rect 14334 8200 14339 8256
rect 10872 8198 14339 8200
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 8702 8060 8708 8124
rect 8772 8122 8778 8124
rect 9489 8122 9555 8125
rect 8772 8120 9555 8122
rect 8772 8064 9494 8120
rect 9550 8064 9555 8120
rect 8772 8062 9555 8064
rect 8772 8060 8778 8062
rect 9489 8059 9555 8062
rect 0 7986 480 8016
rect 6177 7986 6243 7989
rect 0 7984 6243 7986
rect 0 7928 6182 7984
rect 6238 7928 6243 7984
rect 0 7926 6243 7928
rect 0 7896 480 7926
rect 6177 7923 6243 7926
rect 6453 7986 6519 7989
rect 10542 7986 10548 7988
rect 6453 7984 10548 7986
rect 6453 7928 6458 7984
rect 6514 7928 10548 7984
rect 6453 7926 10548 7928
rect 6453 7923 6519 7926
rect 10542 7924 10548 7926
rect 10612 7924 10618 7988
rect 4429 7850 4495 7853
rect 7649 7850 7715 7853
rect 9305 7850 9371 7853
rect 10872 7850 10932 8198
rect 14273 8195 14339 8198
rect 18638 8196 18644 8260
rect 18708 8258 18755 8260
rect 18708 8256 18800 8258
rect 18750 8200 18800 8256
rect 18708 8198 18800 8200
rect 18708 8196 18755 8198
rect 18689 8195 18755 8196
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 11053 8122 11119 8125
rect 13905 8122 13971 8125
rect 11053 8120 13971 8122
rect 11053 8064 11058 8120
rect 11114 8064 13910 8120
rect 13966 8064 13971 8120
rect 11053 8062 13971 8064
rect 11053 8059 11119 8062
rect 13905 8059 13971 8062
rect 17401 8122 17467 8125
rect 18781 8122 18847 8125
rect 17401 8120 18847 8122
rect 17401 8064 17406 8120
rect 17462 8064 18786 8120
rect 18842 8064 18847 8120
rect 17401 8062 18847 8064
rect 17401 8059 17467 8062
rect 18781 8059 18847 8062
rect 16573 7986 16639 7989
rect 22320 7986 22800 8016
rect 4429 7848 4906 7850
rect 4429 7792 4434 7848
rect 4490 7792 4906 7848
rect 4429 7790 4906 7792
rect 4429 7787 4495 7790
rect 0 7714 480 7744
rect 3969 7714 4035 7717
rect 0 7712 4035 7714
rect 0 7656 3974 7712
rect 4030 7656 4035 7712
rect 0 7654 4035 7656
rect 4846 7714 4906 7790
rect 7649 7848 10932 7850
rect 7649 7792 7654 7848
rect 7710 7792 9310 7848
rect 9366 7792 10932 7848
rect 7649 7790 10932 7792
rect 11102 7984 22800 7986
rect 11102 7928 16578 7984
rect 16634 7928 22800 7984
rect 11102 7926 22800 7928
rect 7649 7787 7715 7790
rect 9305 7787 9371 7790
rect 5165 7714 5231 7717
rect 11102 7714 11162 7926
rect 16573 7923 16639 7926
rect 22320 7896 22800 7926
rect 11237 7850 11303 7853
rect 16849 7850 16915 7853
rect 11237 7848 16915 7850
rect 11237 7792 11242 7848
rect 11298 7792 16854 7848
rect 16910 7792 16915 7848
rect 18048 7816 19258 7850
rect 11237 7790 16915 7792
rect 11237 7787 11303 7790
rect 16849 7787 16915 7790
rect 17910 7790 19442 7816
rect 17910 7756 18108 7790
rect 19198 7756 19442 7790
rect 4846 7712 11162 7714
rect 4846 7656 5170 7712
rect 5226 7656 11162 7712
rect 4846 7654 11162 7656
rect 13721 7714 13787 7717
rect 13721 7712 14336 7714
rect 13721 7656 13726 7712
rect 13782 7656 14336 7712
rect 13721 7654 14336 7656
rect 0 7624 480 7654
rect 3969 7651 4035 7654
rect 5165 7651 5231 7654
rect 13721 7651 13787 7654
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 6177 7578 6243 7581
rect 8845 7578 8911 7581
rect 9397 7578 9463 7581
rect 6177 7576 9463 7578
rect 6177 7520 6182 7576
rect 6238 7520 8850 7576
rect 8906 7520 9402 7576
rect 9458 7520 9463 7576
rect 6177 7518 9463 7520
rect 6177 7515 6243 7518
rect 8845 7515 8911 7518
rect 9397 7515 9463 7518
rect 10317 7578 10383 7581
rect 10961 7578 11027 7581
rect 10317 7576 11027 7578
rect 10317 7520 10322 7576
rect 10378 7520 10966 7576
rect 11022 7520 11027 7576
rect 10317 7518 11027 7520
rect 10317 7515 10383 7518
rect 10961 7515 11027 7518
rect 11830 7516 11836 7580
rect 11900 7578 11906 7580
rect 13077 7578 13143 7581
rect 14089 7580 14155 7581
rect 11900 7576 13143 7578
rect 11900 7520 13082 7576
rect 13138 7520 13143 7576
rect 11900 7518 13143 7520
rect 11900 7516 11906 7518
rect 13077 7515 13143 7518
rect 14038 7516 14044 7580
rect 14108 7578 14155 7580
rect 14276 7578 14336 7654
rect 14406 7652 14412 7716
rect 14476 7714 14482 7716
rect 17910 7714 17970 7756
rect 14476 7654 17970 7714
rect 19382 7714 19442 7756
rect 22320 7714 22800 7744
rect 19382 7654 22800 7714
rect 14476 7652 14482 7654
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 22320 7624 22800 7654
rect 18104 7583 18424 7584
rect 15745 7578 15811 7581
rect 14108 7576 14200 7578
rect 14150 7520 14200 7576
rect 14108 7518 14200 7520
rect 14276 7576 15811 7578
rect 14276 7520 15750 7576
rect 15806 7520 15811 7576
rect 14276 7518 15811 7520
rect 14108 7516 14155 7518
rect 14089 7515 14155 7516
rect 15745 7515 15811 7518
rect 4705 7442 4771 7445
rect 7281 7442 7347 7445
rect 4705 7440 7347 7442
rect 4705 7384 4710 7440
rect 4766 7384 7286 7440
rect 7342 7384 7347 7440
rect 4705 7382 7347 7384
rect 4705 7379 4771 7382
rect 7281 7379 7347 7382
rect 7598 7380 7604 7444
rect 7668 7442 7674 7444
rect 11053 7442 11119 7445
rect 18229 7442 18295 7445
rect 7668 7440 11119 7442
rect 7668 7384 11058 7440
rect 11114 7384 11119 7440
rect 7668 7382 11119 7384
rect 7668 7380 7674 7382
rect 11053 7379 11119 7382
rect 11286 7440 18295 7442
rect 11286 7384 18234 7440
rect 18290 7384 18295 7440
rect 11286 7382 18295 7384
rect 0 7306 480 7336
rect 6361 7306 6427 7309
rect 0 7304 6427 7306
rect 0 7248 6366 7304
rect 6422 7248 6427 7304
rect 0 7246 6427 7248
rect 0 7216 480 7246
rect 6361 7243 6427 7246
rect 7046 7244 7052 7308
rect 7116 7306 7122 7308
rect 7414 7306 7420 7308
rect 7116 7246 7420 7306
rect 7116 7244 7122 7246
rect 7414 7244 7420 7246
rect 7484 7306 7490 7308
rect 8845 7306 8911 7309
rect 11145 7306 11211 7309
rect 7484 7246 8264 7306
rect 7484 7244 7490 7246
rect 1761 7170 1827 7173
rect 7230 7170 7236 7172
rect 1761 7168 7236 7170
rect 1761 7112 1766 7168
rect 1822 7112 7236 7168
rect 1761 7110 7236 7112
rect 1761 7107 1827 7110
rect 7230 7108 7236 7110
rect 7300 7108 7306 7172
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 6637 7034 6703 7037
rect 8204 7034 8264 7246
rect 8845 7304 11211 7306
rect 8845 7248 8850 7304
rect 8906 7248 11150 7304
rect 11206 7248 11211 7304
rect 8845 7246 11211 7248
rect 8845 7243 8911 7246
rect 11145 7243 11211 7246
rect 8518 7108 8524 7172
rect 8588 7170 8594 7172
rect 11286 7170 11346 7382
rect 18229 7379 18295 7382
rect 11513 7306 11579 7309
rect 12065 7306 12131 7309
rect 11513 7304 12131 7306
rect 11513 7248 11518 7304
rect 11574 7248 12070 7304
rect 12126 7248 12131 7304
rect 11513 7246 12131 7248
rect 11513 7243 11579 7246
rect 12065 7243 12131 7246
rect 12985 7306 13051 7309
rect 15837 7306 15903 7309
rect 12985 7304 15903 7306
rect 12985 7248 12990 7304
rect 13046 7248 15842 7304
rect 15898 7248 15903 7304
rect 12985 7246 15903 7248
rect 12985 7243 13051 7246
rect 15837 7243 15903 7246
rect 16062 7244 16068 7308
rect 16132 7306 16138 7308
rect 22320 7306 22800 7336
rect 16132 7246 22800 7306
rect 16132 7244 16138 7246
rect 14365 7170 14431 7173
rect 8588 7110 11346 7170
rect 11424 7168 14431 7170
rect 11424 7112 14370 7168
rect 14426 7112 14431 7168
rect 11424 7110 14431 7112
rect 8588 7108 8594 7110
rect 11424 7034 11484 7110
rect 13678 7037 13738 7110
rect 14365 7107 14431 7110
rect 15285 7170 15351 7173
rect 16070 7170 16130 7244
rect 22320 7216 22800 7246
rect 15285 7168 16130 7170
rect 15285 7112 15290 7168
rect 15346 7112 16130 7168
rect 15285 7110 16130 7112
rect 16205 7170 16271 7173
rect 18781 7170 18847 7173
rect 19190 7170 19196 7172
rect 16205 7168 19196 7170
rect 16205 7112 16210 7168
rect 16266 7112 18786 7168
rect 18842 7112 19196 7168
rect 16205 7110 19196 7112
rect 15285 7107 15351 7110
rect 16205 7107 16271 7110
rect 18781 7107 18847 7110
rect 19190 7108 19196 7110
rect 19260 7108 19266 7172
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 6637 7032 7482 7034
rect 6637 6976 6642 7032
rect 6698 6976 7482 7032
rect 6637 6974 7482 6976
rect 8204 6974 11484 7034
rect 12893 7034 12959 7037
rect 13118 7034 13124 7036
rect 12893 7032 13124 7034
rect 12893 6976 12898 7032
rect 12954 6976 13124 7032
rect 12893 6974 13124 6976
rect 6637 6971 6703 6974
rect 0 6898 480 6928
rect 7422 6898 7482 6974
rect 12893 6971 12959 6974
rect 13118 6972 13124 6974
rect 13188 6972 13194 7036
rect 13629 7032 13738 7037
rect 13629 6976 13634 7032
rect 13690 6976 13738 7032
rect 13629 6974 13738 6976
rect 18321 7034 18387 7037
rect 18822 7034 18828 7036
rect 18321 7032 18828 7034
rect 18321 6976 18326 7032
rect 18382 6976 18828 7032
rect 18321 6974 18828 6976
rect 13629 6971 13695 6974
rect 18321 6971 18387 6974
rect 18822 6972 18828 6974
rect 18892 6972 18898 7036
rect 11237 6898 11303 6901
rect 0 6838 1410 6898
rect 7422 6896 11303 6898
rect 7422 6840 11242 6896
rect 11298 6840 11303 6896
rect 7422 6838 11303 6840
rect 0 6808 480 6838
rect 1350 6626 1410 6838
rect 11237 6835 11303 6838
rect 12893 6898 12959 6901
rect 18505 6898 18571 6901
rect 12893 6896 18571 6898
rect 12893 6840 12898 6896
rect 12954 6840 18510 6896
rect 18566 6840 18571 6896
rect 12893 6838 18571 6840
rect 12893 6835 12959 6838
rect 18505 6835 18571 6838
rect 19149 6898 19215 6901
rect 22320 6898 22800 6928
rect 19149 6896 22800 6898
rect 19149 6840 19154 6896
rect 19210 6840 22800 6896
rect 19149 6838 22800 6840
rect 19149 6835 19215 6838
rect 22320 6808 22800 6838
rect 1761 6762 1827 6765
rect 3417 6762 3483 6765
rect 1761 6760 3483 6762
rect 1761 6704 1766 6760
rect 1822 6704 3422 6760
rect 3478 6704 3483 6760
rect 1761 6702 3483 6704
rect 1761 6699 1827 6702
rect 3417 6699 3483 6702
rect 3601 6762 3667 6765
rect 16205 6762 16271 6765
rect 3601 6760 16271 6762
rect 3601 6704 3606 6760
rect 3662 6704 16210 6760
rect 16266 6704 16271 6760
rect 3601 6702 16271 6704
rect 3601 6699 3667 6702
rect 16205 6699 16271 6702
rect 16481 6762 16547 6765
rect 18321 6762 18387 6765
rect 16481 6760 18387 6762
rect 16481 6704 16486 6760
rect 16542 6704 18326 6760
rect 18382 6704 18387 6760
rect 16481 6702 18387 6704
rect 16481 6699 16547 6702
rect 18321 6699 18387 6702
rect 3969 6626 4035 6629
rect 1350 6624 4035 6626
rect 1350 6568 3974 6624
rect 4030 6568 4035 6624
rect 1350 6566 4035 6568
rect 3969 6563 4035 6566
rect 5441 6626 5507 6629
rect 11053 6626 11119 6629
rect 5441 6624 11119 6626
rect 5441 6568 5446 6624
rect 5502 6568 11058 6624
rect 11114 6568 11119 6624
rect 5441 6566 11119 6568
rect 5441 6563 5507 6566
rect 11053 6563 11119 6566
rect 13118 6564 13124 6628
rect 13188 6626 13194 6628
rect 14917 6626 14983 6629
rect 13188 6624 14983 6626
rect 13188 6568 14922 6624
rect 14978 6568 14983 6624
rect 13188 6566 14983 6568
rect 13188 6564 13194 6566
rect 14917 6563 14983 6566
rect 15101 6626 15167 6629
rect 17309 6626 17375 6629
rect 15101 6624 17375 6626
rect 15101 6568 15106 6624
rect 15162 6568 17314 6624
rect 17370 6568 17375 6624
rect 15101 6566 17375 6568
rect 15101 6563 15167 6566
rect 17309 6563 17375 6566
rect 4376 6560 4696 6561
rect 0 6490 480 6520
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 4245 6490 4311 6493
rect 0 6488 4311 6490
rect 0 6432 4250 6488
rect 4306 6432 4311 6488
rect 0 6430 4311 6432
rect 0 6400 480 6430
rect 4245 6427 4311 6430
rect 5717 6490 5783 6493
rect 7649 6490 7715 6493
rect 10358 6490 10364 6492
rect 5717 6488 7715 6490
rect 5717 6432 5722 6488
rect 5778 6432 7654 6488
rect 7710 6432 7715 6488
rect 5717 6430 7715 6432
rect 5717 6427 5783 6430
rect 7649 6427 7715 6430
rect 7790 6430 10364 6490
rect 1577 6354 1643 6357
rect 7790 6354 7850 6430
rect 10358 6428 10364 6430
rect 10428 6428 10434 6492
rect 11881 6490 11947 6493
rect 15193 6490 15259 6493
rect 22320 6490 22800 6520
rect 11881 6488 15259 6490
rect 11881 6432 11886 6488
rect 11942 6432 15198 6488
rect 15254 6432 15259 6488
rect 19382 6456 22800 6490
rect 11881 6430 15259 6432
rect 11881 6427 11947 6430
rect 15193 6427 15259 6430
rect 19198 6430 22800 6456
rect 19198 6396 19442 6430
rect 22320 6400 22800 6430
rect 1577 6352 7850 6354
rect 1577 6296 1582 6352
rect 1638 6296 7850 6352
rect 1577 6294 7850 6296
rect 7925 6354 7991 6357
rect 8569 6354 8635 6357
rect 7925 6352 8635 6354
rect 7925 6296 7930 6352
rect 7986 6296 8574 6352
rect 8630 6296 8635 6352
rect 7925 6294 8635 6296
rect 1577 6291 1643 6294
rect 7925 6291 7991 6294
rect 8569 6291 8635 6294
rect 9397 6354 9463 6357
rect 14089 6354 14155 6357
rect 9397 6352 14155 6354
rect 9397 6296 9402 6352
rect 9458 6296 14094 6352
rect 14150 6296 14155 6352
rect 9397 6294 14155 6296
rect 9397 6291 9463 6294
rect 14089 6291 14155 6294
rect 14917 6354 14983 6357
rect 19198 6354 19258 6396
rect 14917 6352 19258 6354
rect 14917 6296 14922 6352
rect 14978 6296 19258 6352
rect 14917 6294 19258 6296
rect 14917 6291 14983 6294
rect 5073 6218 5139 6221
rect 5717 6218 5783 6221
rect 8569 6218 8635 6221
rect 5073 6216 5783 6218
rect 5073 6160 5078 6216
rect 5134 6160 5722 6216
rect 5778 6160 5783 6216
rect 5073 6158 5783 6160
rect 5073 6155 5139 6158
rect 5717 6155 5783 6158
rect 6456 6158 8264 6218
rect 0 6082 480 6112
rect 6456 6082 6516 6158
rect 0 6022 6516 6082
rect 6637 6082 6703 6085
rect 6862 6082 6868 6084
rect 6637 6080 6868 6082
rect 6637 6024 6642 6080
rect 6698 6024 6868 6080
rect 6637 6022 6868 6024
rect 0 5992 480 6022
rect 6637 6019 6703 6022
rect 6862 6020 6868 6022
rect 6932 6020 6938 6084
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 4705 5946 4771 5949
rect 6545 5946 6611 5949
rect 4705 5944 6611 5946
rect 4705 5888 4710 5944
rect 4766 5888 6550 5944
rect 6606 5888 6611 5944
rect 4705 5886 6611 5888
rect 4705 5883 4771 5886
rect 6545 5883 6611 5886
rect 6821 5946 6887 5949
rect 7189 5946 7255 5949
rect 6821 5944 7255 5946
rect 6821 5888 6826 5944
rect 6882 5888 7194 5944
rect 7250 5888 7255 5944
rect 6821 5886 7255 5888
rect 8204 5946 8264 6158
rect 8569 6216 17234 6218
rect 8569 6160 8574 6216
rect 8630 6160 17234 6216
rect 8569 6158 17234 6160
rect 8569 6155 8635 6158
rect 9581 6082 9647 6085
rect 10501 6082 10567 6085
rect 9581 6080 10567 6082
rect 9581 6024 9586 6080
rect 9642 6024 10506 6080
rect 10562 6024 10567 6080
rect 9581 6022 10567 6024
rect 9581 6019 9647 6022
rect 10501 6019 10567 6022
rect 10777 6082 10843 6085
rect 11830 6082 11836 6084
rect 10777 6080 11836 6082
rect 10777 6024 10782 6080
rect 10838 6024 11836 6080
rect 10777 6022 11836 6024
rect 10777 6019 10843 6022
rect 11830 6020 11836 6022
rect 11900 6020 11906 6084
rect 12433 6082 12499 6085
rect 12566 6082 12572 6084
rect 12433 6080 12572 6082
rect 12433 6024 12438 6080
rect 12494 6024 12572 6080
rect 12433 6022 12572 6024
rect 12433 6019 12499 6022
rect 12566 6020 12572 6022
rect 12636 6082 12642 6084
rect 13905 6082 13971 6085
rect 12636 6080 13971 6082
rect 12636 6024 13910 6080
rect 13966 6024 13971 6080
rect 12636 6022 13971 6024
rect 17174 6082 17234 6158
rect 22320 6082 22800 6112
rect 17174 6022 22800 6082
rect 12636 6020 12642 6022
rect 13905 6019 13971 6022
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 22320 5992 22800 6022
rect 14672 5951 14992 5952
rect 8569 5946 8635 5949
rect 12617 5946 12683 5949
rect 8204 5944 12683 5946
rect 8204 5888 8574 5944
rect 8630 5888 12622 5944
rect 12678 5888 12683 5944
rect 8204 5886 12683 5888
rect 6821 5883 6887 5886
rect 7189 5883 7255 5886
rect 8569 5883 8635 5886
rect 12617 5883 12683 5886
rect 17033 5946 17099 5949
rect 17677 5946 17743 5949
rect 18137 5946 18203 5949
rect 17033 5944 18203 5946
rect 17033 5888 17038 5944
rect 17094 5888 17682 5944
rect 17738 5888 18142 5944
rect 18198 5888 18203 5944
rect 17033 5886 18203 5888
rect 17033 5883 17099 5886
rect 17677 5883 17743 5886
rect 18137 5883 18203 5886
rect 19742 5884 19748 5948
rect 19812 5946 19818 5948
rect 19885 5946 19951 5949
rect 19812 5944 19951 5946
rect 19812 5888 19890 5944
rect 19946 5888 19951 5944
rect 19812 5886 19951 5888
rect 19812 5884 19818 5886
rect 19885 5883 19951 5886
rect 3417 5810 3483 5813
rect 13077 5810 13143 5813
rect 18321 5810 18387 5813
rect 3417 5808 13002 5810
rect 3417 5752 3422 5808
rect 3478 5752 13002 5808
rect 3417 5750 13002 5752
rect 3417 5747 3483 5750
rect 0 5674 480 5704
rect 4981 5674 5047 5677
rect 0 5672 5047 5674
rect 0 5616 4986 5672
rect 5042 5616 5047 5672
rect 0 5614 5047 5616
rect 0 5584 480 5614
rect 4981 5611 5047 5614
rect 10358 5612 10364 5676
rect 10428 5674 10434 5676
rect 12433 5674 12499 5677
rect 10428 5672 12499 5674
rect 10428 5616 12438 5672
rect 12494 5616 12499 5672
rect 10428 5614 12499 5616
rect 12942 5674 13002 5750
rect 13077 5808 18387 5810
rect 13077 5752 13082 5808
rect 13138 5752 18326 5808
rect 18382 5752 18387 5808
rect 13077 5750 18387 5752
rect 13077 5747 13143 5750
rect 18321 5747 18387 5750
rect 15142 5674 15148 5676
rect 12942 5614 15148 5674
rect 10428 5612 10434 5614
rect 12433 5611 12499 5614
rect 15142 5612 15148 5614
rect 15212 5612 15218 5676
rect 15837 5674 15903 5677
rect 22320 5674 22800 5704
rect 15837 5672 22800 5674
rect 15837 5616 15842 5672
rect 15898 5616 22800 5672
rect 15837 5614 22800 5616
rect 15837 5611 15903 5614
rect 22320 5584 22800 5614
rect 1669 5538 1735 5541
rect 4889 5538 4955 5541
rect 5022 5538 5028 5540
rect 1669 5536 4170 5538
rect 1669 5480 1674 5536
rect 1730 5480 4170 5536
rect 1669 5478 4170 5480
rect 1669 5475 1735 5478
rect 0 5266 480 5296
rect 3550 5266 3556 5268
rect 0 5206 3556 5266
rect 0 5176 480 5206
rect 3550 5204 3556 5206
rect 3620 5266 3626 5268
rect 4110 5266 4170 5478
rect 4889 5536 5028 5538
rect 4889 5480 4894 5536
rect 4950 5480 5028 5536
rect 4889 5478 5028 5480
rect 4889 5475 4955 5478
rect 5022 5476 5028 5478
rect 5092 5476 5098 5540
rect 5441 5538 5507 5541
rect 8518 5538 8524 5540
rect 5441 5536 8524 5538
rect 5441 5480 5446 5536
rect 5502 5480 8524 5536
rect 5441 5478 8524 5480
rect 5441 5475 5507 5478
rect 8518 5476 8524 5478
rect 8588 5476 8594 5540
rect 13353 5538 13419 5541
rect 13997 5538 14063 5541
rect 13353 5536 14063 5538
rect 13353 5480 13358 5536
rect 13414 5480 14002 5536
rect 14058 5480 14063 5536
rect 13353 5478 14063 5480
rect 13353 5475 13419 5478
rect 13997 5475 14063 5478
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 5533 5402 5599 5405
rect 9397 5402 9463 5405
rect 13261 5404 13327 5405
rect 13261 5402 13308 5404
rect 5533 5400 9463 5402
rect 5533 5344 5538 5400
rect 5594 5344 9402 5400
rect 9458 5344 9463 5400
rect 5533 5342 9463 5344
rect 13216 5400 13308 5402
rect 13216 5344 13266 5400
rect 13216 5342 13308 5344
rect 5533 5339 5599 5342
rect 9397 5339 9463 5342
rect 13261 5340 13308 5342
rect 13372 5340 13378 5404
rect 13905 5402 13971 5405
rect 16573 5402 16639 5405
rect 13905 5400 16639 5402
rect 13905 5344 13910 5400
rect 13966 5344 16578 5400
rect 16634 5344 16639 5400
rect 13905 5342 16639 5344
rect 13261 5339 13327 5340
rect 13905 5339 13971 5342
rect 16573 5339 16639 5342
rect 5257 5266 5323 5269
rect 15469 5266 15535 5269
rect 3620 5206 4032 5266
rect 4110 5264 15535 5266
rect 4110 5208 5262 5264
rect 5318 5208 15474 5264
rect 15530 5208 15535 5264
rect 4110 5206 15535 5208
rect 3620 5204 3626 5206
rect 3972 5130 4032 5206
rect 5257 5203 5323 5206
rect 15469 5203 15535 5206
rect 15837 5266 15903 5269
rect 22320 5266 22800 5296
rect 15837 5264 22800 5266
rect 15837 5208 15842 5264
rect 15898 5208 22800 5264
rect 15837 5206 22800 5208
rect 15837 5203 15903 5206
rect 22320 5176 22800 5206
rect 7833 5130 7899 5133
rect 3972 5128 7899 5130
rect 3972 5072 7838 5128
rect 7894 5072 7899 5128
rect 3972 5070 7899 5072
rect 7833 5067 7899 5070
rect 9673 5130 9739 5133
rect 9857 5130 9923 5133
rect 9673 5128 9923 5130
rect 9673 5072 9678 5128
rect 9734 5072 9862 5128
rect 9918 5072 9923 5128
rect 9673 5070 9923 5072
rect 9673 5067 9739 5070
rect 9857 5067 9923 5070
rect 10961 5130 11027 5133
rect 11697 5130 11763 5133
rect 10961 5128 11763 5130
rect 10961 5072 10966 5128
rect 11022 5072 11702 5128
rect 11758 5072 11763 5128
rect 10961 5070 11763 5072
rect 10961 5067 11027 5070
rect 11697 5067 11763 5070
rect 13077 5130 13143 5133
rect 19149 5130 19215 5133
rect 13077 5128 19215 5130
rect 13077 5072 13082 5128
rect 13138 5072 19154 5128
rect 19210 5072 19215 5128
rect 13077 5070 19215 5072
rect 13077 5067 13143 5070
rect 19149 5067 19215 5070
rect 1669 4994 1735 4997
rect 4797 4994 4863 4997
rect 1669 4992 4863 4994
rect 1669 4936 1674 4992
rect 1730 4936 4802 4992
rect 4858 4936 4863 4992
rect 1669 4934 4863 4936
rect 1669 4931 1735 4934
rect 4797 4931 4863 4934
rect 4981 4994 5047 4997
rect 5574 4994 5580 4996
rect 4981 4992 5580 4994
rect 4981 4936 4986 4992
rect 5042 4936 5580 4992
rect 4981 4934 5580 4936
rect 4981 4931 5047 4934
rect 5574 4932 5580 4934
rect 5644 4932 5650 4996
rect 8845 4994 8911 4997
rect 10685 4994 10751 4997
rect 8845 4992 10751 4994
rect 8845 4936 8850 4992
rect 8906 4936 10690 4992
rect 10746 4936 10751 4992
rect 8845 4934 10751 4936
rect 8845 4931 8911 4934
rect 10685 4931 10751 4934
rect 11094 4932 11100 4996
rect 11164 4994 11170 4996
rect 12341 4994 12407 4997
rect 11164 4992 12407 4994
rect 11164 4936 12346 4992
rect 12402 4936 12407 4992
rect 11164 4934 12407 4936
rect 11164 4932 11170 4934
rect 12341 4931 12407 4934
rect 12617 4994 12683 4997
rect 14089 4994 14155 4997
rect 14406 4994 14412 4996
rect 12617 4992 13968 4994
rect 12617 4936 12622 4992
rect 12678 4936 13968 4992
rect 12617 4934 13968 4936
rect 12617 4931 12683 4934
rect 7808 4928 8128 4929
rect 0 4858 480 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 10174 4858 10180 4860
rect 0 4798 4906 4858
rect 0 4768 480 4798
rect 4846 4722 4906 4798
rect 9998 4798 10180 4858
rect 9998 4722 10058 4798
rect 10174 4796 10180 4798
rect 10244 4858 10250 4860
rect 13077 4858 13143 4861
rect 10244 4856 13143 4858
rect 10244 4800 13082 4856
rect 13138 4800 13143 4856
rect 10244 4798 13143 4800
rect 13908 4858 13968 4934
rect 14089 4992 14412 4994
rect 14089 4936 14094 4992
rect 14150 4936 14412 4992
rect 14089 4934 14412 4936
rect 14089 4931 14155 4934
rect 14406 4932 14412 4934
rect 14476 4932 14482 4996
rect 17493 4994 17559 4997
rect 19425 4994 19491 4997
rect 17493 4992 19491 4994
rect 17493 4936 17498 4992
rect 17554 4936 19430 4992
rect 19486 4936 19491 4992
rect 17493 4934 19491 4936
rect 17493 4931 17559 4934
rect 19425 4931 19491 4934
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 14089 4858 14155 4861
rect 13908 4856 14155 4858
rect 13908 4800 14094 4856
rect 14150 4800 14155 4856
rect 13908 4798 14155 4800
rect 10244 4796 10250 4798
rect 13077 4795 13143 4798
rect 14089 4795 14155 4798
rect 15101 4858 15167 4861
rect 22320 4858 22800 4888
rect 15101 4856 22800 4858
rect 15101 4800 15106 4856
rect 15162 4800 22800 4856
rect 15101 4798 22800 4800
rect 15101 4795 15167 4798
rect 22320 4768 22800 4798
rect 4846 4662 10058 4722
rect 10133 4722 10199 4725
rect 21817 4722 21883 4725
rect 10133 4720 21883 4722
rect 10133 4664 10138 4720
rect 10194 4664 21822 4720
rect 21878 4664 21883 4720
rect 10133 4662 21883 4664
rect 10133 4659 10199 4662
rect 21817 4659 21883 4662
rect 13261 4586 13327 4589
rect 4248 4584 13327 4586
rect 4248 4528 13266 4584
rect 13322 4528 13327 4584
rect 4248 4526 13327 4528
rect 0 4450 480 4480
rect 4248 4450 4308 4526
rect 13261 4523 13327 4526
rect 13486 4524 13492 4588
rect 13556 4586 13562 4588
rect 13556 4552 19258 4586
rect 13556 4526 19442 4552
rect 13556 4524 13562 4526
rect 19198 4492 19442 4526
rect 8569 4450 8635 4453
rect 0 4390 4308 4450
rect 7652 4448 8635 4450
rect 7652 4392 8574 4448
rect 8630 4392 8635 4448
rect 7652 4390 8635 4392
rect 0 4360 480 4390
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 5441 4314 5507 4317
rect 4846 4312 5507 4314
rect 4846 4256 5446 4312
rect 5502 4256 5507 4312
rect 4846 4254 5507 4256
rect 4337 4178 4403 4181
rect 4846 4178 4906 4254
rect 5441 4251 5507 4254
rect 5993 4314 6059 4317
rect 7652 4314 7712 4390
rect 8569 4387 8635 4390
rect 12801 4450 12867 4453
rect 13629 4450 13695 4453
rect 12801 4448 13695 4450
rect 12801 4392 12806 4448
rect 12862 4392 13634 4448
rect 13690 4392 13695 4448
rect 12801 4390 13695 4392
rect 19382 4450 19442 4492
rect 22320 4450 22800 4480
rect 19382 4390 22800 4450
rect 12801 4387 12867 4390
rect 13629 4387 13695 4390
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 22320 4360 22800 4390
rect 18104 4319 18424 4320
rect 14733 4314 14799 4317
rect 5993 4312 7712 4314
rect 5993 4256 5998 4312
rect 6054 4256 7712 4312
rect 5993 4254 7712 4256
rect 11654 4312 14799 4314
rect 11654 4256 14738 4312
rect 14794 4256 14799 4312
rect 11654 4254 14799 4256
rect 5993 4251 6059 4254
rect 4337 4176 4906 4178
rect 4337 4120 4342 4176
rect 4398 4120 4906 4176
rect 4337 4118 4906 4120
rect 4337 4115 4403 4118
rect 7230 4116 7236 4180
rect 7300 4178 7306 4180
rect 8845 4178 8911 4181
rect 11654 4178 11714 4254
rect 14733 4251 14799 4254
rect 7300 4176 11714 4178
rect 7300 4120 8850 4176
rect 8906 4120 11714 4176
rect 7300 4118 11714 4120
rect 7300 4116 7306 4118
rect 8845 4115 8911 4118
rect 12198 4116 12204 4180
rect 12268 4178 12274 4180
rect 13905 4178 13971 4181
rect 12268 4176 13971 4178
rect 12268 4120 13910 4176
rect 13966 4120 13971 4176
rect 12268 4118 13971 4120
rect 12268 4116 12274 4118
rect 13905 4115 13971 4118
rect 15469 4178 15535 4181
rect 16941 4178 17007 4181
rect 18045 4178 18111 4181
rect 18873 4178 18939 4181
rect 19241 4180 19307 4181
rect 19190 4178 19196 4180
rect 15469 4176 17188 4178
rect 15469 4120 15474 4176
rect 15530 4120 16946 4176
rect 17002 4120 17188 4176
rect 15469 4118 17188 4120
rect 15469 4115 15535 4118
rect 16941 4115 17007 4118
rect 0 4042 480 4072
rect 2998 4042 3004 4044
rect 0 3982 3004 4042
rect 0 3952 480 3982
rect 2998 3980 3004 3982
rect 3068 3980 3074 4044
rect 3693 4042 3759 4045
rect 5533 4042 5599 4045
rect 3693 4040 5599 4042
rect 3693 3984 3698 4040
rect 3754 3984 5538 4040
rect 5594 3984 5599 4040
rect 3693 3982 5599 3984
rect 3693 3979 3759 3982
rect 5533 3979 5599 3982
rect 5993 4042 6059 4045
rect 7414 4042 7420 4044
rect 5993 4040 7420 4042
rect 5993 3984 5998 4040
rect 6054 3984 7420 4040
rect 5993 3982 7420 3984
rect 5993 3979 6059 3982
rect 7414 3980 7420 3982
rect 7484 3980 7490 4044
rect 11094 4042 11100 4044
rect 7606 3982 11100 4042
rect 1117 3906 1183 3909
rect 3785 3906 3851 3909
rect 1117 3904 3851 3906
rect 1117 3848 1122 3904
rect 1178 3848 3790 3904
rect 3846 3848 3851 3904
rect 1117 3846 3851 3848
rect 1117 3843 1183 3846
rect 3785 3843 3851 3846
rect 5022 3844 5028 3908
rect 5092 3906 5098 3908
rect 7606 3906 7666 3982
rect 11094 3980 11100 3982
rect 11164 3980 11170 4044
rect 11973 4042 12039 4045
rect 12617 4042 12683 4045
rect 13813 4042 13879 4045
rect 15193 4042 15259 4045
rect 11973 4040 12683 4042
rect 11973 3984 11978 4040
rect 12034 3984 12622 4040
rect 12678 3984 12683 4040
rect 11973 3982 12683 3984
rect 11973 3979 12039 3982
rect 12617 3979 12683 3982
rect 12758 3982 13324 4042
rect 5092 3846 7666 3906
rect 5092 3844 5098 3846
rect 9438 3844 9444 3908
rect 9508 3906 9514 3908
rect 12758 3906 12818 3982
rect 9508 3846 12818 3906
rect 9508 3844 9514 3846
rect 12934 3844 12940 3908
rect 13004 3906 13010 3908
rect 13077 3906 13143 3909
rect 13004 3904 13143 3906
rect 13004 3848 13082 3904
rect 13138 3848 13143 3904
rect 13004 3846 13143 3848
rect 13264 3906 13324 3982
rect 13813 4040 15259 4042
rect 13813 3984 13818 4040
rect 13874 3984 15198 4040
rect 15254 3984 15259 4040
rect 13813 3982 15259 3984
rect 13813 3979 13879 3982
rect 15193 3979 15259 3982
rect 15653 4042 15719 4045
rect 16941 4042 17007 4045
rect 15653 4040 17007 4042
rect 15653 3984 15658 4040
rect 15714 3984 16946 4040
rect 17002 3984 17007 4040
rect 15653 3982 17007 3984
rect 17128 4042 17188 4118
rect 18045 4176 18939 4178
rect 18045 4120 18050 4176
rect 18106 4120 18878 4176
rect 18934 4120 18939 4176
rect 18045 4118 18939 4120
rect 19150 4118 19196 4178
rect 19260 4176 19307 4180
rect 19302 4120 19307 4176
rect 18045 4115 18111 4118
rect 18873 4115 18939 4118
rect 19190 4116 19196 4118
rect 19260 4116 19307 4120
rect 19241 4115 19307 4116
rect 19977 4178 20043 4181
rect 20897 4178 20963 4181
rect 19977 4176 20963 4178
rect 19977 4120 19982 4176
rect 20038 4120 20902 4176
rect 20958 4120 20963 4176
rect 19977 4118 20963 4120
rect 19977 4115 20043 4118
rect 20897 4115 20963 4118
rect 22320 4042 22800 4072
rect 17128 3982 22800 4042
rect 15653 3979 15719 3982
rect 16941 3979 17007 3982
rect 22320 3952 22800 3982
rect 14457 3906 14523 3909
rect 13264 3904 14523 3906
rect 13264 3848 14462 3904
rect 14518 3848 14523 3904
rect 13264 3846 14523 3848
rect 13004 3844 13010 3846
rect 13077 3843 13143 3846
rect 14457 3843 14523 3846
rect 15377 3906 15443 3909
rect 20478 3906 20484 3908
rect 15377 3904 20484 3906
rect 15377 3848 15382 3904
rect 15438 3848 20484 3904
rect 15377 3846 20484 3848
rect 15377 3843 15443 3846
rect 20478 3844 20484 3846
rect 20548 3844 20554 3908
rect 7808 3840 8128 3841
rect 0 3770 480 3800
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 2773 3770 2839 3773
rect 0 3768 2839 3770
rect 0 3712 2778 3768
rect 2834 3712 2839 3768
rect 0 3710 2839 3712
rect 0 3680 480 3710
rect 2773 3707 2839 3710
rect 5257 3770 5323 3773
rect 12801 3770 12867 3773
rect 13813 3770 13879 3773
rect 5257 3768 7712 3770
rect 5257 3712 5262 3768
rect 5318 3712 7712 3768
rect 5257 3710 7712 3712
rect 5257 3707 5323 3710
rect 933 3634 999 3637
rect 7373 3636 7439 3637
rect 7373 3634 7420 3636
rect 933 3632 7420 3634
rect 7484 3634 7490 3636
rect 7652 3634 7712 3710
rect 8204 3710 12266 3770
rect 8204 3634 8264 3710
rect 933 3576 938 3632
rect 994 3576 7378 3632
rect 933 3574 7420 3576
rect 933 3571 999 3574
rect 7373 3572 7420 3574
rect 7484 3574 7566 3634
rect 7652 3574 8264 3634
rect 7484 3572 7490 3574
rect 8518 3572 8524 3636
rect 8588 3634 8594 3636
rect 11973 3634 12039 3637
rect 8588 3632 12039 3634
rect 8588 3576 11978 3632
rect 12034 3576 12039 3632
rect 8588 3574 12039 3576
rect 12206 3634 12266 3710
rect 12801 3768 13879 3770
rect 12801 3712 12806 3768
rect 12862 3712 13818 3768
rect 13874 3712 13879 3768
rect 12801 3710 13879 3712
rect 12801 3707 12867 3710
rect 13813 3707 13879 3710
rect 15101 3770 15167 3773
rect 20345 3770 20411 3773
rect 15101 3768 20411 3770
rect 15101 3712 15106 3768
rect 15162 3712 20350 3768
rect 20406 3712 20411 3768
rect 15101 3710 20411 3712
rect 15101 3707 15167 3710
rect 20345 3707 20411 3710
rect 21173 3770 21239 3773
rect 22320 3770 22800 3800
rect 21173 3768 22800 3770
rect 21173 3712 21178 3768
rect 21234 3712 22800 3768
rect 21173 3710 22800 3712
rect 21173 3707 21239 3710
rect 22320 3680 22800 3710
rect 14825 3634 14891 3637
rect 12206 3632 14891 3634
rect 12206 3576 14830 3632
rect 14886 3576 14891 3632
rect 12206 3574 14891 3576
rect 8588 3572 8594 3574
rect 7373 3571 7439 3572
rect 11973 3571 12039 3574
rect 14825 3571 14891 3574
rect 15193 3634 15259 3637
rect 18781 3634 18847 3637
rect 20345 3634 20411 3637
rect 15193 3632 18568 3634
rect 15193 3576 15198 3632
rect 15254 3576 18568 3632
rect 15193 3574 18568 3576
rect 15193 3571 15259 3574
rect 3918 3436 3924 3500
rect 3988 3498 3994 3500
rect 4153 3498 4219 3501
rect 3988 3496 4219 3498
rect 3988 3440 4158 3496
rect 4214 3440 4219 3496
rect 3988 3438 4219 3440
rect 3988 3436 3994 3438
rect 4153 3435 4219 3438
rect 4337 3498 4403 3501
rect 5073 3500 5139 3501
rect 4337 3496 4860 3498
rect 4337 3440 4342 3496
rect 4398 3440 4860 3496
rect 4337 3438 4860 3440
rect 4337 3435 4403 3438
rect 0 3362 480 3392
rect 4245 3362 4311 3365
rect 0 3360 4311 3362
rect 0 3304 4250 3360
rect 4306 3304 4311 3360
rect 0 3302 4311 3304
rect 4800 3362 4860 3438
rect 5022 3436 5028 3500
rect 5092 3498 5139 3500
rect 6453 3498 6519 3501
rect 8477 3498 8543 3501
rect 10358 3498 10364 3500
rect 5092 3496 5184 3498
rect 5134 3440 5184 3496
rect 5092 3438 5184 3440
rect 6453 3496 10364 3498
rect 6453 3440 6458 3496
rect 6514 3440 8482 3496
rect 8538 3440 10364 3496
rect 6453 3438 10364 3440
rect 5092 3436 5139 3438
rect 5073 3435 5139 3436
rect 6453 3435 6519 3438
rect 8477 3435 8543 3438
rect 10358 3436 10364 3438
rect 10428 3436 10434 3500
rect 10961 3498 11027 3501
rect 12525 3498 12591 3501
rect 10961 3496 12591 3498
rect 10961 3440 10966 3496
rect 11022 3440 12530 3496
rect 12586 3440 12591 3496
rect 10961 3438 12591 3440
rect 10961 3435 11027 3438
rect 12525 3435 12591 3438
rect 7005 3362 7071 3365
rect 9121 3362 9187 3365
rect 4800 3302 6930 3362
rect 0 3272 480 3302
rect 4245 3299 4311 3302
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 3233 3226 3299 3229
rect 3877 3226 3943 3229
rect 5390 3226 5396 3228
rect 3233 3224 3943 3226
rect 3233 3168 3238 3224
rect 3294 3168 3882 3224
rect 3938 3168 3943 3224
rect 3233 3166 3943 3168
rect 3233 3163 3299 3166
rect 3877 3163 3943 3166
rect 5214 3166 5396 3226
rect 3785 3090 3851 3093
rect 5214 3090 5274 3166
rect 5390 3164 5396 3166
rect 5460 3164 5466 3228
rect 6870 3226 6930 3302
rect 7005 3360 9187 3362
rect 7005 3304 7010 3360
rect 7066 3304 9126 3360
rect 9182 3304 9187 3360
rect 7005 3302 9187 3304
rect 7005 3299 7071 3302
rect 9121 3299 9187 3302
rect 10685 3362 10751 3365
rect 11053 3362 11119 3365
rect 10685 3360 11119 3362
rect 10685 3304 10690 3360
rect 10746 3304 11058 3360
rect 11114 3304 11119 3360
rect 10685 3302 11119 3304
rect 10685 3299 10751 3302
rect 11053 3299 11119 3302
rect 11646 3300 11652 3364
rect 11716 3362 11722 3364
rect 18508 3362 18568 3574
rect 18781 3632 20411 3634
rect 18781 3576 18786 3632
rect 18842 3576 20350 3632
rect 20406 3576 20411 3632
rect 18781 3574 20411 3576
rect 18781 3571 18847 3574
rect 20345 3571 20411 3574
rect 20294 3362 20300 3364
rect 11716 3302 15946 3362
rect 18508 3302 20300 3362
rect 11716 3300 11722 3302
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 7465 3226 7531 3229
rect 6870 3224 7531 3226
rect 6870 3168 7470 3224
rect 7526 3168 7531 3224
rect 6870 3166 7531 3168
rect 7465 3163 7531 3166
rect 8293 3226 8359 3229
rect 9305 3226 9371 3229
rect 11789 3228 11855 3229
rect 11789 3226 11836 3228
rect 8293 3224 9371 3226
rect 8293 3168 8298 3224
rect 8354 3168 9310 3224
rect 9366 3168 9371 3224
rect 8293 3166 9371 3168
rect 11744 3224 11836 3226
rect 11744 3168 11794 3224
rect 11744 3166 11836 3168
rect 8293 3163 8359 3166
rect 9305 3163 9371 3166
rect 11789 3164 11836 3166
rect 11900 3164 11906 3228
rect 14457 3226 14523 3229
rect 15377 3226 15443 3229
rect 14457 3224 15443 3226
rect 14457 3168 14462 3224
rect 14518 3168 15382 3224
rect 15438 3168 15443 3224
rect 14457 3166 15443 3168
rect 11789 3163 11855 3164
rect 14457 3163 14523 3166
rect 15377 3163 15443 3166
rect 3785 3088 5274 3090
rect 3785 3032 3790 3088
rect 3846 3032 5274 3088
rect 3785 3030 5274 3032
rect 5349 3090 5415 3093
rect 8845 3090 8911 3093
rect 13261 3090 13327 3093
rect 5349 3088 8911 3090
rect 5349 3032 5354 3088
rect 5410 3032 8850 3088
rect 8906 3032 8911 3088
rect 5349 3030 8911 3032
rect 3785 3027 3851 3030
rect 5349 3027 5415 3030
rect 8845 3027 8911 3030
rect 9630 3088 13327 3090
rect 9630 3032 13266 3088
rect 13322 3032 13327 3088
rect 9630 3030 13327 3032
rect 0 2954 480 2984
rect 1117 2954 1183 2957
rect 0 2952 1183 2954
rect 0 2896 1122 2952
rect 1178 2896 1183 2952
rect 0 2894 1183 2896
rect 0 2864 480 2894
rect 1117 2891 1183 2894
rect 3693 2954 3759 2957
rect 9630 2954 9690 3030
rect 13261 3027 13327 3030
rect 14917 3090 14983 3093
rect 15326 3090 15332 3092
rect 14917 3088 15332 3090
rect 14917 3032 14922 3088
rect 14978 3032 15332 3088
rect 14917 3030 15332 3032
rect 14917 3027 14983 3030
rect 15326 3028 15332 3030
rect 15396 3028 15402 3092
rect 15886 3090 15946 3302
rect 20294 3300 20300 3302
rect 20364 3300 20370 3364
rect 20713 3362 20779 3365
rect 22320 3362 22800 3392
rect 20713 3360 22800 3362
rect 20713 3304 20718 3360
rect 20774 3304 22800 3360
rect 20713 3302 22800 3304
rect 20713 3299 20779 3302
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 22320 3272 22800 3302
rect 18104 3231 18424 3232
rect 15886 3030 19258 3090
rect 19198 2957 19258 3030
rect 3693 2952 9690 2954
rect 3693 2896 3698 2952
rect 3754 2896 9690 2952
rect 3693 2894 9690 2896
rect 10225 2954 10291 2957
rect 10910 2954 10916 2956
rect 10225 2952 10916 2954
rect 10225 2896 10230 2952
rect 10286 2896 10916 2952
rect 10225 2894 10916 2896
rect 3693 2891 3759 2894
rect 10225 2891 10291 2894
rect 10910 2892 10916 2894
rect 10980 2892 10986 2956
rect 11094 2892 11100 2956
rect 11164 2954 11170 2956
rect 14733 2954 14799 2957
rect 11164 2952 14799 2954
rect 11164 2896 14738 2952
rect 14794 2896 14799 2952
rect 11164 2894 14799 2896
rect 11164 2892 11170 2894
rect 14733 2891 14799 2894
rect 15377 2954 15443 2957
rect 19006 2954 19012 2956
rect 15377 2952 19012 2954
rect 15377 2896 15382 2952
rect 15438 2896 19012 2952
rect 15377 2894 19012 2896
rect 15377 2891 15443 2894
rect 19006 2892 19012 2894
rect 19076 2892 19082 2956
rect 19198 2952 19307 2957
rect 19198 2896 19246 2952
rect 19302 2896 19307 2952
rect 19198 2894 19307 2896
rect 19241 2891 19307 2894
rect 19425 2954 19491 2957
rect 21357 2954 21423 2957
rect 22320 2954 22800 2984
rect 19425 2952 22800 2954
rect 19425 2896 19430 2952
rect 19486 2896 21362 2952
rect 21418 2896 22800 2952
rect 19425 2894 22800 2896
rect 19425 2891 19491 2894
rect 21357 2891 21423 2894
rect 22320 2864 22800 2894
rect 1761 2818 1827 2821
rect 2681 2818 2747 2821
rect 1761 2816 2747 2818
rect 1761 2760 1766 2816
rect 1822 2760 2686 2816
rect 2742 2760 2747 2816
rect 1761 2758 2747 2760
rect 1761 2755 1827 2758
rect 2681 2755 2747 2758
rect 4245 2818 4311 2821
rect 9121 2820 9187 2821
rect 4838 2818 4844 2820
rect 4245 2816 4844 2818
rect 4245 2760 4250 2816
rect 4306 2760 4844 2816
rect 4245 2758 4844 2760
rect 4245 2755 4311 2758
rect 4838 2756 4844 2758
rect 4908 2756 4914 2820
rect 9070 2756 9076 2820
rect 9140 2818 9187 2820
rect 9765 2818 9831 2821
rect 11789 2818 11855 2821
rect 9140 2816 9232 2818
rect 9182 2760 9232 2816
rect 9140 2758 9232 2760
rect 9765 2816 11855 2818
rect 9765 2760 9770 2816
rect 9826 2760 11794 2816
rect 11850 2760 11855 2816
rect 9765 2758 11855 2760
rect 9140 2756 9187 2758
rect 9121 2755 9187 2756
rect 9765 2755 9831 2758
rect 11789 2755 11855 2758
rect 12985 2818 13051 2821
rect 13118 2818 13124 2820
rect 12985 2816 13124 2818
rect 12985 2760 12990 2816
rect 13046 2760 13124 2816
rect 12985 2758 13124 2760
rect 12985 2755 13051 2758
rect 13118 2756 13124 2758
rect 13188 2756 13194 2820
rect 21173 2818 21239 2821
rect 15104 2816 21239 2818
rect 15104 2760 21178 2816
rect 21234 2760 21239 2816
rect 15104 2758 21239 2760
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 2405 2682 2471 2685
rect 7097 2682 7163 2685
rect 10317 2684 10383 2685
rect 10317 2682 10364 2684
rect 2405 2680 7163 2682
rect 2405 2624 2410 2680
rect 2466 2624 7102 2680
rect 7158 2624 7163 2680
rect 2405 2622 7163 2624
rect 10272 2680 10364 2682
rect 10272 2624 10322 2680
rect 10272 2622 10364 2624
rect 2405 2619 2471 2622
rect 7097 2619 7163 2622
rect 10317 2620 10364 2622
rect 10428 2620 10434 2684
rect 14222 2682 14228 2684
rect 11884 2622 14228 2682
rect 10317 2619 10383 2620
rect 0 2546 480 2576
rect 1945 2546 2011 2549
rect 0 2544 2011 2546
rect 0 2488 1950 2544
rect 2006 2488 2011 2544
rect 0 2486 2011 2488
rect 0 2456 480 2486
rect 1945 2483 2011 2486
rect 4153 2546 4219 2549
rect 11884 2546 11944 2622
rect 14222 2620 14228 2622
rect 14292 2620 14298 2684
rect 4153 2544 11944 2546
rect 4153 2488 4158 2544
rect 4214 2488 11944 2544
rect 4153 2486 11944 2488
rect 13077 2546 13143 2549
rect 15104 2546 15164 2758
rect 21173 2755 21239 2758
rect 17125 2682 17191 2685
rect 17902 2682 17908 2684
rect 17125 2680 17908 2682
rect 17125 2624 17130 2680
rect 17186 2624 17908 2680
rect 17125 2622 17908 2624
rect 17125 2619 17191 2622
rect 17902 2620 17908 2622
rect 17972 2620 17978 2684
rect 20110 2682 20116 2684
rect 18278 2622 20116 2682
rect 13077 2544 15164 2546
rect 13077 2488 13082 2544
rect 13138 2488 15164 2544
rect 13077 2486 15164 2488
rect 16849 2546 16915 2549
rect 18278 2546 18338 2622
rect 20110 2620 20116 2622
rect 20180 2620 20186 2684
rect 16849 2544 18338 2546
rect 16849 2488 16854 2544
rect 16910 2488 18338 2544
rect 16849 2486 18338 2488
rect 4153 2483 4219 2486
rect 13077 2483 13143 2486
rect 16849 2483 16915 2486
rect 18822 2484 18828 2548
rect 18892 2546 18898 2548
rect 22320 2546 22800 2576
rect 18892 2486 22800 2546
rect 18892 2484 18898 2486
rect 22320 2456 22800 2486
rect 4337 2410 4403 2413
rect 14457 2410 14523 2413
rect 17166 2410 17172 2412
rect 4337 2408 12864 2410
rect 4337 2352 4342 2408
rect 4398 2352 12864 2408
rect 4337 2350 12864 2352
rect 4337 2347 4403 2350
rect 5574 2212 5580 2276
rect 5644 2274 5650 2276
rect 9121 2274 9187 2277
rect 5644 2272 9187 2274
rect 5644 2216 9126 2272
rect 9182 2216 9187 2272
rect 5644 2214 9187 2216
rect 12804 2274 12864 2350
rect 14457 2408 17172 2410
rect 14457 2352 14462 2408
rect 14518 2352 17172 2408
rect 14457 2350 17172 2352
rect 14457 2347 14523 2350
rect 17166 2348 17172 2350
rect 17236 2348 17242 2412
rect 17677 2410 17743 2413
rect 19558 2410 19564 2412
rect 17677 2408 19564 2410
rect 17677 2352 17682 2408
rect 17738 2352 19564 2408
rect 17677 2350 19564 2352
rect 17677 2347 17743 2350
rect 19558 2348 19564 2350
rect 19628 2348 19634 2412
rect 15377 2274 15443 2277
rect 12804 2272 15443 2274
rect 12804 2216 15382 2272
rect 15438 2216 15443 2272
rect 12804 2214 15443 2216
rect 5644 2212 5650 2214
rect 9121 2211 9187 2214
rect 15377 2211 15443 2214
rect 18597 2274 18663 2277
rect 20805 2274 20871 2277
rect 18597 2272 20871 2274
rect 18597 2216 18602 2272
rect 18658 2216 20810 2272
rect 20866 2216 20871 2272
rect 18597 2214 20871 2216
rect 18597 2211 18663 2214
rect 20805 2211 20871 2214
rect 4376 2208 4696 2209
rect 0 2138 480 2168
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 2957 2138 3023 2141
rect 0 2136 3023 2138
rect 0 2080 2962 2136
rect 3018 2080 3023 2136
rect 0 2078 3023 2080
rect 0 2048 480 2078
rect 2957 2075 3023 2078
rect 7373 2138 7439 2141
rect 8334 2138 8340 2140
rect 7373 2136 8340 2138
rect 7373 2080 7378 2136
rect 7434 2080 8340 2136
rect 7373 2078 8340 2080
rect 7373 2075 7439 2078
rect 8334 2076 8340 2078
rect 8404 2076 8410 2140
rect 19057 2138 19123 2141
rect 22320 2138 22800 2168
rect 19057 2136 22800 2138
rect 19057 2080 19062 2136
rect 19118 2080 22800 2136
rect 19057 2078 22800 2080
rect 19057 2075 19123 2078
rect 22320 2048 22800 2078
rect 6361 2002 6427 2005
rect 8518 2002 8524 2004
rect 6361 2000 8524 2002
rect 6361 1944 6366 2000
rect 6422 1944 8524 2000
rect 6361 1942 8524 1944
rect 6361 1939 6427 1942
rect 8518 1940 8524 1942
rect 8588 1940 8594 2004
rect 12014 1940 12020 2004
rect 12084 2002 12090 2004
rect 13629 2002 13695 2005
rect 12084 2000 13695 2002
rect 12084 1944 13634 2000
rect 13690 1944 13695 2000
rect 12084 1942 13695 1944
rect 12084 1940 12090 1942
rect 13629 1939 13695 1942
rect 16297 2002 16363 2005
rect 19374 2002 19380 2004
rect 16297 2000 19380 2002
rect 16297 1944 16302 2000
rect 16358 1944 19380 2000
rect 16297 1942 19380 1944
rect 16297 1939 16363 1942
rect 19374 1940 19380 1942
rect 19444 1940 19450 2004
rect 3693 1866 3759 1869
rect 17718 1866 17724 1868
rect 3693 1864 17724 1866
rect 3693 1808 3698 1864
rect 3754 1808 17724 1864
rect 3693 1806 17724 1808
rect 3693 1803 3759 1806
rect 17718 1804 17724 1806
rect 17788 1804 17794 1868
rect 0 1730 480 1760
rect 3049 1730 3115 1733
rect 0 1728 3115 1730
rect 0 1672 3054 1728
rect 3110 1672 3115 1728
rect 0 1670 3115 1672
rect 0 1640 480 1670
rect 3049 1667 3115 1670
rect 7281 1730 7347 1733
rect 8702 1730 8708 1732
rect 7281 1728 8708 1730
rect 7281 1672 7286 1728
rect 7342 1672 8708 1728
rect 7281 1670 8708 1672
rect 7281 1667 7347 1670
rect 8702 1668 8708 1670
rect 8772 1668 8778 1732
rect 17350 1668 17356 1732
rect 17420 1730 17426 1732
rect 18873 1730 18939 1733
rect 17420 1728 18939 1730
rect 17420 1672 18878 1728
rect 18934 1672 18939 1728
rect 17420 1670 18939 1672
rect 17420 1668 17426 1670
rect 18873 1667 18939 1670
rect 20805 1730 20871 1733
rect 22320 1730 22800 1760
rect 20805 1728 22800 1730
rect 20805 1672 20810 1728
rect 20866 1672 22800 1728
rect 20805 1670 22800 1672
rect 20805 1667 20871 1670
rect 22320 1640 22800 1670
rect 6177 1594 6243 1597
rect 6310 1594 6316 1596
rect 6177 1592 6316 1594
rect 6177 1536 6182 1592
rect 6238 1536 6316 1592
rect 6177 1534 6316 1536
rect 6177 1531 6243 1534
rect 6310 1532 6316 1534
rect 6380 1532 6386 1596
rect 8017 1594 8083 1597
rect 9438 1594 9444 1596
rect 8017 1592 9444 1594
rect 8017 1536 8022 1592
rect 8078 1536 9444 1592
rect 8017 1534 9444 1536
rect 8017 1531 8083 1534
rect 9438 1532 9444 1534
rect 9508 1532 9514 1596
rect 0 1322 480 1352
rect 4153 1322 4219 1325
rect 0 1320 4219 1322
rect 0 1264 4158 1320
rect 4214 1264 4219 1320
rect 0 1262 4219 1264
rect 0 1232 480 1262
rect 4153 1259 4219 1262
rect 18638 1260 18644 1324
rect 18708 1322 18714 1324
rect 19149 1322 19215 1325
rect 22320 1322 22800 1352
rect 18708 1320 22800 1322
rect 18708 1264 19154 1320
rect 19210 1264 22800 1320
rect 18708 1262 22800 1264
rect 18708 1260 18714 1262
rect 19149 1259 19215 1262
rect 22320 1232 22800 1262
rect 0 914 480 944
rect 3601 914 3667 917
rect 0 912 3667 914
rect 0 856 3606 912
rect 3662 856 3667 912
rect 0 854 3667 856
rect 0 824 480 854
rect 3601 851 3667 854
rect 21265 914 21331 917
rect 22320 914 22800 944
rect 21265 912 22800 914
rect 21265 856 21270 912
rect 21326 856 22800 912
rect 21265 854 22800 856
rect 21265 851 21331 854
rect 22320 824 22800 854
rect 0 506 480 536
rect 6085 506 6151 509
rect 0 504 6151 506
rect 0 448 6090 504
rect 6146 448 6151 504
rect 0 446 6151 448
rect 0 416 480 446
rect 6085 443 6151 446
rect 16481 506 16547 509
rect 22320 506 22800 536
rect 16481 504 22800 506
rect 16481 448 16486 504
rect 16542 448 22800 504
rect 16481 446 22800 448
rect 16481 443 16547 446
rect 22320 416 22800 446
rect 0 234 480 264
rect 3969 234 4035 237
rect 0 232 4035 234
rect 0 176 3974 232
rect 4030 176 4035 232
rect 0 174 4035 176
rect 0 144 480 174
rect 3969 171 4035 174
rect 19190 172 19196 236
rect 19260 234 19266 236
rect 22320 234 22800 264
rect 19260 174 22800 234
rect 19260 172 19266 174
rect 22320 144 22800 174
<< via3 >>
rect 7052 22204 7116 22268
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 14228 19408 14292 19412
rect 14228 19352 14242 19408
rect 14242 19352 14292 19408
rect 14228 19348 14292 19352
rect 12204 19076 12268 19140
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 11836 18940 11900 19004
rect 16436 18940 16500 19004
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 9628 18864 9692 18868
rect 9628 18808 9678 18864
rect 9678 18808 9692 18864
rect 9628 18804 9692 18808
rect 10548 18804 10612 18868
rect 8892 18668 8956 18732
rect 12756 18668 12820 18732
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 9628 18396 9692 18460
rect 13860 18396 13924 18460
rect 7052 17988 7116 18052
rect 8524 17988 8588 18052
rect 10364 17988 10428 18052
rect 15148 17988 15212 18052
rect 17356 17988 17420 18052
rect 17908 17988 17972 18052
rect 18644 17988 18708 18052
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 5764 17716 5828 17780
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 16252 17580 16316 17644
rect 12388 17444 12452 17508
rect 15700 17444 15764 17508
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 5212 17172 5276 17236
rect 11652 17036 11716 17100
rect 12020 17096 12084 17100
rect 12020 17040 12034 17096
rect 12034 17040 12084 17096
rect 12020 17036 12084 17040
rect 9076 16900 9140 16964
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 3556 16628 3620 16692
rect 4844 16492 4908 16556
rect 17724 16628 17788 16692
rect 19196 16688 19260 16692
rect 19196 16632 19246 16688
rect 19246 16632 19260 16688
rect 19196 16628 19260 16632
rect 19564 16688 19628 16692
rect 19564 16632 19578 16688
rect 19578 16632 19628 16688
rect 19564 16628 19628 16632
rect 20116 16688 20180 16692
rect 20116 16632 20130 16688
rect 20130 16632 20180 16688
rect 20116 16628 20180 16632
rect 10916 16356 10980 16420
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 12940 16084 13004 16148
rect 19748 16280 19812 16284
rect 19748 16224 19762 16280
rect 19762 16224 19812 16280
rect 19748 16220 19812 16224
rect 8340 15948 8404 16012
rect 16436 15948 16500 16012
rect 19012 15948 19076 16012
rect 15332 15812 15396 15876
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 12572 15676 12636 15740
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 16436 15540 16500 15604
rect 16988 15540 17052 15604
rect 6684 15464 6748 15468
rect 6684 15408 6698 15464
rect 6698 15408 6748 15464
rect 6684 15404 6748 15408
rect 13308 15404 13372 15468
rect 19380 15328 19444 15332
rect 19380 15272 19430 15328
rect 19430 15272 19444 15328
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 19380 15268 19444 15272
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 18828 15132 18892 15196
rect 17172 14724 17236 14788
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 15700 14588 15764 14652
rect 18828 14588 18892 14652
rect 8340 14452 8404 14516
rect 16620 14452 16684 14516
rect 17540 14452 17604 14516
rect 19748 14452 19812 14516
rect 9076 14316 9140 14380
rect 11100 14316 11164 14380
rect 16252 14180 16316 14244
rect 18828 14180 18892 14244
rect 19748 14180 19812 14244
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 9444 13772 9508 13836
rect 20300 13772 20364 13836
rect 20484 13832 20548 13836
rect 20484 13776 20534 13832
rect 20534 13776 20548 13832
rect 20484 13772 20548 13776
rect 6684 13696 6748 13700
rect 6684 13640 6734 13696
rect 6734 13640 6748 13696
rect 6684 13636 6748 13640
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 14412 13500 14476 13564
rect 16804 13500 16868 13564
rect 19748 13228 19812 13292
rect 15516 13092 15580 13156
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 10732 12956 10796 13020
rect 16620 12956 16684 13020
rect 17540 12880 17604 12884
rect 17540 12824 17590 12880
rect 17590 12824 17604 12880
rect 17540 12820 17604 12824
rect 5580 12684 5644 12748
rect 14044 12684 14108 12748
rect 15838 12684 15902 12748
rect 7236 12548 7300 12612
rect 11836 12608 11900 12612
rect 11836 12552 11886 12608
rect 11886 12552 11900 12608
rect 11836 12548 11900 12552
rect 16252 12548 16316 12612
rect 17540 12684 17604 12748
rect 18644 12684 18708 12748
rect 18644 12548 18708 12612
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 8708 12412 8772 12476
rect 9628 12472 9692 12476
rect 9628 12416 9642 12472
rect 9642 12416 9692 12472
rect 9628 12412 9692 12416
rect 9812 12412 9876 12476
rect 10180 12472 10244 12476
rect 10180 12416 10194 12472
rect 10194 12416 10244 12472
rect 10180 12412 10244 12416
rect 7236 12276 7300 12340
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 19748 12472 19812 12476
rect 19748 12416 19798 12472
rect 19798 12416 19812 12472
rect 19748 12412 19812 12416
rect 13124 12276 13188 12340
rect 10180 12140 10244 12204
rect 11836 12140 11900 12204
rect 8340 12004 8404 12068
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 5396 11928 5460 11932
rect 5396 11872 5410 11928
rect 5410 11872 5460 11928
rect 5396 11868 5460 11872
rect 15332 12004 15396 12068
rect 18828 12004 18892 12068
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 8340 11792 8404 11796
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 15700 11868 15764 11932
rect 16620 11868 16684 11932
rect 16988 11868 17052 11932
rect 8340 11736 8354 11792
rect 8354 11736 8404 11792
rect 8340 11732 8404 11736
rect 4844 11520 4908 11524
rect 4844 11464 4858 11520
rect 4858 11464 4908 11520
rect 4844 11460 4908 11464
rect 13124 11596 13188 11660
rect 10732 11460 10796 11524
rect 15332 11460 15396 11524
rect 16068 11520 16132 11524
rect 16068 11464 16118 11520
rect 16118 11464 16132 11520
rect 16068 11460 16132 11464
rect 16252 11460 16316 11524
rect 16804 11460 16868 11524
rect 19932 11460 19996 11524
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 9260 11324 9324 11388
rect 12756 11324 12820 11388
rect 13676 11324 13740 11388
rect 3004 11052 3068 11116
rect 5580 10976 5644 10980
rect 5580 10920 5594 10976
rect 5594 10920 5644 10976
rect 5580 10916 5644 10920
rect 12388 11052 12452 11116
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 10180 10840 10244 10844
rect 10180 10784 10194 10840
rect 10194 10784 10244 10840
rect 10180 10780 10244 10784
rect 12204 10780 12268 10844
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 18644 10780 18708 10844
rect 5212 10644 5276 10708
rect 5764 10644 5828 10708
rect 3556 10508 3620 10572
rect 17540 10644 17604 10708
rect 19748 10508 19812 10572
rect 8340 10432 8404 10436
rect 8340 10376 8390 10432
rect 8390 10376 8404 10432
rect 8340 10372 8404 10376
rect 8708 10432 8772 10436
rect 8708 10376 8722 10432
rect 8722 10376 8772 10432
rect 8708 10372 8772 10376
rect 9076 10432 9140 10436
rect 9076 10376 9090 10432
rect 9090 10376 9140 10432
rect 9076 10372 9140 10376
rect 9628 10372 9692 10436
rect 12204 10372 12268 10436
rect 12940 10372 13004 10436
rect 15516 10372 15580 10436
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4844 10296 4908 10300
rect 4844 10240 4894 10296
rect 4894 10240 4908 10296
rect 4844 10236 4908 10240
rect 7052 10296 7116 10300
rect 7052 10240 7066 10296
rect 7066 10240 7116 10296
rect 7052 10236 7116 10240
rect 16436 10100 16500 10164
rect 7236 9828 7300 9892
rect 9812 9828 9876 9892
rect 11100 9828 11164 9892
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 10180 9692 10244 9756
rect 7236 9556 7300 9620
rect 12020 9692 12084 9756
rect 18828 9828 18892 9892
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 13860 9556 13924 9620
rect 6316 9480 6380 9484
rect 6316 9424 6330 9480
rect 6330 9424 6380 9480
rect 6316 9420 6380 9424
rect 6868 9420 6932 9484
rect 10180 9420 10244 9484
rect 13492 9420 13556 9484
rect 3924 9284 3988 9348
rect 13676 9284 13740 9348
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 12204 9148 12268 9212
rect 5580 8876 5644 8940
rect 9076 8876 9140 8940
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 9444 8740 9508 8804
rect 11100 8740 11164 8804
rect 12940 8876 13004 8940
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 8892 8604 8956 8668
rect 12020 8392 12084 8396
rect 12020 8336 12034 8392
rect 12034 8336 12084 8392
rect 12020 8332 12084 8336
rect 16068 8332 16132 8396
rect 5396 8196 5460 8260
rect 8340 8196 8404 8260
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 8708 8060 8772 8124
rect 10548 7924 10612 7988
rect 18644 8256 18708 8260
rect 18644 8200 18694 8256
rect 18694 8200 18708 8256
rect 18644 8196 18708 8200
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 11836 7516 11900 7580
rect 14044 7576 14108 7580
rect 14412 7652 14476 7716
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 14044 7520 14094 7576
rect 14094 7520 14108 7576
rect 14044 7516 14108 7520
rect 7604 7380 7668 7444
rect 7052 7244 7116 7308
rect 7420 7244 7484 7308
rect 7236 7108 7300 7172
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 8524 7108 8588 7172
rect 16068 7244 16132 7308
rect 19196 7108 19260 7172
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 13124 6972 13188 7036
rect 18828 6972 18892 7036
rect 13124 6564 13188 6628
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 10364 6428 10428 6492
rect 6868 6020 6932 6084
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 11836 6020 11900 6084
rect 12572 6020 12636 6084
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 19748 5884 19812 5948
rect 10364 5612 10428 5676
rect 15148 5612 15212 5676
rect 3556 5204 3620 5268
rect 5028 5476 5092 5540
rect 8524 5476 8588 5540
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 13308 5400 13372 5404
rect 13308 5344 13322 5400
rect 13322 5344 13372 5400
rect 13308 5340 13372 5344
rect 5580 4932 5644 4996
rect 11100 4932 11164 4996
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 10180 4796 10244 4860
rect 14412 4932 14476 4996
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 13492 4524 13556 4588
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7236 4116 7300 4180
rect 12204 4116 12268 4180
rect 3004 3980 3068 4044
rect 7420 3980 7484 4044
rect 5028 3844 5092 3908
rect 11100 3980 11164 4044
rect 9444 3844 9508 3908
rect 12940 3844 13004 3908
rect 19196 4176 19260 4180
rect 19196 4120 19246 4176
rect 19246 4120 19260 4176
rect 19196 4116 19260 4120
rect 20484 3844 20548 3908
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 7420 3632 7484 3636
rect 7420 3576 7434 3632
rect 7434 3576 7484 3632
rect 7420 3572 7484 3576
rect 8524 3572 8588 3636
rect 3924 3436 3988 3500
rect 5028 3496 5092 3500
rect 5028 3440 5078 3496
rect 5078 3440 5092 3496
rect 5028 3436 5092 3440
rect 10364 3436 10428 3500
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 5396 3164 5460 3228
rect 11652 3300 11716 3364
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 11836 3224 11900 3228
rect 11836 3168 11850 3224
rect 11850 3168 11900 3224
rect 11836 3164 11900 3168
rect 15332 3028 15396 3092
rect 20300 3300 20364 3364
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 10916 2892 10980 2956
rect 11100 2892 11164 2956
rect 19012 2892 19076 2956
rect 4844 2756 4908 2820
rect 9076 2816 9140 2820
rect 9076 2760 9126 2816
rect 9126 2760 9140 2816
rect 9076 2756 9140 2760
rect 13124 2756 13188 2820
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 10364 2680 10428 2684
rect 10364 2624 10378 2680
rect 10378 2624 10428 2680
rect 10364 2620 10428 2624
rect 14228 2620 14292 2684
rect 17908 2620 17972 2684
rect 20116 2620 20180 2684
rect 18828 2484 18892 2548
rect 5580 2212 5644 2276
rect 17172 2348 17236 2412
rect 19564 2348 19628 2412
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
rect 8340 2076 8404 2140
rect 8524 1940 8588 2004
rect 12020 1940 12084 2004
rect 19380 1940 19444 2004
rect 17724 1804 17788 1868
rect 8708 1668 8772 1732
rect 17356 1668 17420 1732
rect 6316 1532 6380 1596
rect 9444 1532 9508 1596
rect 18644 1260 18708 1324
rect 19196 172 19260 236
<< metal4 >>
rect 7051 22268 7117 22269
rect 7051 22204 7052 22268
rect 7116 22204 7117 22268
rect 7051 22203 7117 22204
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 7054 18053 7114 22203
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7051 18052 7117 18053
rect 7051 17988 7052 18052
rect 7116 17988 7117 18052
rect 7051 17987 7117 17988
rect 7808 17984 8128 19008
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 9627 18868 9693 18869
rect 9627 18804 9628 18868
rect 9692 18804 9693 18868
rect 9627 18803 9693 18804
rect 10547 18868 10613 18869
rect 10547 18804 10548 18868
rect 10612 18804 10613 18868
rect 10547 18803 10613 18804
rect 8891 18732 8957 18733
rect 8891 18668 8892 18732
rect 8956 18668 8957 18732
rect 8891 18667 8957 18668
rect 8523 18052 8589 18053
rect 8523 17988 8524 18052
rect 8588 17988 8589 18052
rect 8523 17987 8589 17988
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 5763 17780 5829 17781
rect 5763 17716 5764 17780
rect 5828 17716 5829 17780
rect 5763 17715 5829 17716
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 3555 16692 3621 16693
rect 3555 16628 3556 16692
rect 3620 16628 3621 16692
rect 3555 16627 3621 16628
rect 3003 11116 3069 11117
rect 3003 11052 3004 11116
rect 3068 11052 3069 11116
rect 3003 11051 3069 11052
rect 3006 4045 3066 11051
rect 3558 10573 3618 16627
rect 4376 16352 4696 17376
rect 5211 17236 5277 17237
rect 5211 17172 5212 17236
rect 5276 17172 5277 17236
rect 5211 17171 5277 17172
rect 4843 16556 4909 16557
rect 4843 16492 4844 16556
rect 4908 16492 4909 16556
rect 4843 16491 4909 16492
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4846 11525 4906 16491
rect 4843 11524 4909 11525
rect 4843 11460 4844 11524
rect 4908 11460 4909 11524
rect 4843 11459 4909 11460
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 3555 10572 3621 10573
rect 3555 10508 3556 10572
rect 3620 10508 3621 10572
rect 3555 10507 3621 10508
rect 3558 5269 3618 10507
rect 4376 9824 4696 10848
rect 5214 10709 5274 17171
rect 5579 12748 5645 12749
rect 5579 12684 5580 12748
rect 5644 12684 5645 12748
rect 5579 12683 5645 12684
rect 5395 11932 5461 11933
rect 5395 11868 5396 11932
rect 5460 11868 5461 11932
rect 5395 11867 5461 11868
rect 5211 10708 5277 10709
rect 5211 10644 5212 10708
rect 5276 10644 5277 10708
rect 5211 10643 5277 10644
rect 4843 10300 4909 10301
rect 4843 10236 4844 10300
rect 4908 10236 4909 10300
rect 4843 10235 4909 10236
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 3923 9348 3989 9349
rect 3923 9284 3924 9348
rect 3988 9284 3989 9348
rect 3923 9283 3989 9284
rect 3555 5268 3621 5269
rect 3555 5204 3556 5268
rect 3620 5204 3621 5268
rect 3555 5203 3621 5204
rect 3003 4044 3069 4045
rect 3003 3980 3004 4044
rect 3068 3980 3069 4044
rect 3003 3979 3069 3980
rect 3926 3501 3986 9283
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 3923 3500 3989 3501
rect 3923 3436 3924 3500
rect 3988 3436 3989 3500
rect 3923 3435 3989 3436
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4846 2821 4906 10235
rect 5398 8261 5458 11867
rect 5582 10981 5642 12683
rect 5579 10980 5645 10981
rect 5579 10916 5580 10980
rect 5644 10916 5645 10980
rect 5579 10915 5645 10916
rect 5766 10709 5826 17715
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 8339 16012 8405 16013
rect 8339 15948 8340 16012
rect 8404 16010 8405 16012
rect 8526 16010 8586 17987
rect 8404 15950 8586 16010
rect 8404 15948 8405 15950
rect 8339 15947 8405 15948
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 6683 15468 6749 15469
rect 6683 15404 6684 15468
rect 6748 15404 6749 15468
rect 6683 15403 6749 15404
rect 6686 13701 6746 15403
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 6683 13700 6749 13701
rect 6683 13636 6684 13700
rect 6748 13636 6749 13700
rect 6683 13635 6749 13636
rect 7808 13632 8128 14656
rect 8339 14516 8405 14517
rect 8339 14452 8340 14516
rect 8404 14452 8405 14516
rect 8339 14451 8405 14452
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7235 12612 7301 12613
rect 7235 12548 7236 12612
rect 7300 12548 7301 12612
rect 7235 12547 7301 12548
rect 7238 12341 7298 12547
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7235 12340 7301 12341
rect 7235 12276 7236 12340
rect 7300 12276 7301 12340
rect 7235 12275 7301 12276
rect 7808 11456 8128 12480
rect 8342 12069 8402 14451
rect 8339 12068 8405 12069
rect 8339 12004 8340 12068
rect 8404 12004 8405 12068
rect 8339 12003 8405 12004
rect 8339 11796 8405 11797
rect 8339 11732 8340 11796
rect 8404 11732 8405 11796
rect 8339 11731 8405 11732
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 5763 10708 5829 10709
rect 5763 10644 5764 10708
rect 5828 10644 5829 10708
rect 5763 10643 5829 10644
rect 7808 10368 8128 11392
rect 8342 10437 8402 11731
rect 8339 10436 8405 10437
rect 8339 10372 8340 10436
rect 8404 10372 8405 10436
rect 8339 10371 8405 10372
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7051 10300 7117 10301
rect 7051 10236 7052 10300
rect 7116 10236 7117 10300
rect 7051 10235 7117 10236
rect 6315 9484 6381 9485
rect 6315 9420 6316 9484
rect 6380 9420 6381 9484
rect 6315 9419 6381 9420
rect 6867 9484 6933 9485
rect 6867 9420 6868 9484
rect 6932 9420 6933 9484
rect 6867 9419 6933 9420
rect 5579 8940 5645 8941
rect 5579 8876 5580 8940
rect 5644 8876 5645 8940
rect 5579 8875 5645 8876
rect 5395 8260 5461 8261
rect 5395 8196 5396 8260
rect 5460 8196 5461 8260
rect 5395 8195 5461 8196
rect 5027 5540 5093 5541
rect 5027 5476 5028 5540
rect 5092 5476 5093 5540
rect 5027 5475 5093 5476
rect 5030 3909 5090 5475
rect 5027 3908 5093 3909
rect 5027 3844 5028 3908
rect 5092 3844 5093 3908
rect 5027 3843 5093 3844
rect 5030 3501 5090 3843
rect 5027 3500 5093 3501
rect 5027 3436 5028 3500
rect 5092 3436 5093 3500
rect 5027 3435 5093 3436
rect 5398 3229 5458 8195
rect 5582 4997 5642 8875
rect 5579 4996 5645 4997
rect 5579 4932 5580 4996
rect 5644 4932 5645 4996
rect 5579 4931 5645 4932
rect 5395 3228 5461 3229
rect 5395 3164 5396 3228
rect 5460 3164 5461 3228
rect 5395 3163 5461 3164
rect 4843 2820 4909 2821
rect 4843 2756 4844 2820
rect 4908 2756 4909 2820
rect 4843 2755 4909 2756
rect 5582 2277 5642 4931
rect 5579 2276 5645 2277
rect 5579 2212 5580 2276
rect 5644 2212 5645 2276
rect 5579 2211 5645 2212
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 6318 1597 6378 9419
rect 6870 6085 6930 9419
rect 7054 7309 7114 10235
rect 7235 9892 7301 9893
rect 7235 9828 7236 9892
rect 7300 9828 7301 9892
rect 7235 9827 7301 9828
rect 7238 9621 7298 9827
rect 7235 9620 7301 9621
rect 7235 9556 7236 9620
rect 7300 9556 7301 9620
rect 7235 9555 7301 9556
rect 7051 7308 7117 7309
rect 7051 7244 7052 7308
rect 7116 7244 7117 7308
rect 7051 7243 7117 7244
rect 7238 7173 7298 9555
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 8339 8260 8405 8261
rect 8339 8196 8340 8260
rect 8404 8196 8405 8260
rect 8339 8195 8405 8196
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7603 7444 7669 7445
rect 7603 7380 7604 7444
rect 7668 7380 7669 7444
rect 7603 7379 7669 7380
rect 7419 7308 7485 7309
rect 7419 7244 7420 7308
rect 7484 7244 7485 7308
rect 7419 7243 7485 7244
rect 7235 7172 7301 7173
rect 7235 7108 7236 7172
rect 7300 7108 7301 7172
rect 7235 7107 7301 7108
rect 6867 6084 6933 6085
rect 6867 6020 6868 6084
rect 6932 6020 6933 6084
rect 6867 6019 6933 6020
rect 7238 4181 7298 7107
rect 7235 4180 7301 4181
rect 7235 4116 7236 4180
rect 7300 4116 7301 4180
rect 7235 4115 7301 4116
rect 7422 4045 7482 7243
rect 7419 4044 7485 4045
rect 7419 3980 7420 4044
rect 7484 3980 7485 4044
rect 7419 3979 7485 3980
rect 7606 3770 7666 7379
rect 7422 3710 7666 3770
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7422 3637 7482 3710
rect 7419 3636 7485 3637
rect 7419 3572 7420 3636
rect 7484 3572 7485 3636
rect 7419 3571 7485 3572
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 8342 2141 8402 8195
rect 8526 7173 8586 15950
rect 8707 12476 8773 12477
rect 8707 12412 8708 12476
rect 8772 12412 8773 12476
rect 8707 12411 8773 12412
rect 8710 10437 8770 12411
rect 8707 10436 8773 10437
rect 8707 10372 8708 10436
rect 8772 10372 8773 10436
rect 8707 10371 8773 10372
rect 8894 8669 8954 18667
rect 9630 18461 9690 18803
rect 9627 18460 9693 18461
rect 9627 18396 9628 18460
rect 9692 18396 9693 18460
rect 9627 18395 9693 18396
rect 10363 18052 10429 18053
rect 10363 17988 10364 18052
rect 10428 17988 10429 18052
rect 10363 17987 10429 17988
rect 9075 16964 9141 16965
rect 9075 16900 9076 16964
rect 9140 16900 9141 16964
rect 9075 16899 9141 16900
rect 9078 14381 9138 16899
rect 9075 14380 9141 14381
rect 9075 14316 9076 14380
rect 9140 14316 9141 14380
rect 9075 14315 9141 14316
rect 9078 10437 9138 14315
rect 9443 13836 9509 13837
rect 9443 13772 9444 13836
rect 9508 13772 9509 13836
rect 9443 13771 9509 13772
rect 9259 11388 9325 11389
rect 9259 11324 9260 11388
rect 9324 11324 9325 11388
rect 9259 11323 9325 11324
rect 9075 10436 9141 10437
rect 9075 10372 9076 10436
rect 9140 10372 9141 10436
rect 9075 10371 9141 10372
rect 9075 8940 9141 8941
rect 9075 8876 9076 8940
rect 9140 8876 9141 8940
rect 9075 8875 9141 8876
rect 8891 8668 8957 8669
rect 8891 8604 8892 8668
rect 8956 8604 8957 8668
rect 8891 8603 8957 8604
rect 8707 8124 8773 8125
rect 8707 8060 8708 8124
rect 8772 8060 8773 8124
rect 8707 8059 8773 8060
rect 8523 7172 8589 7173
rect 8523 7108 8524 7172
rect 8588 7108 8589 7172
rect 8523 7107 8589 7108
rect 8526 5541 8586 7107
rect 8523 5540 8589 5541
rect 8523 5476 8524 5540
rect 8588 5476 8589 5540
rect 8523 5475 8589 5476
rect 8523 3636 8589 3637
rect 8523 3572 8524 3636
rect 8588 3572 8589 3636
rect 8523 3571 8589 3572
rect 8339 2140 8405 2141
rect 8339 2076 8340 2140
rect 8404 2076 8405 2140
rect 8339 2075 8405 2076
rect 8526 2005 8586 3571
rect 8523 2004 8589 2005
rect 8523 1940 8524 2004
rect 8588 1940 8589 2004
rect 8523 1939 8589 1940
rect 8710 1733 8770 8059
rect 9078 2821 9138 8875
rect 9262 8666 9322 11323
rect 9446 8805 9506 13771
rect 9627 12476 9693 12477
rect 9627 12412 9628 12476
rect 9692 12412 9693 12476
rect 9627 12411 9693 12412
rect 9811 12476 9877 12477
rect 9811 12412 9812 12476
rect 9876 12412 9877 12476
rect 9811 12411 9877 12412
rect 10179 12476 10245 12477
rect 10179 12412 10180 12476
rect 10244 12412 10245 12476
rect 10179 12411 10245 12412
rect 9630 10437 9690 12411
rect 9627 10436 9693 10437
rect 9627 10372 9628 10436
rect 9692 10372 9693 10436
rect 9627 10371 9693 10372
rect 9814 9893 9874 12411
rect 10182 12205 10242 12411
rect 10179 12204 10245 12205
rect 10179 12140 10180 12204
rect 10244 12140 10245 12204
rect 10179 12139 10245 12140
rect 10179 10844 10245 10845
rect 10179 10780 10180 10844
rect 10244 10780 10245 10844
rect 10179 10779 10245 10780
rect 9811 9892 9877 9893
rect 9811 9828 9812 9892
rect 9876 9828 9877 9892
rect 9811 9827 9877 9828
rect 10182 9757 10242 10779
rect 10179 9756 10245 9757
rect 10179 9692 10180 9756
rect 10244 9692 10245 9756
rect 10179 9691 10245 9692
rect 10179 9484 10245 9485
rect 10179 9420 10180 9484
rect 10244 9420 10245 9484
rect 10179 9419 10245 9420
rect 9443 8804 9509 8805
rect 9443 8740 9444 8804
rect 9508 8740 9509 8804
rect 9443 8739 9509 8740
rect 9262 8606 9506 8666
rect 9446 3909 9506 8606
rect 10182 4861 10242 9419
rect 10366 6493 10426 17987
rect 10550 7989 10610 18803
rect 11240 18528 11560 19552
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14227 19412 14293 19413
rect 14227 19348 14228 19412
rect 14292 19348 14293 19412
rect 14227 19347 14293 19348
rect 12203 19140 12269 19141
rect 12203 19076 12204 19140
rect 12268 19076 12269 19140
rect 12203 19075 12269 19076
rect 11835 19004 11901 19005
rect 11835 18940 11836 19004
rect 11900 18940 11901 19004
rect 11835 18939 11901 18940
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 10915 16420 10981 16421
rect 10915 16356 10916 16420
rect 10980 16356 10981 16420
rect 10915 16355 10981 16356
rect 10731 13020 10797 13021
rect 10731 12956 10732 13020
rect 10796 12956 10797 13020
rect 10731 12955 10797 12956
rect 10734 11525 10794 12955
rect 10731 11524 10797 11525
rect 10731 11460 10732 11524
rect 10796 11460 10797 11524
rect 10731 11459 10797 11460
rect 10547 7988 10613 7989
rect 10547 7924 10548 7988
rect 10612 7924 10613 7988
rect 10547 7923 10613 7924
rect 10363 6492 10429 6493
rect 10363 6428 10364 6492
rect 10428 6428 10429 6492
rect 10363 6427 10429 6428
rect 10363 5676 10429 5677
rect 10363 5612 10364 5676
rect 10428 5612 10429 5676
rect 10363 5611 10429 5612
rect 10179 4860 10245 4861
rect 10179 4796 10180 4860
rect 10244 4796 10245 4860
rect 10179 4795 10245 4796
rect 9443 3908 9509 3909
rect 9443 3844 9444 3908
rect 9508 3844 9509 3908
rect 9443 3843 9509 3844
rect 9075 2820 9141 2821
rect 9075 2756 9076 2820
rect 9140 2756 9141 2820
rect 9075 2755 9141 2756
rect 8707 1732 8773 1733
rect 8707 1668 8708 1732
rect 8772 1668 8773 1732
rect 8707 1667 8773 1668
rect 9446 1597 9506 3843
rect 10366 3501 10426 5611
rect 10363 3500 10429 3501
rect 10363 3436 10364 3500
rect 10428 3436 10429 3500
rect 10363 3435 10429 3436
rect 10366 2685 10426 3435
rect 10918 2957 10978 16355
rect 11240 16352 11560 17376
rect 11651 17100 11717 17101
rect 11651 17036 11652 17100
rect 11716 17036 11717 17100
rect 11651 17035 11717 17036
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11099 14380 11165 14381
rect 11099 14316 11100 14380
rect 11164 14316 11165 14380
rect 11099 14315 11165 14316
rect 11102 9893 11162 14315
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11099 9892 11165 9893
rect 11099 9828 11100 9892
rect 11164 9828 11165 9892
rect 11099 9827 11165 9828
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11099 8804 11165 8805
rect 11099 8740 11100 8804
rect 11164 8740 11165 8804
rect 11099 8739 11165 8740
rect 11102 4997 11162 8739
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11099 4996 11165 4997
rect 11099 4932 11100 4996
rect 11164 4932 11165 4996
rect 11099 4931 11165 4932
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11099 4044 11165 4045
rect 11099 3980 11100 4044
rect 11164 3980 11165 4044
rect 11099 3979 11165 3980
rect 11102 2957 11162 3979
rect 11240 3296 11560 4320
rect 11654 3365 11714 17035
rect 11838 12613 11898 18939
rect 12019 17100 12085 17101
rect 12019 17036 12020 17100
rect 12084 17036 12085 17100
rect 12019 17035 12085 17036
rect 11835 12612 11901 12613
rect 11835 12548 11836 12612
rect 11900 12548 11901 12612
rect 11835 12547 11901 12548
rect 11835 12204 11901 12205
rect 11835 12140 11836 12204
rect 11900 12140 11901 12204
rect 11835 12139 11901 12140
rect 11838 7581 11898 12139
rect 12022 9757 12082 17035
rect 12206 10845 12266 19075
rect 12755 18732 12821 18733
rect 12755 18668 12756 18732
rect 12820 18668 12821 18732
rect 12755 18667 12821 18668
rect 12387 17508 12453 17509
rect 12387 17444 12388 17508
rect 12452 17444 12453 17508
rect 12387 17443 12453 17444
rect 12390 11117 12450 17443
rect 12571 15740 12637 15741
rect 12571 15676 12572 15740
rect 12636 15676 12637 15740
rect 12571 15675 12637 15676
rect 12387 11116 12453 11117
rect 12387 11052 12388 11116
rect 12452 11052 12453 11116
rect 12387 11051 12453 11052
rect 12203 10844 12269 10845
rect 12203 10780 12204 10844
rect 12268 10780 12269 10844
rect 12203 10779 12269 10780
rect 12203 10436 12269 10437
rect 12203 10372 12204 10436
rect 12268 10372 12269 10436
rect 12203 10371 12269 10372
rect 12019 9756 12085 9757
rect 12019 9692 12020 9756
rect 12084 9692 12085 9756
rect 12019 9691 12085 9692
rect 12206 9213 12266 10371
rect 12203 9212 12269 9213
rect 12203 9148 12204 9212
rect 12268 9148 12269 9212
rect 12203 9147 12269 9148
rect 12019 8396 12085 8397
rect 12019 8332 12020 8396
rect 12084 8332 12085 8396
rect 12019 8331 12085 8332
rect 11835 7580 11901 7581
rect 11835 7516 11836 7580
rect 11900 7516 11901 7580
rect 11835 7515 11901 7516
rect 11835 6084 11901 6085
rect 11835 6020 11836 6084
rect 11900 6020 11901 6084
rect 11835 6019 11901 6020
rect 11651 3364 11717 3365
rect 11651 3300 11652 3364
rect 11716 3300 11717 3364
rect 11651 3299 11717 3300
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 10915 2956 10981 2957
rect 10915 2892 10916 2956
rect 10980 2892 10981 2956
rect 10915 2891 10981 2892
rect 11099 2956 11165 2957
rect 11099 2892 11100 2956
rect 11164 2892 11165 2956
rect 11099 2891 11165 2892
rect 10363 2684 10429 2685
rect 10363 2620 10364 2684
rect 10428 2620 10429 2684
rect 10363 2619 10429 2620
rect 11240 2208 11560 3232
rect 11838 3229 11898 6019
rect 11835 3228 11901 3229
rect 11835 3164 11836 3228
rect 11900 3164 11901 3228
rect 11835 3163 11901 3164
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 12022 2005 12082 8331
rect 12206 4181 12266 9147
rect 12574 6085 12634 15675
rect 12758 11389 12818 18667
rect 13859 18460 13925 18461
rect 13859 18396 13860 18460
rect 13924 18396 13925 18460
rect 13859 18395 13925 18396
rect 12939 16148 13005 16149
rect 12939 16084 12940 16148
rect 13004 16084 13005 16148
rect 12939 16083 13005 16084
rect 12755 11388 12821 11389
rect 12755 11324 12756 11388
rect 12820 11324 12821 11388
rect 12755 11323 12821 11324
rect 12942 10437 13002 16083
rect 13307 15468 13373 15469
rect 13307 15404 13308 15468
rect 13372 15404 13373 15468
rect 13307 15403 13373 15404
rect 13123 12340 13189 12341
rect 13123 12276 13124 12340
rect 13188 12276 13189 12340
rect 13123 12275 13189 12276
rect 13126 11661 13186 12275
rect 13123 11660 13189 11661
rect 13123 11596 13124 11660
rect 13188 11596 13189 11660
rect 13123 11595 13189 11596
rect 12939 10436 13005 10437
rect 12939 10372 12940 10436
rect 13004 10372 13005 10436
rect 12939 10371 13005 10372
rect 12939 8940 13005 8941
rect 12939 8876 12940 8940
rect 13004 8876 13005 8940
rect 12939 8875 13005 8876
rect 12571 6084 12637 6085
rect 12571 6020 12572 6084
rect 12636 6020 12637 6084
rect 12571 6019 12637 6020
rect 12203 4180 12269 4181
rect 12203 4116 12204 4180
rect 12268 4116 12269 4180
rect 12203 4115 12269 4116
rect 12942 3909 13002 8875
rect 13123 7036 13189 7037
rect 13123 6972 13124 7036
rect 13188 6972 13189 7036
rect 13123 6971 13189 6972
rect 13126 6629 13186 6971
rect 13123 6628 13189 6629
rect 13123 6564 13124 6628
rect 13188 6564 13189 6628
rect 13123 6563 13189 6564
rect 12939 3908 13005 3909
rect 12939 3844 12940 3908
rect 13004 3844 13005 3908
rect 12939 3843 13005 3844
rect 13126 2821 13186 6563
rect 13310 5405 13370 15403
rect 13675 11388 13741 11389
rect 13675 11324 13676 11388
rect 13740 11324 13741 11388
rect 13675 11323 13741 11324
rect 13491 9484 13557 9485
rect 13491 9420 13492 9484
rect 13556 9420 13557 9484
rect 13491 9419 13557 9420
rect 13307 5404 13373 5405
rect 13307 5340 13308 5404
rect 13372 5340 13373 5404
rect 13307 5339 13373 5340
rect 13494 4589 13554 9419
rect 13678 9349 13738 11323
rect 13862 9621 13922 18395
rect 14043 12748 14109 12749
rect 14043 12684 14044 12748
rect 14108 12684 14109 12748
rect 14043 12683 14109 12684
rect 13859 9620 13925 9621
rect 13859 9556 13860 9620
rect 13924 9556 13925 9620
rect 13859 9555 13925 9556
rect 13675 9348 13741 9349
rect 13675 9284 13676 9348
rect 13740 9284 13741 9348
rect 13675 9283 13741 9284
rect 14046 7581 14106 12683
rect 14043 7580 14109 7581
rect 14043 7516 14044 7580
rect 14108 7516 14109 7580
rect 14043 7515 14109 7516
rect 13491 4588 13557 4589
rect 13491 4524 13492 4588
rect 13556 4524 13557 4588
rect 13491 4523 13557 4524
rect 13123 2820 13189 2821
rect 13123 2756 13124 2820
rect 13188 2756 13189 2820
rect 13123 2755 13189 2756
rect 14230 2685 14290 19347
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 16435 19004 16501 19005
rect 16435 18940 16436 19004
rect 16500 18940 16501 19004
rect 16435 18939 16501 18940
rect 15147 18052 15213 18053
rect 15147 17988 15148 18052
rect 15212 17988 15213 18052
rect 15147 17987 15213 17988
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14411 13564 14477 13565
rect 14411 13500 14412 13564
rect 14476 13500 14477 13564
rect 14411 13499 14477 13500
rect 14414 7717 14474 13499
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14411 7716 14477 7717
rect 14411 7652 14412 7716
rect 14476 7652 14477 7716
rect 14411 7651 14477 7652
rect 14414 4997 14474 7651
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14411 4996 14477 4997
rect 14411 4932 14412 4996
rect 14476 4932 14477 4996
rect 14411 4931 14477 4932
rect 14672 4928 14992 5952
rect 15150 5677 15210 17987
rect 16251 17644 16317 17645
rect 16251 17580 16252 17644
rect 16316 17580 16317 17644
rect 16251 17579 16317 17580
rect 15699 17508 15765 17509
rect 15699 17444 15700 17508
rect 15764 17444 15765 17508
rect 15699 17443 15765 17444
rect 15331 15876 15397 15877
rect 15331 15812 15332 15876
rect 15396 15812 15397 15876
rect 15331 15811 15397 15812
rect 15334 12069 15394 15811
rect 15702 14653 15762 17443
rect 15699 14652 15765 14653
rect 15699 14588 15700 14652
rect 15764 14588 15765 14652
rect 15699 14587 15765 14588
rect 15515 13156 15581 13157
rect 15515 13092 15516 13156
rect 15580 13092 15581 13156
rect 15515 13091 15581 13092
rect 15331 12068 15397 12069
rect 15331 12004 15332 12068
rect 15396 12004 15397 12068
rect 15331 12003 15397 12004
rect 15331 11524 15397 11525
rect 15331 11460 15332 11524
rect 15396 11460 15397 11524
rect 15331 11459 15397 11460
rect 15147 5676 15213 5677
rect 15147 5612 15148 5676
rect 15212 5612 15213 5676
rect 15147 5611 15213 5612
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 15334 3093 15394 11459
rect 15518 10437 15578 13091
rect 15702 11933 15762 14587
rect 16254 14245 16314 17579
rect 16438 16013 16498 18939
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 17355 18052 17421 18053
rect 17355 17988 17356 18052
rect 17420 17988 17421 18052
rect 17355 17987 17421 17988
rect 17907 18052 17973 18053
rect 17907 17988 17908 18052
rect 17972 17988 17973 18052
rect 17907 17987 17973 17988
rect 16435 16012 16501 16013
rect 16435 15948 16436 16012
rect 16500 15948 16501 16012
rect 16435 15947 16501 15948
rect 16435 15604 16501 15605
rect 16435 15540 16436 15604
rect 16500 15540 16501 15604
rect 16435 15539 16501 15540
rect 16987 15604 17053 15605
rect 16987 15540 16988 15604
rect 17052 15540 17053 15604
rect 16987 15539 17053 15540
rect 16251 14244 16317 14245
rect 16251 14180 16252 14244
rect 16316 14180 16317 14244
rect 16251 14179 16317 14180
rect 15837 12748 15903 12749
rect 15837 12684 15838 12748
rect 15902 12746 15903 12748
rect 15902 12684 15946 12746
rect 15837 12683 15946 12684
rect 15699 11932 15765 11933
rect 15699 11868 15700 11932
rect 15764 11868 15765 11932
rect 15699 11867 15765 11868
rect 15515 10436 15581 10437
rect 15515 10372 15516 10436
rect 15580 10372 15581 10436
rect 15515 10371 15581 10372
rect 15886 7306 15946 12683
rect 16251 12612 16317 12613
rect 16251 12548 16252 12612
rect 16316 12548 16317 12612
rect 16251 12547 16317 12548
rect 16254 11525 16314 12547
rect 16067 11524 16133 11525
rect 16067 11460 16068 11524
rect 16132 11460 16133 11524
rect 16067 11459 16133 11460
rect 16251 11524 16317 11525
rect 16251 11460 16252 11524
rect 16316 11460 16317 11524
rect 16251 11459 16317 11460
rect 16070 8397 16130 11459
rect 16438 10165 16498 15539
rect 16619 14516 16685 14517
rect 16619 14452 16620 14516
rect 16684 14452 16685 14516
rect 16619 14451 16685 14452
rect 16622 13021 16682 14451
rect 16803 13564 16869 13565
rect 16803 13500 16804 13564
rect 16868 13500 16869 13564
rect 16803 13499 16869 13500
rect 16619 13020 16685 13021
rect 16619 12956 16620 13020
rect 16684 12956 16685 13020
rect 16619 12955 16685 12956
rect 16622 11933 16682 12955
rect 16619 11932 16685 11933
rect 16619 11868 16620 11932
rect 16684 11868 16685 11932
rect 16619 11867 16685 11868
rect 16806 11525 16866 13499
rect 16990 11933 17050 15539
rect 17171 14788 17237 14789
rect 17171 14724 17172 14788
rect 17236 14724 17237 14788
rect 17171 14723 17237 14724
rect 16987 11932 17053 11933
rect 16987 11868 16988 11932
rect 17052 11868 17053 11932
rect 16987 11867 17053 11868
rect 16803 11524 16869 11525
rect 16803 11460 16804 11524
rect 16868 11460 16869 11524
rect 16803 11459 16869 11460
rect 16435 10164 16501 10165
rect 16435 10100 16436 10164
rect 16500 10100 16501 10164
rect 16435 10099 16501 10100
rect 16067 8396 16133 8397
rect 16067 8332 16068 8396
rect 16132 8332 16133 8396
rect 16067 8331 16133 8332
rect 16067 7308 16133 7309
rect 16067 7306 16068 7308
rect 15886 7246 16068 7306
rect 16067 7244 16068 7246
rect 16132 7244 16133 7308
rect 16067 7243 16133 7244
rect 15331 3092 15397 3093
rect 15331 3028 15332 3092
rect 15396 3028 15397 3092
rect 15331 3027 15397 3028
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14227 2684 14293 2685
rect 14227 2620 14228 2684
rect 14292 2620 14293 2684
rect 14227 2619 14293 2620
rect 14672 2128 14992 2688
rect 17174 2413 17234 14723
rect 17171 2412 17237 2413
rect 17171 2348 17172 2412
rect 17236 2348 17237 2412
rect 17171 2347 17237 2348
rect 12019 2004 12085 2005
rect 12019 1940 12020 2004
rect 12084 1940 12085 2004
rect 12019 1939 12085 1940
rect 17358 1733 17418 17987
rect 17723 16692 17789 16693
rect 17723 16628 17724 16692
rect 17788 16628 17789 16692
rect 17723 16627 17789 16628
rect 17539 14516 17605 14517
rect 17539 14452 17540 14516
rect 17604 14452 17605 14516
rect 17539 14451 17605 14452
rect 17542 12885 17602 14451
rect 17539 12884 17605 12885
rect 17539 12820 17540 12884
rect 17604 12820 17605 12884
rect 17539 12819 17605 12820
rect 17539 12748 17605 12749
rect 17539 12684 17540 12748
rect 17604 12684 17605 12748
rect 17539 12683 17605 12684
rect 17542 10709 17602 12683
rect 17539 10708 17605 10709
rect 17539 10644 17540 10708
rect 17604 10644 17605 10708
rect 17539 10643 17605 10644
rect 17726 1869 17786 16627
rect 17910 2685 17970 17987
rect 18104 17440 18424 18464
rect 18643 18052 18709 18053
rect 18643 17988 18644 18052
rect 18708 17988 18709 18052
rect 18643 17987 18709 17988
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18646 12749 18706 17987
rect 19195 16692 19261 16693
rect 19195 16628 19196 16692
rect 19260 16628 19261 16692
rect 19195 16627 19261 16628
rect 19563 16692 19629 16693
rect 19563 16628 19564 16692
rect 19628 16628 19629 16692
rect 19563 16627 19629 16628
rect 20115 16692 20181 16693
rect 20115 16628 20116 16692
rect 20180 16628 20181 16692
rect 20115 16627 20181 16628
rect 19011 16012 19077 16013
rect 19011 15948 19012 16012
rect 19076 15948 19077 16012
rect 19011 15947 19077 15948
rect 18827 15196 18893 15197
rect 18827 15132 18828 15196
rect 18892 15132 18893 15196
rect 18827 15131 18893 15132
rect 18830 14653 18890 15131
rect 18827 14652 18893 14653
rect 18827 14588 18828 14652
rect 18892 14588 18893 14652
rect 18827 14587 18893 14588
rect 18827 14244 18893 14245
rect 18827 14180 18828 14244
rect 18892 14180 18893 14244
rect 18827 14179 18893 14180
rect 18643 12748 18709 12749
rect 18643 12684 18644 12748
rect 18708 12684 18709 12748
rect 18643 12683 18709 12684
rect 18643 12612 18709 12613
rect 18643 12548 18644 12612
rect 18708 12548 18709 12612
rect 18643 12547 18709 12548
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18646 10845 18706 12547
rect 18830 12069 18890 14179
rect 18827 12068 18893 12069
rect 18827 12004 18828 12068
rect 18892 12004 18893 12068
rect 18827 12003 18893 12004
rect 18643 10844 18709 10845
rect 18643 10780 18644 10844
rect 18708 10780 18709 10844
rect 18643 10779 18709 10780
rect 18827 9892 18893 9893
rect 18827 9828 18828 9892
rect 18892 9828 18893 9892
rect 18827 9827 18893 9828
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18643 8260 18709 8261
rect 18643 8196 18644 8260
rect 18708 8196 18709 8260
rect 18643 8195 18709 8196
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 17907 2684 17973 2685
rect 17907 2620 17908 2684
rect 17972 2620 17973 2684
rect 17907 2619 17973 2620
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
rect 17723 1868 17789 1869
rect 17723 1804 17724 1868
rect 17788 1804 17789 1868
rect 17723 1803 17789 1804
rect 17355 1732 17421 1733
rect 17355 1668 17356 1732
rect 17420 1668 17421 1732
rect 17355 1667 17421 1668
rect 6315 1596 6381 1597
rect 6315 1532 6316 1596
rect 6380 1532 6381 1596
rect 6315 1531 6381 1532
rect 9443 1596 9509 1597
rect 9443 1532 9444 1596
rect 9508 1532 9509 1596
rect 9443 1531 9509 1532
rect 18646 1325 18706 8195
rect 18830 7037 18890 9827
rect 18827 7036 18893 7037
rect 18827 6972 18828 7036
rect 18892 6972 18893 7036
rect 18827 6971 18893 6972
rect 18830 2549 18890 6971
rect 19014 2957 19074 15947
rect 19198 7173 19258 16627
rect 19379 15332 19445 15333
rect 19379 15268 19380 15332
rect 19444 15268 19445 15332
rect 19379 15267 19445 15268
rect 19195 7172 19261 7173
rect 19195 7108 19196 7172
rect 19260 7108 19261 7172
rect 19195 7107 19261 7108
rect 19195 4180 19261 4181
rect 19195 4116 19196 4180
rect 19260 4116 19261 4180
rect 19195 4115 19261 4116
rect 19011 2956 19077 2957
rect 19011 2892 19012 2956
rect 19076 2892 19077 2956
rect 19011 2891 19077 2892
rect 18827 2548 18893 2549
rect 18827 2484 18828 2548
rect 18892 2484 18893 2548
rect 18827 2483 18893 2484
rect 18643 1324 18709 1325
rect 18643 1260 18644 1324
rect 18708 1260 18709 1324
rect 18643 1259 18709 1260
rect 19198 237 19258 4115
rect 19382 2005 19442 15267
rect 19566 2413 19626 16627
rect 19747 16284 19813 16285
rect 19747 16220 19748 16284
rect 19812 16220 19813 16284
rect 19747 16219 19813 16220
rect 19750 14517 19810 16219
rect 19747 14516 19813 14517
rect 19747 14452 19748 14516
rect 19812 14452 19813 14516
rect 19747 14451 19813 14452
rect 19747 14244 19813 14245
rect 19747 14180 19748 14244
rect 19812 14180 19813 14244
rect 19747 14179 19813 14180
rect 19750 13293 19810 14179
rect 19747 13292 19813 13293
rect 19747 13228 19748 13292
rect 19812 13228 19813 13292
rect 19747 13227 19813 13228
rect 19750 12610 19810 13227
rect 19750 12550 19994 12610
rect 19747 12476 19813 12477
rect 19747 12412 19748 12476
rect 19812 12412 19813 12476
rect 19747 12411 19813 12412
rect 19750 10573 19810 12411
rect 19934 11525 19994 12550
rect 19931 11524 19997 11525
rect 19931 11460 19932 11524
rect 19996 11460 19997 11524
rect 19931 11459 19997 11460
rect 19747 10572 19813 10573
rect 19747 10508 19748 10572
rect 19812 10508 19813 10572
rect 19747 10507 19813 10508
rect 19750 5949 19810 10507
rect 19747 5948 19813 5949
rect 19747 5884 19748 5948
rect 19812 5884 19813 5948
rect 19747 5883 19813 5884
rect 20118 2685 20178 16627
rect 20299 13836 20365 13837
rect 20299 13772 20300 13836
rect 20364 13772 20365 13836
rect 20299 13771 20365 13772
rect 20483 13836 20549 13837
rect 20483 13772 20484 13836
rect 20548 13772 20549 13836
rect 20483 13771 20549 13772
rect 20302 3365 20362 13771
rect 20486 3909 20546 13771
rect 20483 3908 20549 3909
rect 20483 3844 20484 3908
rect 20548 3844 20549 3908
rect 20483 3843 20549 3844
rect 20299 3364 20365 3365
rect 20299 3300 20300 3364
rect 20364 3300 20365 3364
rect 20299 3299 20365 3300
rect 20115 2684 20181 2685
rect 20115 2620 20116 2684
rect 20180 2620 20181 2684
rect 20115 2619 20181 2620
rect 19563 2412 19629 2413
rect 19563 2348 19564 2412
rect 19628 2348 19629 2412
rect 19563 2347 19629 2348
rect 19379 2004 19445 2005
rect 19379 1940 19380 2004
rect 19444 1940 19445 2004
rect 19379 1939 19445 1940
rect 19195 236 19261 237
rect 19195 172 19196 236
rect 19260 172 19261 236
rect 19195 171 19261 172
use sky130_fd_sc_hd__decap_3  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606256979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1606256979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1656 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1606256979
transform 1 0 1932 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18
timestamp 1606256979
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1606256979
transform 1 0 2668 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2944 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3496 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3864 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4416 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 3128 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1606256979
transform 1 0 4232 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32
timestamp 1606256979
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1606256979
transform 1 0 5336 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_2_
timestamp 1606256979
transform 1 0 5704 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_4_
timestamp 1606256979
transform 1 0 5888 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606256979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1606256979
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8464 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1606256979
transform 1 0 7912 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_4_
timestamp 1606256979
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1606256979
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_78
timestamp 1606256979
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _138_
timestamp 1606256979
transform 1 0 10120 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _145_
timestamp 1606256979
transform 1 0 9108 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 10672 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1606256979
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606256979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1606256979
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1606256979
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_96
timestamp 1606256979
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1606256979
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 11776 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1606256979
transform 1 0 10764 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606256979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1606256979
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1606256979
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1606256979
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 14076 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13432 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13616 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1606256979
transform 1 0 14352 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1606256979
transform 1 0 14352 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1606256979
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_142
timestamp 1606256979
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1606256979
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_140
timestamp 1606256979
transform 1 0 13984 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1606256979
transform 1 0 15640 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15824 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15180 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_3_
timestamp 1606256979
transform 1 0 16192 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606256979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1606256979
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156
timestamp 1606256979
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_162
timestamp 1606256979
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_159
timestamp 1606256979
transform 1 0 15732 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_176
timestamp 1606256979
transform 1 0 17296 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_173
timestamp 1606256979
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_2_
timestamp 1606256979
transform 1 0 17204 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_184
timestamp 1606256979
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1606256979
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1606256979
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606256979
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1606256979
transform 1 0 18216 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1606256979
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1606256979
transform 1 0 19504 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 19320 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_196
timestamp 1606256979
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_207
timestamp 1606256979
transform 1 0 20148 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1606256979
transform 1 0 19044 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_199
timestamp 1606256979
transform 1 0 19412 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_S_FTB01
timestamp 1606256979
transform 1 0 20516 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_S_FTB01
timestamp 1606256979
transform 1 0 20332 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606256979
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1606256979
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1606256979
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1606256979
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_217
timestamp 1606256979
transform 1 0 21068 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 2116 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1380 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1606256979
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1606256979
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4416 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1606256979
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_32
timestamp 1606256979
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_5_
timestamp 1606256979
transform 1 0 6624 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5428 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1606256979
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_56
timestamp 1606256979
transform 1 0 6256 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1606256979
transform 1 0 7636 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_69
timestamp 1606256979
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1606256979
transform 1 0 8464 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 8832 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1606256979
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_102
timestamp 1606256979
transform 1 0 10488 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 10764 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1606256979
transform 1 0 12420 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_121
timestamp 1606256979
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1606256979
transform 1 0 13432 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_132
timestamp 1606256979
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_143
timestamp 1606256979
transform 1 0 14260 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_S_FTB01
timestamp 1606256979
transform 1 0 16376 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1606256979
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1606256979
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1606256979
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_165
timestamp 1606256979
transform 1 0 16284 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 17112 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_172
timestamp 1606256979
transform 1 0 16928 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 18768 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1606256979
transform 1 0 19780 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_190
timestamp 1606256979
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_201
timestamp 1606256979
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_212
timestamp 1606256979
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1606256979
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1606256979
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 2668 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 1656 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1606256979
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1606256979
transform 1 0 4508 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_4_
timestamp 1606256979
transform 1 0 3680 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_26
timestamp 1606256979
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_41
timestamp 1606256979
transform 1 0 4876 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1606256979
transform 1 0 6164 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l5_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1606256979
transform 1 0 4968 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1606256979
transform 1 0 5796 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606256979
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1606256979
transform 1 0 8096 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8648 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_71
timestamp 1606256979
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_75
timestamp 1606256979
transform 1 0 8004 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_80
timestamp 1606256979
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 10304 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_98
timestamp 1606256979
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1606256979
transform 1 0 12512 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1606256979
transform 1 0 11224 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_106
timestamp 1606256979
transform 1 0 10856 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1606256979
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1606256979
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13064 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_128
timestamp 1606256979
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 14720 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15732 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1606256979
transform 1 0 16284 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_146
timestamp 1606256979
transform 1 0 14536 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_157
timestamp 1606256979
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1606256979
transform 1 0 17480 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 18032 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1606256979
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_174
timestamp 1606256979
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1606256979
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1606256979
transform 1 0 19688 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1606256979
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1606256979
transform 1 0 20700 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_211
timestamp 1606256979
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp 1606256979
transform 1 0 21068 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 1472 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_5_
timestamp 1606256979
transform 1 0 2944 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1606256979
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1606256979
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1606256979
transform 1 0 4600 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1606256979
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_36
timestamp 1606256979
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 5704 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_4_47
timestamp 1606256979
transform 1 0 5428 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8372 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 7360 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1606256979
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_77
timestamp 1606256979
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _148_
timestamp 1606256979
transform 1 0 9936 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10488 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1606256979
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_93
timestamp 1606256979
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_100
timestamp 1606256979
transform 1 0 10304 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12512 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 11500 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_111
timestamp 1606256979
transform 1 0 11316 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_122
timestamp 1606256979
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13524 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_133
timestamp 1606256979
transform 1 0 13340 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_144
timestamp 1606256979
transform 1 0 14352 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1606256979
transform 1 0 14628 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_4_
timestamp 1606256979
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16376 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1606256979
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_163
timestamp 1606256979
transform 1 0 16100 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 17388 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_175
timestamp 1606256979
transform 1 0 17204 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_186
timestamp 1606256979
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1606256979
transform 1 0 20148 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_2_S_FTB01
timestamp 1606256979
transform 1 0 18400 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1606256979
transform 1 0 19136 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1606256979
transform 1 0 18952 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_205
timestamp 1606256979
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1606256979
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_211
timestamp 1606256979
transform 1 0 20516 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_218
timestamp 1606256979
transform 1 0 21160 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1606256979
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 1932 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_7
timestamp 1606256979
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1606256979
transform 1 0 4600 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1606256979
transform 1 0 3588 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_25
timestamp 1606256979
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_36
timestamp 1606256979
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606256979
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_1_
timestamp 1606256979
transform 1 0 5704 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_47
timestamp 1606256979
transform 1 0 5428 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606256979
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8740 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1606256979
transform 1 0 8280 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_82
timestamp 1606256979
transform 1 0 8648 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1606256979
transform 1 0 10396 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_99
timestamp 1606256979
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1606256979
transform 1 0 10948 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_4_
timestamp 1606256979
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_105
timestamp 1606256979
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_116
timestamp 1606256979
transform 1 0 11776 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13708 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1606256979
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_134
timestamp 1606256979
transform 1 0 13432 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 15824 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_4_
timestamp 1606256979
transform 1 0 14812 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_5_146
timestamp 1606256979
transform 1 0 14536 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_158
timestamp 1606256979
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1606256979
transform 1 0 17480 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1606256979
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_176
timestamp 1606256979
transform 1 0 17296 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1606256979
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 18860 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_188
timestamp 1606256979
transform 1 0 18400 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_192
timestamp 1606256979
transform 1 0 18768 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 20516 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_209
timestamp 1606256979
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_217
timestamp 1606256979
transform 1 0 21068 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1606256979
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1606256979
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1564 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1606256979
transform 1 0 1932 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1606256979
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_18
timestamp 1606256979
transform 1 0 2760 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1606256979
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1606256979
transform 1 0 2852 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 2300 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4048 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_3_
timestamp 1606256979
transform 1 0 4048 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1606256979
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1606256979
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_28
timestamp 1606256979
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_41
timestamp 1606256979
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1606256979
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1606256979
transform 1 0 5704 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1606256979
transform 1 0 6164 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1606256979
transform 1 0 5888 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5060 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_48
timestamp 1606256979
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_53
timestamp 1606256979
transform 1 0 5980 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 7820 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_6_
timestamp 1606256979
transform 1 0 8188 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_7_
timestamp 1606256979
transform 1 0 7176 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1606256979
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_64
timestamp 1606256979
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_75
timestamp 1606256979
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_65
timestamp 1606256979
transform 1 0 7084 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_82
timestamp 1606256979
transform 1 0 8648 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1606256979
transform 1 0 9200 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9752 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_86
timestamp 1606256979
transform 1 0 9016 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1606256979
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_110
timestamp 1606256979
transform 1 0 11224 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1606256979
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1606256979
transform 1 0 11316 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1606256979
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1606256979
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_120
timestamp 1606256979
transform 1 0 12144 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _141_
timestamp 1606256979
transform 1 0 12512 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1606256979
transform 1 0 11776 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 12604 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1606256979
transform 1 0 14444 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13064 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_128
timestamp 1606256979
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_141
timestamp 1606256979
transform 1 0 14076 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1606256979
transform 1 0 14720 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 14996 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1606256979
transform 1 0 15456 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_146
timestamp 1606256979
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1606256979
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1606256979
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_165
timestamp 1606256979
transform 1 0 16284 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_149
timestamp 1606256979
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 16744 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1606256979
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1606256979
transform 1 0 16928 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_169
timestamp 1606256979
transform 1 0 16652 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_186
timestamp 1606256979
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_167
timestamp 1606256979
transform 1 0 16468 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_171
timestamp 1606256979
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1606256979
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 19320 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 19412 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1606256979
transform 1 0 18400 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1606256979
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_208
timestamp 1606256979
transform 1 0 20240 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_193
timestamp 1606256979
transform 1 0 18860 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_197
timestamp 1606256979
transform 1 0 19228 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606256979
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606256979
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_214
timestamp 1606256979
transform 1 0 20792 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1606256979
transform 1 0 1564 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1606256979
transform 1 0 2116 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1606256979
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_9
timestamp 1606256979
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_20
timestamp 1606256979
transform 1 0 2944 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1606256979
transform 1 0 3404 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1606256979
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_24
timestamp 1606256979
transform 1 0 3312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1606256979
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_41
timestamp 1606256979
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_3_
timestamp 1606256979
transform 1 0 5060 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6256 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1606256979
transform 1 0 6072 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_52
timestamp 1606256979
transform 1 0 5888 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_3_
timestamp 1606256979
transform 1 0 8556 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 7544 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 7268 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_65
timestamp 1606256979
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_79
timestamp 1606256979
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9844 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1606256979
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1606256979
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_104
timestamp 1606256979
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10856 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1606256979
transform 1 0 11868 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_115
timestamp 1606256979
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12880 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 14168 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1606256979
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_126
timestamp 1606256979
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1606256979
transform 1 0 13708 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1606256979
transform 1 0 16284 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1606256979
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1606256979
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1606256979
transform 1 0 17848 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 16836 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_169
timestamp 1606256979
transform 1 0 16652 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_180
timestamp 1606256979
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 19136 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_191
timestamp 1606256979
transform 1 0 18676 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1606256979
transform 1 0 19044 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1606256979
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1606256979
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_218
timestamp 1606256979
transform 1 0 21160 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1748 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 3772 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_9_23
timestamp 1606256979
transform 1 0 3220 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1606256979
transform 1 0 5428 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_45
timestamp 1606256979
transform 1 0 5244 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_56
timestamp 1606256979
transform 1 0 6256 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1606256979
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_62
timestamp 1606256979
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7084 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_9_81
timestamp 1606256979
transform 1 0 8556 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1606256979
transform 1 0 8832 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1606256979
transform 1 0 9844 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_93
timestamp 1606256979
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_104
timestamp 1606256979
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1606256979
transform 1 0 11868 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12420 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10856 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_115
timestamp 1606256979
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1606256979
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_4_
timestamp 1606256979
transform 1 0 14076 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_139
timestamp 1606256979
transform 1 0 13892 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1606256979
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 15364 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 15088 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_150
timestamp 1606256979
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_164
timestamp 1606256979
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1606256979
transform 1 0 17388 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1606256979
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1606256979
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1606256979
transform 1 0 20056 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1606256979
transform 1 0 19044 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1606256979
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_204
timestamp 1606256979
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_215
timestamp 1606256979
transform 1 0 20884 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1606256979
transform 1 0 21252 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 2300 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1564 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1606256979
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1606256979
transform 1 0 2116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1606256979
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1606256979
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1606256979
transform 1 0 6348 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 5060 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 6072 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_52
timestamp 1606256979
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_61
timestamp 1606256979
transform 1 0 6716 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7912 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6900 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_72
timestamp 1606256979
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1606256979
transform 1 0 9936 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10580 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1606256979
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_93
timestamp 1606256979
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_100
timestamp 1606256979
transform 1 0 10304 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1606256979
transform 1 0 12236 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_119
timestamp 1606256979
transform 1 0 12052 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13524 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 13248 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_130
timestamp 1606256979
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1606256979
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1606256979
transform 1 0 16100 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1606256979
transform 1 0 16468 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 17020 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_171
timestamp 1606256979
transform 1 0 16836 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1606256979
transform 1 0 19688 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1606256979
transform 1 0 18676 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_189
timestamp 1606256979
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_200
timestamp 1606256979
transform 1 0 19504 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_211
timestamp 1606256979
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1606256979
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1606256979
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1606256979
transform 1 0 1380 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_5_
timestamp 1606256979
transform 1 0 2392 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_12
timestamp 1606256979
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _146_
timestamp 1606256979
transform 1 0 3404 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4048 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_23
timestamp 1606256979
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_29
timestamp 1606256979
transform 1 0 3772 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_48
timestamp 1606256979
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606256979
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1606256979
transform 1 0 8464 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_78
timestamp 1606256979
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10488 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9476 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_89
timestamp 1606256979
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_100
timestamp 1606256979
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1606256979
transform 1 0 11776 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_111
timestamp 1606256979
transform 1 0 11316 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_115
timestamp 1606256979
transform 1 0 11684 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1606256979
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1606256979
transform 1 0 13432 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1606256979
transform 1 0 14444 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_132
timestamp 1606256979
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_143
timestamp 1606256979
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1606256979
transform 1 0 15548 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16100 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_11_154
timestamp 1606256979
transform 1 0 15272 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_161
timestamp 1606256979
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1606256979
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1606256979
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1606256979
transform 1 0 20056 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1606256979
transform 1 0 19044 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1606256979
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_204
timestamp 1606256979
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_215
timestamp 1606256979
transform 1 0 20884 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_219
timestamp 1606256979
transform 1 0 21252 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1606256979
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_7_
timestamp 1606256979
transform 1 0 2944 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_1_
timestamp 1606256979
transform 1 0 1932 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1606256979
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_18
timestamp 1606256979
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_4_
timestamp 1606256979
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1606256979
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1606256979
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5060 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6716 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1606256979
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 7820 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_12_70
timestamp 1606256979
transform 1 0 7544 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1606256979
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_89
timestamp 1606256979
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_102
timestamp 1606256979
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 10856 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l4_in_0_
timestamp 1606256979
transform 1 0 12512 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_122
timestamp 1606256979
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1606256979
transform 1 0 13524 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1606256979
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_144
timestamp 1606256979
transform 1 0 14352 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _143_
timestamp 1606256979
transform 1 0 14628 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1606256979
transform 1 0 16284 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_4_
timestamp 1606256979
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1606256979
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1606256979
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 18216 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 17480 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_174
timestamp 1606256979
transform 1 0 17112 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_184
timestamp 1606256979
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19872 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_202
timestamp 1606256979
transform 1 0 19688 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1606256979
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606256979
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1606256979
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_8
timestamp 1606256979
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1606256979
transform 1 0 1380 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_9
timestamp 1606256979
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1606256979
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1606256979
transform 1 0 1564 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1606256979
transform 1 0 1472 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_19
timestamp 1606256979
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_3_
timestamp 1606256979
transform 1 0 2024 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_2_
timestamp 1606256979
transform 1 0 2116 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_20
timestamp 1606256979
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1606256979
transform 1 0 3036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4048 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1606256979
transform 1 0 4876 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_6_
timestamp 1606256979
transform 1 0 3128 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4048 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_31
timestamp 1606256979
transform 1 0 3956 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_25
timestamp 1606256979
transform 1 0 3404 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1606256979
transform 1 0 6808 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5980 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 5704 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606256979
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_48
timestamp 1606256979
transform 1 0 5520 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_52
timestamp 1606256979
transform 1 0 5888 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1606256979
transform 1 0 8004 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8740 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7084 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1606256979
transform 1 0 8556 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 7728 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1606256979
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_71
timestamp 1606256979
transform 1 0 7636 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_79
timestamp 1606256979
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1606256979
transform 1 0 10396 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_3_
timestamp 1606256979
transform 1 0 10672 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1606256979
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1606256979
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1606256979
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1606256979
transform 1 0 11776 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _147_
timestamp 1606256979
transform 1 0 11868 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1606256979
transform 1 0 12420 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_110
timestamp 1606256979
transform 1 0 11224 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1606256979
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_113
timestamp 1606256979
transform 1 0 11500 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_121
timestamp 1606256979
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 14352 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1606256979
transform 1 0 13432 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 14076 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_139
timestamp 1606256979
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_132
timestamp 1606256979
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_143
timestamp 1606256979
transform 1 0 14260 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1606256979
transform 1 0 15364 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1606256979
transform 1 0 14628 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 15824 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_153
timestamp 1606256979
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_158
timestamp 1606256979
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1606256979
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_173
timestamp 1606256979
transform 1 0 17020 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_176
timestamp 1606256979
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1606256979
transform 1 0 17204 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1606256979
transform 1 0 16744 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_186
timestamp 1606256979
transform 1 0 18216 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1606256979
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_3_
timestamp 1606256979
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1606256979
transform 1 0 17388 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1606256979
transform 1 0 17480 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1606256979
transform 1 0 18492 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606256979
transform 1 0 19044 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1606256979
transform 1 0 20056 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19044 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_193
timestamp 1606256979
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_204
timestamp 1606256979
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_193
timestamp 1606256979
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606256979
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1606256979
transform 1 0 20884 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_219
timestamp 1606256979
transform 1 0 21252 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1606256979
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606256979
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1606256979
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1606256979
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 1840 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_6
timestamp 1606256979
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1606256979
transform 1 0 3496 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1606256979
transform 1 0 3956 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1606256979
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_30
timestamp 1606256979
transform 1 0 3864 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_40
timestamp 1606256979
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1606256979
transform 1 0 6164 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1606256979
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606256979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1606256979
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1606256979
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1606256979
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_62 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6808 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1606256979
transform 1 0 7820 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1606256979
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_70
timestamp 1606256979
transform 1 0 7544 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_82
timestamp 1606256979
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9752 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_1_
timestamp 1606256979
transform 1 0 8832 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_93
timestamp 1606256979
transform 1 0 9660 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1606256979
transform 1 0 11868 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _144_
timestamp 1606256979
transform 1 0 11500 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606256979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_110
timestamp 1606256979
transform 1 0 11224 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1606256979
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1606256979
transform 1 0 13432 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1606256979
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_143
timestamp 1606256979
transform 1 0 14260 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_3_
timestamp 1606256979
transform 1 0 15824 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1606256979
transform 1 0 14812 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_158
timestamp 1606256979
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18032 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1606256979
transform 1 0 16928 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606256979
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_169
timestamp 1606256979
transform 1 0 16652 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1606256979
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_2_
timestamp 1606256979
transform 1 0 19872 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1606256979
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1606256979
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_213
timestamp 1606256979
transform 1 0 20700 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_219
timestamp 1606256979
transform 1 0 21252 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1606256979
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606256979
transform 1 0 1840 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_6
timestamp 1606256979
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1606256979
transform 1 0 3496 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606256979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_24
timestamp 1606256979
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1606256979
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 1606256979
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1606256979
transform 1 0 5060 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 5704 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_47
timestamp 1606256979
transform 1 0 5428 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7360 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_66
timestamp 1606256979
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _126_
timestamp 1606256979
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _149_
timestamp 1606256979
transform 1 0 9660 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606256979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 10396 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_16_84
timestamp 1606256979
transform 1 0 8832 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_97
timestamp 1606256979
transform 1 0 10028 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12420 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_121
timestamp 1606256979
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_1_
timestamp 1606256979
transform 1 0 14076 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_139
timestamp 1606256979
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1606256979
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606256979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1606256979
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1606256979
transform 1 0 16100 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1606256979
transform 1 0 16560 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1606256979
transform 1 0 17572 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_167
timestamp 1606256979
transform 1 0 16468 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_177
timestamp 1606256979
transform 1 0 17388 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1606256979
transform 1 0 18584 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 19136 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_188
timestamp 1606256979
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1606256979
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606256979
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1606256979
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606256979
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606256979
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l5_in_0_
timestamp 1606256979
transform 1 0 2116 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_9
timestamp 1606256979
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_20
timestamp 1606256979
transform 1 0 2944 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1606256979
transform 1 0 4876 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 3220 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_39
timestamp 1606256979
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1606256979
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1606256979
transform 1 0 5520 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606256979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_45
timestamp 1606256979
transform 1 0 5244 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1606256979
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1606256979
transform 1 0 7820 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_71
timestamp 1606256979
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_82
timestamp 1606256979
transform 1 0 8648 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10672 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9844 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_2_
timestamp 1606256979
transform 1 0 9016 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l4_in_0_
timestamp 1606256979
transform 1 0 11500 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606256979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 14352 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 14076 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1606256979
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1606256979
transform 1 0 16376 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 16008 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_160
timestamp 1606256979
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_165
timestamp 1606256979
transform 1 0 16284 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 18032 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16928 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606256979
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_170
timestamp 1606256979
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1606256979
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l4_in_0_
timestamp 1606256979
transform 1 0 19688 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1606256979
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1606256979
transform 1 0 20700 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_211
timestamp 1606256979
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_217
timestamp 1606256979
transform 1 0 21068 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1606256979
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1606256979
transform 1 0 2944 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1606256979
transform 1 0 1932 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_7
timestamp 1606256979
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_18
timestamp 1606256979
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1606256979
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4692 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606256979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1606256979
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_36
timestamp 1606256979
transform 1 0 4416 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6348 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_55
timestamp 1606256979
transform 1 0 6164 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8372 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l4_in_0_
timestamp 1606256979
transform 1 0 7360 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_66
timestamp 1606256979
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_77
timestamp 1606256979
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 9752 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606256979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1606256979
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1606256979
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 11408 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_110
timestamp 1606256979
transform 1 0 11224 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1606256979
transform 1 0 13064 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_3_
timestamp 1606256979
transform 1 0 14076 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_128
timestamp 1606256979
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_139
timestamp 1606256979
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15456 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606256979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_150
timestamp 1606256979
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1606256979
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_165
timestamp 1606256979
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16468 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 18216 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_183
timestamp 1606256979
transform 1 0 17940 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19872 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_202
timestamp 1606256979
transform 1 0 19688 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1606256979
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606256979
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1606256979
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_218
timestamp 1606256979
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1606256979
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1606256979
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1564 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1606256979
transform 1 0 1564 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1606256979
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_14
timestamp 1606256979
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 2300 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 2576 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1606256979
transform 1 0 4232 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4140 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606256979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_32
timestamp 1606256979
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1606256979
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_32
timestamp 1606256979
transform 1 0 4048 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_42
timestamp 1606256979
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_43
timestamp 1606256979
transform 1 0 5060 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1606256979
transform 1 0 5152 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5428 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_59
timestamp 1606256979
transform 1 0 6532 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_53
timestamp 1606256979
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_56
timestamp 1606256979
transform 1 0 6256 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606256979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1606256979
transform 1 0 6164 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1606256979
transform 1 0 6808 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1606256979
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7268 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7820 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1606256979
transform 1 0 7084 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_83
timestamp 1606256979
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_71
timestamp 1606256979
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1606256979
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1606256979
transform 1 0 10672 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _142_
timestamp 1606256979
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9936 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1606256979
transform 1 0 8924 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1606256979
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606256979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_94
timestamp 1606256979
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1606256979
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1606256979
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_108
timestamp 1606256979
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_105
timestamp 1606256979
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1606256979
transform 1 0 10948 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1606256979
transform 1 0 11224 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_123
timestamp 1606256979
transform 1 0 12420 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_119
timestamp 1606256979
transform 1 0 12052 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_123
timestamp 1606256979
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1606256979
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_116
timestamp 1606256979
transform 1 0 11776 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606256979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1606256979
transform 1 0 11868 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12512 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13524 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12696 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1606256979
transform 1 0 14352 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_142
timestamp 1606256979
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_133
timestamp 1606256979
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1606256979
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_153
timestamp 1606256979
transform 1 0 15180 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 15272 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606256979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_163
timestamp 1606256979
transform 1 0 16100 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_161
timestamp 1606256979
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1606256979
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1606256979
transform 1 0 16284 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1606256979
transform 1 0 15548 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1606256979
transform 1 0 16376 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1606256979
transform 1 0 17388 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_1_
timestamp 1606256979
transform 1 0 17388 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18124 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606256979
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_174
timestamp 1606256979
transform 1 0 17112 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1606256979
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_184
timestamp 1606256979
transform 1 0 18032 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_175
timestamp 1606256979
transform 1 0 17204 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_186
timestamp 1606256979
transform 1 0 18216 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_1_
timestamp 1606256979
transform 1 0 19412 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_2_
timestamp 1606256979
transform 1 0 18400 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_3_
timestamp 1606256979
transform 1 0 18860 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_1_
timestamp 1606256979
transform 1 0 19872 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_191
timestamp 1606256979
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_202
timestamp 1606256979
transform 1 0 19688 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1606256979
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_208
timestamp 1606256979
transform 1 0 20240 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606256979
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_213
timestamp 1606256979
transform 1 0 20700 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_219
timestamp 1606256979
transform 1 0 21252 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606256979
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606256979
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1606256979
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_1_
timestamp 1606256979
transform 1 0 2852 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 1840 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_6
timestamp 1606256979
transform 1 0 1656 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_17
timestamp 1606256979
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 3864 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_28
timestamp 1606256979
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1606256979
transform 1 0 5704 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 6808 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606256979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_46
timestamp 1606256979
transform 1 0 5336 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1606256979
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7728 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_68
timestamp 1606256979
transform 1 0 7360 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _140_
timestamp 1606256979
transform 1 0 9384 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1606256979
transform 1 0 9936 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_88
timestamp 1606256979
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_94
timestamp 1606256979
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1606256979
transform 1 0 10948 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606256979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1606256979
transform 1 0 10764 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_116
timestamp 1606256979
transform 1 0 11776 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_123
timestamp 1606256979
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 12788 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_21_143
timestamp 1606256979
transform 1 0 14260 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1606256979
transform 1 0 14536 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15088 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_150
timestamp 1606256979
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18032 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16744 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606256979
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_168
timestamp 1606256979
transform 1 0 16560 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1606256979
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1606256979
transform 1 0 19688 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1606256979
transform 1 0 19504 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1606256979
transform 1 0 20700 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_211
timestamp 1606256979
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_217
timestamp 1606256979
transform 1 0 21068 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1606256979
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_3_
timestamp 1606256979
transform 1 0 1840 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2852 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_6
timestamp 1606256979
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_17
timestamp 1606256979
transform 1 0 2668 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4232 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606256979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_28
timestamp 1606256979
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1606256979
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1606256979
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5888 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_43
timestamp 1606256979
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_49
timestamp 1606256979
transform 1 0 5612 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1606256979
transform 1 0 7544 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8556 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_68
timestamp 1606256979
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_79
timestamp 1606256979
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _139_
timestamp 1606256979
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10304 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606256979
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1606256979
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_97
timestamp 1606256979
transform 1 0 10028 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1606256979
transform 1 0 11316 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1606256979
transform 1 0 12328 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_109
timestamp 1606256979
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_120
timestamp 1606256979
transform 1 0 12144 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14444 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1606256979
transform 1 0 13340 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_131
timestamp 1606256979
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_142
timestamp 1606256979
transform 1 0 14168 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1606256979
transform 1 0 16008 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15272 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606256979
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1606256979
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_160
timestamp 1606256979
transform 1 0 15824 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 17020 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_171
timestamp 1606256979
transform 1 0 16836 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_3_
timestamp 1606256979
transform 1 0 19688 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_2_
timestamp 1606256979
transform 1 0 18492 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1606256979
transform 1 0 19504 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_198
timestamp 1606256979
transform 1 0 19320 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1606256979
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606256979
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_211
timestamp 1606256979
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_218
timestamp 1606256979
transform 1 0 21160 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1656 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606256979
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1606256979
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 3312 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_22
timestamp 1606256979
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_40
timestamp 1606256979
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4968 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1606256979
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606256979
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_58
timestamp 1606256979
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1606256979
transform 1 0 7820 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 8648 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 8372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1606256979
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_77
timestamp 1606256979
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 10304 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_98
timestamp 1606256979
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606256979
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_116
timestamp 1606256979
transform 1 0 11776 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1606256979
transform 1 0 13524 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 14076 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_23_132
timestamp 1606256979
transform 1 0 13248 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_139
timestamp 1606256979
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1606256979
transform 1 0 15732 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 16192 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_157
timestamp 1606256979
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_162
timestamp 1606256979
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606256979
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1606256979
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_184
timestamp 1606256979
transform 1 0 18032 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_2_
timestamp 1606256979
transform 1 0 19044 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1606256979
transform 1 0 20056 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606256979
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_192
timestamp 1606256979
transform 1 0 18768 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_204
timestamp 1606256979
transform 1 0 19872 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606256979
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1606256979
transform 1 0 20884 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1606256979
transform 1 0 21252 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1606256979
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_2_
timestamp 1606256979
transform 1 0 2944 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_3_
timestamp 1606256979
transform 1 0 1932 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606256979
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1606256979
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_18
timestamp 1606256979
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1606256979
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1606256979
transform 1 0 4508 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606256979
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1606256979
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_35
timestamp 1606256979
transform 1 0 4324 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1606256979
transform 1 0 5520 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 6532 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_46
timestamp 1606256979
transform 1 0 5336 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_57
timestamp 1606256979
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_62
timestamp 1606256979
transform 1 0 6808 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 6900 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1606256979
transform 1 0 8556 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_79
timestamp 1606256979
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1606256979
transform 1 0 10672 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_4_
timestamp 1606256979
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606256979
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1606256979
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_102
timestamp 1606256979
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11132 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_107
timestamp 1606256979
transform 1 0 10948 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_125
timestamp 1606256979
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  clk_3_E_FTB01
timestamp 1606256979
transform 1 0 14444 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12788 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_143
timestamp 1606256979
transform 1 0 14260 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1606256979
transform 1 0 16376 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_2_
timestamp 1606256979
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606256979
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1606256979
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1606256979
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_165
timestamp 1606256979
transform 1 0 16284 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_3_
timestamp 1606256979
transform 1 0 17388 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l4_in_0_
timestamp 1606256979
transform 1 0 18216 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_175
timestamp 1606256979
transform 1 0 17204 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1606256979
transform 1 0 19412 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_195
timestamp 1606256979
transform 1 0 19044 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_208
timestamp 1606256979
transform 1 0 20240 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606256979
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606256979
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606256979
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606256979
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1606256979
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1840 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1606256979
transform 1 0 2576 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606256979
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1606256979
transform 1 0 1748 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_14
timestamp 1606256979
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1606256979
transform 1 0 4784 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_3_
timestamp 1606256979
transform 1 0 3772 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_25
timestamp 1606256979
transform 1 0 3404 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_38
timestamp 1606256979
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1606256979
transform 1 0 6256 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 6808 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5244 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606256979
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_43
timestamp 1606256979
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1606256979
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1606256979
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _137_
timestamp 1606256979
transform 1 0 8648 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_78
timestamp 1606256979
transform 1 0 8280 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10396 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1606256979
transform 1 0 9384 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1606256979
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_86
timestamp 1606256979
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_99
timestamp 1606256979
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606256979
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_117
timestamp 1606256979
transform 1 0 11868 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1606256979
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_3_
timestamp 1606256979
transform 1 0 13432 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1606256979
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_143
timestamp 1606256979
transform 1 0 14260 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1606256979
transform 1 0 15824 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_3_
timestamp 1606256979
transform 1 0 14812 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_158
timestamp 1606256979
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_1_
timestamp 1606256979
transform 1 0 16836 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18216 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606256979
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1606256979
transform 1 0 16652 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1606256979
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_184
timestamp 1606256979
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_1_
timestamp 1606256979
transform 1 0 19044 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l5_in_0_
timestamp 1606256979
transform 1 0 20056 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_204
timestamp 1606256979
transform 1 0 19872 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606256979
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1606256979
transform 1 0 20884 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1606256979
transform 1 0 21252 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_9
timestamp 1606256979
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1606256979
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1606256979
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606256979
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606256979
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_5_
timestamp 1606256979
transform 1 0 1932 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1380 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_18
timestamp 1606256979
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_6_
timestamp 1606256979
transform 1 0 2944 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 2116 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_7_
timestamp 1606256979
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_2_
timestamp 1606256979
transform 1 0 4048 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606256979
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1606256979
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1606256979
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1606256979
transform 1 0 3588 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_31
timestamp 1606256979
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_41
timestamp 1606256979
transform 1 0 4876 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_43
timestamp 1606256979
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1606256979
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_4_
timestamp 1606256979
transform 1 0 5244 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1606256979
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1606256979
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_61
timestamp 1606256979
transform 1 0 6716 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606256979
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1606256979
transform 1 0 6256 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5244 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _136_
timestamp 1606256979
transform 1 0 7820 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7912 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 6900 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8372 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_72
timestamp 1606256979
transform 1 0 7728 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_71
timestamp 1606256979
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_77
timestamp 1606256979
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_88
timestamp 1606256979
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_93
timestamp 1606256979
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1606256979
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606256979
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1606256979
transform 1 0 9384 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_99
timestamp 1606256979
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_100
timestamp 1606256979
transform 1 0 10304 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1606256979
transform 1 0 10396 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _134_
timestamp 1606256979
transform 1 0 9936 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10488 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _130_
timestamp 1606256979
transform 1 0 11776 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1606256979
transform 1 0 12236 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606256979
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_118
timestamp 1606256979
transform 1 0 11960 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_110
timestamp 1606256979
transform 1 0 11224 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1606256979
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13708 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12972 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_26_127
timestamp 1606256979
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_145
timestamp 1606256979
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_132
timestamp 1606256979
transform 1 0 13248 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_136
timestamp 1606256979
transform 1 0 13616 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1606256979
transform 1 0 14628 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 15364 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1606256979
transform 1 0 15548 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606256979
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1606256979
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1606256979
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_166
timestamp 1606256979
transform 1 0 16376 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_153
timestamp 1606256979
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1606256979
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 17572 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1606256979
transform 1 0 16560 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1606256979
transform 1 0 17112 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606256979
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_177
timestamp 1606256979
transform 1 0 17388 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_171
timestamp 1606256979
transform 1 0 16836 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_7_
timestamp 1606256979
transform 1 0 20056 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 19596 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1606256979
transform 1 0 18584 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1606256979
transform 1 0 19044 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_188
timestamp 1606256979
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_199
timestamp 1606256979
transform 1 0 19412 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_193
timestamp 1606256979
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_204
timestamp 1606256979
transform 1 0 19872 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1606256979
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606256979
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606256979
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606256979
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1606256979
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_218
timestamp 1606256979
transform 1 0 21160 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1606256979
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1606256979
transform 1 0 21252 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 1380 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1606256979
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606256979
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_12
timestamp 1606256979
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1606256979
transform 1 0 3404 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606256979
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1606256979
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1606256979
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_41
timestamp 1606256979
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_1_
timestamp 1606256979
transform 1 0 5060 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6256 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_52
timestamp 1606256979
transform 1 0 5888 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1606256979
transform 1 0 7268 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1606256979
transform 1 0 8556 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_65
timestamp 1606256979
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_76
timestamp 1606256979
transform 1 0 8096 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_80
timestamp 1606256979
transform 1 0 8464 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9936 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606256979
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1606256979
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_93
timestamp 1606256979
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _131_
timestamp 1606256979
transform 1 0 11132 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1606256979
transform 1 0 11684 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_105
timestamp 1606256979
transform 1 0 10764 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_113
timestamp 1606256979
transform 1 0 11500 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_124
timestamp 1606256979
transform 1 0 12512 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _128_
timestamp 1606256979
transform 1 0 12788 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1606256979
transform 1 0 14168 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_W_FTB01
timestamp 1606256979
transform 1 0 13432 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_28_131
timestamp 1606256979
transform 1 0 13156 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_140
timestamp 1606256979
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1606256979
transform 1 0 16284 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1606256979
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606256979
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1606256979
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_163
timestamp 1606256979
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1606256979
transform 1 0 17296 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1606256979
transform 1 0 18308 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_174
timestamp 1606256979
transform 1 0 17112 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_185
timestamp 1606256979
transform 1 0 18124 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18492 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_4_
timestamp 1606256979
transform 1 0 19504 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_198
timestamp 1606256979
transform 1 0 19320 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606256979
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606256979
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1606256979
transform 1 0 20332 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1606256979
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1606256979
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1606256979
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1606256979
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 2392 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606256979
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1606256979
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_11
timestamp 1606256979
transform 1 0 2116 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4048 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_30
timestamp 1606256979
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_41
timestamp 1606256979
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5060 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606256979
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606256979
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_62
timestamp 1606256979
transform 1 0 6808 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _135_
timestamp 1606256979
transform 1 0 6900 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 8464 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1606256979
transform 1 0 7452 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_67
timestamp 1606256979
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 1606256979
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 10672 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9476 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_89
timestamp 1606256979
transform 1 0 9292 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_100
timestamp 1606256979
transform 1 0 10304 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l4_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606256979
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1606256979
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13432 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_132
timestamp 1606256979
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_143
timestamp 1606256979
transform 1 0 14260 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1606256979
transform 1 0 15732 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l4_in_0_
timestamp 1606256979
transform 1 0 14720 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_147
timestamp 1606256979
transform 1 0 14628 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_157
timestamp 1606256979
transform 1 0 15548 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01
timestamp 1606256979
transform 1 0 17204 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1606256979
transform 1 0 16836 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1606256979
transform 1 0 18032 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606256979
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_168
timestamp 1606256979
transform 1 0 16560 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1606256979
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1606256979
transform 1 0 20240 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_6_
timestamp 1606256979
transform 1 0 18400 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_E_FTB01
timestamp 1606256979
transform 1 0 19504 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_197
timestamp 1606256979
transform 1 0 19228 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_206
timestamp 1606256979
transform 1 0 20056 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606256979
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_217
timestamp 1606256979
transform 1 0 21068 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1606256979
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1606256979
transform 1 0 1932 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l5_in_0_
timestamp 1606256979
transform 1 0 2944 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606256979
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1606256979
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1606256979
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606256979
transform 1 0 4048 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606256979
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1606256979
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _133_
timestamp 1606256979
transform 1 0 6716 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5704 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_48
timestamp 1606256979
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_59
timestamp 1606256979
transform 1 0 6532 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7360 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_30_65
timestamp 1606256979
transform 1 0 7084 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _132_
timestamp 1606256979
transform 1 0 9016 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 10672 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606256979
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_84
timestamp 1606256979
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1606256979
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1606256979
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 11408 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_110
timestamp 1606256979
transform 1 0 11224 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13064 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_128
timestamp 1606256979
transform 1 0 12880 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1606256979
transform 1 0 15272 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 15824 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606256979
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_146
timestamp 1606256979
transform 1 0 14536 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1606256979
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_158
timestamp 1606256979
transform 1 0 15640 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1606256979
transform 1 0 17480 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_1_E_FTB01
timestamp 1606256979
transform 1 0 18032 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_176
timestamp 1606256979
transform 1 0 17296 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_182
timestamp 1606256979
transform 1 0 17848 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1606256979
transform 1 0 19780 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1606256979
transform 1 0 18768 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_190
timestamp 1606256979
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_201
timestamp 1606256979
transform 1 0 19596 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606256979
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606256979
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1606256979
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606256979
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606256979
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_W_FTB01
timestamp 1606256979
transform 1 0 1656 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_W_FTB01
timestamp 1606256979
transform 1 0 2392 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606256979
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1606256979
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_12
timestamp 1606256979
transform 1 0 2208 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_20
timestamp 1606256979
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1606256979
transform 1 0 3128 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4784 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 3772 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_31_26
timestamp 1606256979
transform 1 0 3496 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_38
timestamp 1606256979
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606256979
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_56
timestamp 1606256979
transform 1 0 6256 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_60
timestamp 1606256979
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1606256979
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 6992 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_80
timestamp 1606256979
transform 1 0 8464 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8832 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 10488 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_100
timestamp 1606256979
transform 1 0 10304 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1606256979
transform 1 0 11316 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606256979
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_108
timestamp 1606256979
transform 1 0 11040 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1606256979
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _127_
timestamp 1606256979
transform 1 0 13432 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14352 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_132
timestamp 1606256979
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_138
timestamp 1606256979
transform 1 0 13800 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1606256979
transform 1 0 15640 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _129_
timestamp 1606256979
transform 1 0 15088 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16192 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_150
timestamp 1606256979
transform 1 0 14904 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_156
timestamp 1606256979
transform 1 0 15456 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_162
timestamp 1606256979
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1606256979
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_1_W_FTB01
timestamp 1606256979
transform 1 0 17204 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606256979
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_173
timestamp 1606256979
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1606256979
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 20148 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 18584 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_188
timestamp 1606256979
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_202
timestamp 1606256979
transform 1 0 19688 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_206
timestamp 1606256979
transform 1 0 20056 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606256979
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_216
timestamp 1606256979
transform 1 0 20976 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_2_W_FTB01
timestamp 1606256979
transform 1 0 1656 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_W_FTB01
timestamp 1606256979
transform 1 0 2392 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606256979
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1606256979
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_12
timestamp 1606256979
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_20
timestamp 1606256979
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 3220 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606256979
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1606256979
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_41
timestamp 1606256979
transform 1 0 4876 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 6072 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5060 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606256979
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_52
timestamp 1606256979
transform 1 0 5888 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_60
timestamp 1606256979
transform 1 0 6624 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6900 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_32_79
timestamp 1606256979
transform 1 0 8372 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9752 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606256979
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_90
timestamp 1606256979
transform 1 0 9384 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_103
timestamp 1606256979
transform 1 0 10580 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  clk_2_N_FTB01
timestamp 1606256979
transform 1 0 10764 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_1_
timestamp 1606256979
transform 1 0 11500 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 12604 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606256979
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_111
timestamp 1606256979
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1606256979
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1606256979
transform 1 0 13708 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_32_131
timestamp 1606256979
transform 1 0 13156 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1606256979
transform 1 0 14812 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1606256979
transform 1 0 15456 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606256979
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_146
timestamp 1606256979
transform 1 0 14536 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_153
timestamp 1606256979
transform 1 0 15180 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_165
timestamp 1606256979
transform 1 0 16284 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1606256979
transform 1 0 18308 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_2_E_FTB01
timestamp 1606256979
transform 1 0 16744 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1606256979
transform 1 0 17480 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606256979
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_169
timestamp 1606256979
transform 1 0 16652 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_176
timestamp 1606256979
transform 1 0 17296 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1606256979
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_E_FTB01
timestamp 1606256979
transform 1 0 19596 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_N_FTB01
timestamp 1606256979
transform 1 0 18860 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_191
timestamp 1606256979
transform 1 0 18676 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_199
timestamp 1606256979
transform 1 0 19412 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_207
timestamp 1606256979
transform 1 0 20148 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_E_FTB01
timestamp 1606256979
transform 1 0 20332 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606256979
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606256979
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1606256979
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606256979
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 18418 22320 18474 22800 6 Test_en_N_out
port 0 nsew default tristate
rlabel metal2 s 18878 0 18934 480 6 Test_en_S_in
port 1 nsew default input
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 2 nsew default input
rlabel metal2 s 570 0 626 480 6 bottom_left_grid_pin_43_
port 3 nsew default input
rlabel metal2 s 938 0 994 480 6 bottom_left_grid_pin_44_
port 4 nsew default input
rlabel metal2 s 1306 0 1362 480 6 bottom_left_grid_pin_45_
port 5 nsew default input
rlabel metal2 s 1674 0 1730 480 6 bottom_left_grid_pin_46_
port 6 nsew default input
rlabel metal2 s 2042 0 2098 480 6 bottom_left_grid_pin_47_
port 7 nsew default input
rlabel metal2 s 2410 0 2466 480 6 bottom_left_grid_pin_48_
port 8 nsew default input
rlabel metal2 s 2778 0 2834 480 6 bottom_left_grid_pin_49_
port 9 nsew default input
rlabel metal2 s 3146 0 3202 480 6 ccff_head
port 10 nsew default input
rlabel metal2 s 3514 0 3570 480 6 ccff_tail
port 11 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_in[0]
port 12 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[10]
port 13 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[11]
port 14 nsew default input
rlabel metal3 s 0 7896 480 8016 6 chanx_left_in[12]
port 15 nsew default input
rlabel metal3 s 0 8304 480 8424 6 chanx_left_in[13]
port 16 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[14]
port 17 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[15]
port 18 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_left_in[16]
port 19 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[17]
port 20 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[18]
port 21 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[19]
port 22 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[1]
port 23 nsew default input
rlabel metal3 s 0 3952 480 4072 6 chanx_left_in[2]
port 24 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[3]
port 25 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[4]
port 26 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_left_in[5]
port 27 nsew default input
rlabel metal3 s 0 5584 480 5704 6 chanx_left_in[6]
port 28 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[7]
port 29 nsew default input
rlabel metal3 s 0 6400 480 6520 6 chanx_left_in[8]
port 30 nsew default input
rlabel metal3 s 0 6808 480 6928 6 chanx_left_in[9]
port 31 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_left_out[0]
port 32 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 chanx_left_out[10]
port 33 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[11]
port 34 nsew default tristate
rlabel metal3 s 0 15784 480 15904 6 chanx_left_out[12]
port 35 nsew default tristate
rlabel metal3 s 0 16192 480 16312 6 chanx_left_out[13]
port 36 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[14]
port 37 nsew default tristate
rlabel metal3 s 0 17008 480 17128 6 chanx_left_out[15]
port 38 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 chanx_left_out[16]
port 39 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[17]
port 40 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[18]
port 41 nsew default tristate
rlabel metal3 s 0 18640 480 18760 6 chanx_left_out[19]
port 42 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[1]
port 43 nsew default tristate
rlabel metal3 s 0 11840 480 11960 6 chanx_left_out[2]
port 44 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_left_out[3]
port 45 nsew default tristate
rlabel metal3 s 0 12656 480 12776 6 chanx_left_out[4]
port 46 nsew default tristate
rlabel metal3 s 0 13064 480 13184 6 chanx_left_out[5]
port 47 nsew default tristate
rlabel metal3 s 0 13472 480 13592 6 chanx_left_out[6]
port 48 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[7]
port 49 nsew default tristate
rlabel metal3 s 0 14288 480 14408 6 chanx_left_out[8]
port 50 nsew default tristate
rlabel metal3 s 0 14696 480 14816 6 chanx_left_out[9]
port 51 nsew default tristate
rlabel metal3 s 22320 3272 22800 3392 6 chanx_right_in[0]
port 52 nsew default input
rlabel metal3 s 22320 7216 22800 7336 6 chanx_right_in[10]
port 53 nsew default input
rlabel metal3 s 22320 7624 22800 7744 6 chanx_right_in[11]
port 54 nsew default input
rlabel metal3 s 22320 7896 22800 8016 6 chanx_right_in[12]
port 55 nsew default input
rlabel metal3 s 22320 8304 22800 8424 6 chanx_right_in[13]
port 56 nsew default input
rlabel metal3 s 22320 8712 22800 8832 6 chanx_right_in[14]
port 57 nsew default input
rlabel metal3 s 22320 9120 22800 9240 6 chanx_right_in[15]
port 58 nsew default input
rlabel metal3 s 22320 9528 22800 9648 6 chanx_right_in[16]
port 59 nsew default input
rlabel metal3 s 22320 9936 22800 10056 6 chanx_right_in[17]
port 60 nsew default input
rlabel metal3 s 22320 10344 22800 10464 6 chanx_right_in[18]
port 61 nsew default input
rlabel metal3 s 22320 10752 22800 10872 6 chanx_right_in[19]
port 62 nsew default input
rlabel metal3 s 22320 3680 22800 3800 6 chanx_right_in[1]
port 63 nsew default input
rlabel metal3 s 22320 3952 22800 4072 6 chanx_right_in[2]
port 64 nsew default input
rlabel metal3 s 22320 4360 22800 4480 6 chanx_right_in[3]
port 65 nsew default input
rlabel metal3 s 22320 4768 22800 4888 6 chanx_right_in[4]
port 66 nsew default input
rlabel metal3 s 22320 5176 22800 5296 6 chanx_right_in[5]
port 67 nsew default input
rlabel metal3 s 22320 5584 22800 5704 6 chanx_right_in[6]
port 68 nsew default input
rlabel metal3 s 22320 5992 22800 6112 6 chanx_right_in[7]
port 69 nsew default input
rlabel metal3 s 22320 6400 22800 6520 6 chanx_right_in[8]
port 70 nsew default input
rlabel metal3 s 22320 6808 22800 6928 6 chanx_right_in[9]
port 71 nsew default input
rlabel metal3 s 22320 11160 22800 11280 6 chanx_right_out[0]
port 72 nsew default tristate
rlabel metal3 s 22320 15104 22800 15224 6 chanx_right_out[10]
port 73 nsew default tristate
rlabel metal3 s 22320 15376 22800 15496 6 chanx_right_out[11]
port 74 nsew default tristate
rlabel metal3 s 22320 15784 22800 15904 6 chanx_right_out[12]
port 75 nsew default tristate
rlabel metal3 s 22320 16192 22800 16312 6 chanx_right_out[13]
port 76 nsew default tristate
rlabel metal3 s 22320 16600 22800 16720 6 chanx_right_out[14]
port 77 nsew default tristate
rlabel metal3 s 22320 17008 22800 17128 6 chanx_right_out[15]
port 78 nsew default tristate
rlabel metal3 s 22320 17416 22800 17536 6 chanx_right_out[16]
port 79 nsew default tristate
rlabel metal3 s 22320 17824 22800 17944 6 chanx_right_out[17]
port 80 nsew default tristate
rlabel metal3 s 22320 18232 22800 18352 6 chanx_right_out[18]
port 81 nsew default tristate
rlabel metal3 s 22320 18640 22800 18760 6 chanx_right_out[19]
port 82 nsew default tristate
rlabel metal3 s 22320 11568 22800 11688 6 chanx_right_out[1]
port 83 nsew default tristate
rlabel metal3 s 22320 11840 22800 11960 6 chanx_right_out[2]
port 84 nsew default tristate
rlabel metal3 s 22320 12248 22800 12368 6 chanx_right_out[3]
port 85 nsew default tristate
rlabel metal3 s 22320 12656 22800 12776 6 chanx_right_out[4]
port 86 nsew default tristate
rlabel metal3 s 22320 13064 22800 13184 6 chanx_right_out[5]
port 87 nsew default tristate
rlabel metal3 s 22320 13472 22800 13592 6 chanx_right_out[6]
port 88 nsew default tristate
rlabel metal3 s 22320 13880 22800 14000 6 chanx_right_out[7]
port 89 nsew default tristate
rlabel metal3 s 22320 14288 22800 14408 6 chanx_right_out[8]
port 90 nsew default tristate
rlabel metal3 s 22320 14696 22800 14816 6 chanx_right_out[9]
port 91 nsew default tristate
rlabel metal2 s 3882 0 3938 480 6 chany_bottom_in[0]
port 92 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chany_bottom_in[10]
port 93 nsew default input
rlabel metal2 s 8022 0 8078 480 6 chany_bottom_in[11]
port 94 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[12]
port 95 nsew default input
rlabel metal2 s 8758 0 8814 480 6 chany_bottom_in[13]
port 96 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[14]
port 97 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[15]
port 98 nsew default input
rlabel metal2 s 9862 0 9918 480 6 chany_bottom_in[16]
port 99 nsew default input
rlabel metal2 s 10230 0 10286 480 6 chany_bottom_in[17]
port 100 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[18]
port 101 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[19]
port 102 nsew default input
rlabel metal2 s 4250 0 4306 480 6 chany_bottom_in[1]
port 103 nsew default input
rlabel metal2 s 4618 0 4674 480 6 chany_bottom_in[2]
port 104 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[3]
port 105 nsew default input
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_in[4]
port 106 nsew default input
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_in[5]
port 107 nsew default input
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_in[6]
port 108 nsew default input
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_in[7]
port 109 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[8]
port 110 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chany_bottom_in[9]
port 111 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_out[0]
port 112 nsew default tristate
rlabel metal2 s 15106 0 15162 480 6 chany_bottom_out[10]
port 113 nsew default tristate
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_out[11]
port 114 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_out[12]
port 115 nsew default tristate
rlabel metal2 s 16210 0 16266 480 6 chany_bottom_out[13]
port 116 nsew default tristate
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_out[14]
port 117 nsew default tristate
rlabel metal2 s 16946 0 17002 480 6 chany_bottom_out[15]
port 118 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_out[16]
port 119 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 chany_bottom_out[17]
port 120 nsew default tristate
rlabel metal2 s 18142 0 18198 480 6 chany_bottom_out[18]
port 121 nsew default tristate
rlabel metal2 s 18510 0 18566 480 6 chany_bottom_out[19]
port 122 nsew default tristate
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_out[1]
port 123 nsew default tristate
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_out[2]
port 124 nsew default tristate
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_out[3]
port 125 nsew default tristate
rlabel metal2 s 12898 0 12954 480 6 chany_bottom_out[4]
port 126 nsew default tristate
rlabel metal2 s 13266 0 13322 480 6 chany_bottom_out[5]
port 127 nsew default tristate
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_out[6]
port 128 nsew default tristate
rlabel metal2 s 14002 0 14058 480 6 chany_bottom_out[7]
port 129 nsew default tristate
rlabel metal2 s 14370 0 14426 480 6 chany_bottom_out[8]
port 130 nsew default tristate
rlabel metal2 s 14738 0 14794 480 6 chany_bottom_out[9]
port 131 nsew default tristate
rlabel metal2 s 3238 22320 3294 22800 6 chany_top_in[0]
port 132 nsew default input
rlabel metal2 s 7010 22320 7066 22800 6 chany_top_in[10]
port 133 nsew default input
rlabel metal2 s 7378 22320 7434 22800 6 chany_top_in[11]
port 134 nsew default input
rlabel metal2 s 7746 22320 7802 22800 6 chany_top_in[12]
port 135 nsew default input
rlabel metal2 s 8114 22320 8170 22800 6 chany_top_in[13]
port 136 nsew default input
rlabel metal2 s 8482 22320 8538 22800 6 chany_top_in[14]
port 137 nsew default input
rlabel metal2 s 8942 22320 8998 22800 6 chany_top_in[15]
port 138 nsew default input
rlabel metal2 s 9310 22320 9366 22800 6 chany_top_in[16]
port 139 nsew default input
rlabel metal2 s 9678 22320 9734 22800 6 chany_top_in[17]
port 140 nsew default input
rlabel metal2 s 10046 22320 10102 22800 6 chany_top_in[18]
port 141 nsew default input
rlabel metal2 s 10414 22320 10470 22800 6 chany_top_in[19]
port 142 nsew default input
rlabel metal2 s 3606 22320 3662 22800 6 chany_top_in[1]
port 143 nsew default input
rlabel metal2 s 3974 22320 4030 22800 6 chany_top_in[2]
port 144 nsew default input
rlabel metal2 s 4342 22320 4398 22800 6 chany_top_in[3]
port 145 nsew default input
rlabel metal2 s 4710 22320 4766 22800 6 chany_top_in[4]
port 146 nsew default input
rlabel metal2 s 5078 22320 5134 22800 6 chany_top_in[5]
port 147 nsew default input
rlabel metal2 s 5446 22320 5502 22800 6 chany_top_in[6]
port 148 nsew default input
rlabel metal2 s 5906 22320 5962 22800 6 chany_top_in[7]
port 149 nsew default input
rlabel metal2 s 6274 22320 6330 22800 6 chany_top_in[8]
port 150 nsew default input
rlabel metal2 s 6642 22320 6698 22800 6 chany_top_in[9]
port 151 nsew default input
rlabel metal2 s 10782 22320 10838 22800 6 chany_top_out[0]
port 152 nsew default tristate
rlabel metal2 s 14646 22320 14702 22800 6 chany_top_out[10]
port 153 nsew default tristate
rlabel metal2 s 15014 22320 15070 22800 6 chany_top_out[11]
port 154 nsew default tristate
rlabel metal2 s 15382 22320 15438 22800 6 chany_top_out[12]
port 155 nsew default tristate
rlabel metal2 s 15750 22320 15806 22800 6 chany_top_out[13]
port 156 nsew default tristate
rlabel metal2 s 16118 22320 16174 22800 6 chany_top_out[14]
port 157 nsew default tristate
rlabel metal2 s 16486 22320 16542 22800 6 chany_top_out[15]
port 158 nsew default tristate
rlabel metal2 s 16854 22320 16910 22800 6 chany_top_out[16]
port 159 nsew default tristate
rlabel metal2 s 17314 22320 17370 22800 6 chany_top_out[17]
port 160 nsew default tristate
rlabel metal2 s 17682 22320 17738 22800 6 chany_top_out[18]
port 161 nsew default tristate
rlabel metal2 s 18050 22320 18106 22800 6 chany_top_out[19]
port 162 nsew default tristate
rlabel metal2 s 11150 22320 11206 22800 6 chany_top_out[1]
port 163 nsew default tristate
rlabel metal2 s 11610 22320 11666 22800 6 chany_top_out[2]
port 164 nsew default tristate
rlabel metal2 s 11978 22320 12034 22800 6 chany_top_out[3]
port 165 nsew default tristate
rlabel metal2 s 12346 22320 12402 22800 6 chany_top_out[4]
port 166 nsew default tristate
rlabel metal2 s 12714 22320 12770 22800 6 chany_top_out[5]
port 167 nsew default tristate
rlabel metal2 s 13082 22320 13138 22800 6 chany_top_out[6]
port 168 nsew default tristate
rlabel metal2 s 13450 22320 13506 22800 6 chany_top_out[7]
port 169 nsew default tristate
rlabel metal2 s 13818 22320 13874 22800 6 chany_top_out[8]
port 170 nsew default tristate
rlabel metal2 s 14186 22320 14242 22800 6 chany_top_out[9]
port 171 nsew default tristate
rlabel metal3 s 22320 20544 22800 20664 6 clk_1_E_out
port 172 nsew default tristate
rlabel metal2 s 18786 22320 18842 22800 6 clk_1_N_in
port 173 nsew default input
rlabel metal2 s 19246 0 19302 480 6 clk_1_S_in
port 174 nsew default input
rlabel metal3 s 0 19048 480 19168 6 clk_1_W_out
port 175 nsew default tristate
rlabel metal3 s 22320 19048 22800 19168 6 clk_2_E_in
port 176 nsew default input
rlabel metal3 s 22320 20952 22800 21072 6 clk_2_E_out
port 177 nsew default tristate
rlabel metal2 s 19154 22320 19210 22800 6 clk_2_N_in
port 178 nsew default input
rlabel metal2 s 21454 22320 21510 22800 6 clk_2_N_out
port 179 nsew default tristate
rlabel metal2 s 19614 0 19670 480 6 clk_2_S_in
port 180 nsew default input
rlabel metal2 s 20350 0 20406 480 6 clk_2_S_out
port 181 nsew default tristate
rlabel metal3 s 0 21360 480 21480 6 clk_2_W_in
port 182 nsew default input
rlabel metal3 s 0 19320 480 19440 6 clk_2_W_out
port 183 nsew default tristate
rlabel metal3 s 22320 19320 22800 19440 6 clk_3_E_in
port 184 nsew default input
rlabel metal3 s 22320 21360 22800 21480 6 clk_3_E_out
port 185 nsew default tristate
rlabel metal2 s 19522 22320 19578 22800 6 clk_3_N_in
port 186 nsew default input
rlabel metal2 s 21822 22320 21878 22800 6 clk_3_N_out
port 187 nsew default tristate
rlabel metal2 s 19982 0 20038 480 6 clk_3_S_in
port 188 nsew default input
rlabel metal2 s 20718 0 20774 480 6 clk_3_S_out
port 189 nsew default tristate
rlabel metal3 s 0 21768 480 21888 6 clk_3_W_in
port 190 nsew default input
rlabel metal3 s 0 19728 480 19848 6 clk_3_W_out
port 191 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 192 nsew default input
rlabel metal3 s 0 416 480 536 6 left_bottom_grid_pin_35_
port 193 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_36_
port 194 nsew default input
rlabel metal3 s 0 1232 480 1352 6 left_bottom_grid_pin_37_
port 195 nsew default input
rlabel metal3 s 0 1640 480 1760 6 left_bottom_grid_pin_38_
port 196 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_39_
port 197 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_40_
port 198 nsew default input
rlabel metal3 s 0 2864 480 2984 6 left_bottom_grid_pin_41_
port 199 nsew default input
rlabel metal2 s 19890 22320 19946 22800 6 prog_clk_0_N_in
port 200 nsew default input
rlabel metal3 s 22320 21768 22800 21888 6 prog_clk_1_E_out
port 201 nsew default tristate
rlabel metal2 s 20350 22320 20406 22800 6 prog_clk_1_N_in
port 202 nsew default input
rlabel metal2 s 21086 0 21142 480 6 prog_clk_1_S_in
port 203 nsew default input
rlabel metal3 s 0 20136 480 20256 6 prog_clk_1_W_out
port 204 nsew default tristate
rlabel metal3 s 22320 19728 22800 19848 6 prog_clk_2_E_in
port 205 nsew default input
rlabel metal3 s 22320 22176 22800 22296 6 prog_clk_2_E_out
port 206 nsew default tristate
rlabel metal2 s 20718 22320 20774 22800 6 prog_clk_2_N_in
port 207 nsew default input
rlabel metal2 s 22190 22320 22246 22800 6 prog_clk_2_N_out
port 208 nsew default tristate
rlabel metal2 s 21454 0 21510 480 6 prog_clk_2_S_in
port 209 nsew default input
rlabel metal2 s 22190 0 22246 480 6 prog_clk_2_S_out
port 210 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 prog_clk_2_W_in
port 211 nsew default input
rlabel metal3 s 0 20544 480 20664 6 prog_clk_2_W_out
port 212 nsew default tristate
rlabel metal3 s 22320 20136 22800 20256 6 prog_clk_3_E_in
port 213 nsew default input
rlabel metal3 s 22320 22584 22800 22704 6 prog_clk_3_E_out
port 214 nsew default tristate
rlabel metal2 s 21086 22320 21142 22800 6 prog_clk_3_N_in
port 215 nsew default input
rlabel metal2 s 22558 22320 22614 22800 6 prog_clk_3_N_out
port 216 nsew default tristate
rlabel metal2 s 21822 0 21878 480 6 prog_clk_3_S_in
port 217 nsew default input
rlabel metal2 s 22558 0 22614 480 6 prog_clk_3_S_out
port 218 nsew default tristate
rlabel metal3 s 0 22584 480 22704 6 prog_clk_3_W_in
port 219 nsew default input
rlabel metal3 s 0 20952 480 21072 6 prog_clk_3_W_out
port 220 nsew default tristate
rlabel metal3 s 22320 144 22800 264 6 right_bottom_grid_pin_34_
port 221 nsew default input
rlabel metal3 s 22320 416 22800 536 6 right_bottom_grid_pin_35_
port 222 nsew default input
rlabel metal3 s 22320 824 22800 944 6 right_bottom_grid_pin_36_
port 223 nsew default input
rlabel metal3 s 22320 1232 22800 1352 6 right_bottom_grid_pin_37_
port 224 nsew default input
rlabel metal3 s 22320 1640 22800 1760 6 right_bottom_grid_pin_38_
port 225 nsew default input
rlabel metal3 s 22320 2048 22800 2168 6 right_bottom_grid_pin_39_
port 226 nsew default input
rlabel metal3 s 22320 2456 22800 2576 6 right_bottom_grid_pin_40_
port 227 nsew default input
rlabel metal3 s 22320 2864 22800 2984 6 right_bottom_grid_pin_41_
port 228 nsew default input
rlabel metal2 s 202 22320 258 22800 6 top_left_grid_pin_42_
port 229 nsew default input
rlabel metal2 s 570 22320 626 22800 6 top_left_grid_pin_43_
port 230 nsew default input
rlabel metal2 s 938 22320 994 22800 6 top_left_grid_pin_44_
port 231 nsew default input
rlabel metal2 s 1306 22320 1362 22800 6 top_left_grid_pin_45_
port 232 nsew default input
rlabel metal2 s 1674 22320 1730 22800 6 top_left_grid_pin_46_
port 233 nsew default input
rlabel metal2 s 2042 22320 2098 22800 6 top_left_grid_pin_47_
port 234 nsew default input
rlabel metal2 s 2410 22320 2466 22800 6 top_left_grid_pin_48_
port 235 nsew default input
rlabel metal2 s 2778 22320 2834 22800 6 top_left_grid_pin_49_
port 236 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 237 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 238 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
