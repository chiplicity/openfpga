VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__0_
  CLASS BLOCK ;
  FOREIGN cbx_1__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 80.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 2.400 2.680 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 2.400 6.760 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 77.600 9.110 80.000 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 2.400 11.520 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 2.760 200.000 3.360 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 8.200 200.000 8.800 ;
    END
  END address[6]
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 13.640 200.000 14.240 ;
    END
  END bottom_grid_pin_0_
  PIN bottom_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.170 77.600 45.450 80.000 ;
    END
  END bottom_grid_pin_10_
  PIN bottom_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 2.400 16.280 ;
    END
  END bottom_grid_pin_12_
  PIN bottom_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 2.400 21.040 ;
    END
  END bottom_grid_pin_14_
  PIN bottom_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 2.400 ;
    END
  END bottom_grid_pin_2_
  PIN bottom_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 2.400 ;
    END
  END bottom_grid_pin_4_
  PIN bottom_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.770 77.600 27.050 80.000 ;
    END
  END bottom_grid_pin_6_
  PIN bottom_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 19.760 200.000 20.360 ;
    END
  END bottom_grid_pin_8_
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 25.200 200.000 25.800 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.110 77.600 63.390 80.000 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 31.320 200.000 31.920 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 2.400 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 2.400 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 2.400 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 2.400 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 2.400 30.560 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 2.400 35.320 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 36.760 200.000 37.360 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 42.880 200.000 43.480 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 2.400 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.510 77.600 81.790 80.000 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.450 77.600 99.730 80.000 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 48.320 200.000 48.920 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 2.400 40.080 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 2.400 44.840 ;
    END
  END chanx_left_out[8]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 2.400 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 2.400 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 2.400 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.850 77.600 118.130 80.000 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 2.400 49.600 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 77.600 136.070 80.000 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 154.190 77.600 154.470 80.000 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 53.760 200.000 54.360 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 2.400 54.360 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 2.400 59.120 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 2.400 63.880 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 2.400 68.640 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 172.130 77.600 172.410 80.000 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 59.880 200.000 60.480 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 65.320 200.000 65.920 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 71.440 200.000 72.040 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 2.400 78.160 ;
    END
  END chanx_right_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END enable
  PIN top_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.530 77.600 190.810 80.000 ;
    END
  END top_grid_pin_14_
  PIN top_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 76.880 200.000 77.480 ;
    END
  END top_grid_pin_2_
  PIN top_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 2.400 ;
    END
  END top_grid_pin_6_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 38.055 10.640 39.655 68.240 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 71.385 10.640 72.985 68.240 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 68.085 ;
      LAYER met1 ;
        RECT 0.070 0.380 198.190 68.240 ;
      LAYER met2 ;
        RECT 0.090 77.320 8.550 77.930 ;
        RECT 9.390 77.320 26.490 77.930 ;
        RECT 27.330 77.320 44.890 77.930 ;
        RECT 45.730 77.320 62.830 77.930 ;
        RECT 63.670 77.320 81.230 77.930 ;
        RECT 82.070 77.320 99.170 77.930 ;
        RECT 100.010 77.320 117.570 77.930 ;
        RECT 118.410 77.320 135.510 77.930 ;
        RECT 136.350 77.320 153.910 77.930 ;
        RECT 154.750 77.320 171.850 77.930 ;
        RECT 172.690 77.320 190.250 77.930 ;
        RECT 191.090 77.320 198.170 77.930 ;
        RECT 0.090 2.680 198.170 77.320 ;
        RECT 0.090 0.270 6.710 2.680 ;
        RECT 7.550 0.270 20.970 2.680 ;
        RECT 21.810 0.270 35.230 2.680 ;
        RECT 36.070 0.270 49.490 2.680 ;
        RECT 50.330 0.270 63.750 2.680 ;
        RECT 64.590 0.270 78.010 2.680 ;
        RECT 78.850 0.270 92.270 2.680 ;
        RECT 93.110 0.270 106.530 2.680 ;
        RECT 107.370 0.270 120.790 2.680 ;
        RECT 121.630 0.270 135.050 2.680 ;
        RECT 135.890 0.270 149.310 2.680 ;
        RECT 150.150 0.270 163.570 2.680 ;
        RECT 164.410 0.270 177.830 2.680 ;
        RECT 178.670 0.270 192.090 2.680 ;
        RECT 192.930 0.270 198.170 2.680 ;
      LAYER met3 ;
        RECT 2.800 77.160 197.200 77.560 ;
        RECT 0.270 76.480 197.200 77.160 ;
        RECT 0.270 73.800 198.450 76.480 ;
        RECT 2.800 72.440 198.450 73.800 ;
        RECT 2.800 72.400 197.200 72.440 ;
        RECT 0.270 71.040 197.200 72.400 ;
        RECT 0.270 69.040 198.450 71.040 ;
        RECT 2.800 67.640 198.450 69.040 ;
        RECT 0.270 66.320 198.450 67.640 ;
        RECT 0.270 64.920 197.200 66.320 ;
        RECT 0.270 64.280 198.450 64.920 ;
        RECT 2.800 62.880 198.450 64.280 ;
        RECT 0.270 60.880 198.450 62.880 ;
        RECT 0.270 59.520 197.200 60.880 ;
        RECT 2.800 59.480 197.200 59.520 ;
        RECT 2.800 58.120 198.450 59.480 ;
        RECT 0.270 54.760 198.450 58.120 ;
        RECT 2.800 53.360 197.200 54.760 ;
        RECT 0.270 50.000 198.450 53.360 ;
        RECT 2.800 49.320 198.450 50.000 ;
        RECT 2.800 48.600 197.200 49.320 ;
        RECT 0.270 47.920 197.200 48.600 ;
        RECT 0.270 45.240 198.450 47.920 ;
        RECT 2.800 43.880 198.450 45.240 ;
        RECT 2.800 43.840 197.200 43.880 ;
        RECT 0.270 42.480 197.200 43.840 ;
        RECT 0.270 40.480 198.450 42.480 ;
        RECT 2.800 39.080 198.450 40.480 ;
        RECT 0.270 37.760 198.450 39.080 ;
        RECT 0.270 36.360 197.200 37.760 ;
        RECT 0.270 35.720 198.450 36.360 ;
        RECT 2.800 34.320 198.450 35.720 ;
        RECT 0.270 32.320 198.450 34.320 ;
        RECT 0.270 30.960 197.200 32.320 ;
        RECT 2.800 30.920 197.200 30.960 ;
        RECT 2.800 29.560 198.450 30.920 ;
        RECT 0.270 26.200 198.450 29.560 ;
        RECT 2.800 24.800 197.200 26.200 ;
        RECT 0.270 21.440 198.450 24.800 ;
        RECT 2.800 20.760 198.450 21.440 ;
        RECT 2.800 20.040 197.200 20.760 ;
        RECT 0.270 19.360 197.200 20.040 ;
        RECT 0.270 16.680 198.450 19.360 ;
        RECT 2.800 15.280 198.450 16.680 ;
        RECT 0.270 14.640 198.450 15.280 ;
        RECT 0.270 13.240 197.200 14.640 ;
        RECT 0.270 11.920 198.450 13.240 ;
        RECT 2.800 10.520 198.450 11.920 ;
        RECT 0.270 9.200 198.450 10.520 ;
        RECT 0.270 7.800 197.200 9.200 ;
        RECT 0.270 7.160 198.450 7.800 ;
        RECT 2.800 5.760 198.450 7.160 ;
        RECT 0.270 3.760 198.450 5.760 ;
        RECT 0.270 3.080 197.200 3.760 ;
        RECT 2.800 2.360 197.200 3.080 ;
        RECT 2.800 1.680 198.450 2.360 ;
        RECT 0.270 0.855 198.450 1.680 ;
      LAYER met4 ;
        RECT 0.295 10.640 37.655 68.240 ;
        RECT 40.055 10.640 70.985 68.240 ;
        RECT 73.385 10.640 198.425 68.240 ;
  END
END cbx_1__0_
END LIBRARY

